module top(n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n78245, n78246, n78247, n78248, n78249, n78250, n78251, n78252, n78253, n78254, n78255, n78256, n78257, n78258, n78259, n78260, n78261, n78262, n78263, n78264, n78265, n78266, n78267, n78268, n78269, n78270, n78271, n78272, n78273, n78274, n78275, n78276, n78277, n78278, n78279, n78280, n78281, n78282, n78283, n78284, n78285, n78286, n78287, n78288, n78289, n78290, n78291, n78292, n78293, n78294, n78295, n78296, n78297, n78298, n78299, n78300, n78301, n78302, n78303, n78304, n78305, n78306, n78307, n78308, n78309, n78310, n78311, n78312, n78313, n78314, n78315, n78316, n78317, n78318, n78319, n78320, n78321, n78322, n78323, n78324, n78325, n78326, n78327, n78328, n78329, n78330, n78331, n78332, n78333, n78334, n78335, n78336, n78337, n78338, n78339, n78340, n78341, n78342, n78343, n78344, n78345, n78346, n78347, n78348, n78349, n78350, n78351, n78352, n78353, n78354, n78355, n78356, n78357, n78358, n78359, n78360, n78361, n78362, n78363, n78364, n78365, n78366, n78367, n78368, n78369, n78370, n78371, n78372);
  input n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511;
  output n78245, n78246, n78247, n78248, n78249, n78250, n78251, n78252, n78253, n78254, n78255, n78256, n78257, n78258, n78259, n78260, n78261, n78262, n78263, n78264, n78265, n78266, n78267, n78268, n78269, n78270, n78271, n78272, n78273, n78274, n78275, n78276, n78277, n78278, n78279, n78280, n78281, n78282, n78283, n78284, n78285, n78286, n78287, n78288, n78289, n78290, n78291, n78292, n78293, n78294, n78295, n78296, n78297, n78298, n78299, n78300, n78301, n78302, n78303, n78304, n78305, n78306, n78307, n78308, n78309, n78310, n78311, n78312, n78313, n78314, n78315, n78316, n78317, n78318, n78319, n78320, n78321, n78322, n78323, n78324, n78325, n78326, n78327, n78328, n78329, n78330, n78331, n78332, n78333, n78334, n78335, n78336, n78337, n78338, n78339, n78340, n78341, n78342, n78343, n78344, n78345, n78346, n78347, n78348, n78349, n78350, n78351, n78352, n78353, n78354, n78355, n78356, n78357, n78358, n78359, n78360, n78361, n78362, n78363, n78364, n78365, n78366, n78367, n78368, n78369, n78370, n78371, n78372;
  wire n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105, n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249, n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273, n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281, n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289, n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353, n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425, n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489, n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537, n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601, n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609, n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633, n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705, n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777, n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849, n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321, n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681, n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753, n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801, n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809, n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873, n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945, n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969, n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977, n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985, n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993, n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001, n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025, n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041, n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049, n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081, n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089, n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097, n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113, n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121, n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153, n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161, n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169, n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185, n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193, n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201, n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225, n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233, n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257, n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265, n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289, n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297, n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321, n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329, n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337, n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353, n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369, n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377, n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401, n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409, n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425, n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441, n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449, n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473, n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481, n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505, n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513, n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545, n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553, n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697, n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713, n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729, n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777, n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801, n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825, n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857, n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865, n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873, n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897, n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905, n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921, n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929, n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945, n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953, n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977, n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001, n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017, n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025, n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041, n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049, n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065, n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073, n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089, n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097, n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121, n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145, n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161, n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185, n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193, n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201, n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209, n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217, n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225, n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233, n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241, n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257, n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273, n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281, n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289, n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297, n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305, n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313, n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337, n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345, n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353, n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361, n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369, n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377, n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385, n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393, n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401, n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409, n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417, n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425, n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433, n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441, n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449, n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457, n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465, n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473, n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481, n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489, n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497, n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505, n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513, n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529, n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537, n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545, n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553, n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561, n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569, n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577, n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585, n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593, n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601, n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609, n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617, n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625, n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633, n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641, n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649, n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657, n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665, n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673, n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681, n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689, n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697, n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705, n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713, n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721, n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729, n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737, n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745, n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753, n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761, n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769, n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777, n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785, n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793, n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801, n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809, n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817, n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825, n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833, n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841, n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849, n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857, n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865, n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873, n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881, n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889, n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897, n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905, n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913, n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921, n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929, n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937, n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945, n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953, n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961, n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969, n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985, n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993, n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001, n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009, n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017, n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025, n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033, n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041, n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049, n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057, n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065, n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073, n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081, n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089, n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097, n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105, n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113, n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121, n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129, n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137, n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145, n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153, n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161, n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169, n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177, n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185, n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193, n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201, n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209, n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217, n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225, n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233, n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241, n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249, n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257, n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265, n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273, n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281, n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289, n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297, n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305, n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313, n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321, n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329, n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337, n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345, n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353, n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361, n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369, n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377, n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385, n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393, n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401, n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409, n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417, n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425, n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433, n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441, n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449, n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457, n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465, n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473, n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489, n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497, n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505, n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513, n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521, n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529, n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537, n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545, n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561, n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569, n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577, n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585, n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593, n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601, n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609, n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617, n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625, n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633, n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641, n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649, n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657, n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665, n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673, n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681, n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689, n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697, n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705, n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713, n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721, n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729, n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737, n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745, n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753, n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761, n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769, n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777, n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785, n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793, n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801, n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809, n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817, n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825, n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833, n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841, n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849, n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857, n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865, n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873, n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881, n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889, n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897, n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905, n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913, n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921, n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929, n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937, n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945, n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953, n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961, n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969, n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977, n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985, n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993, n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001, n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009, n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017, n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025, n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033, n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041, n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049, n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057, n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065, n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073, n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081, n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089, n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097, n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105, n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113, n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121, n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129, n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137, n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145, n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153, n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161, n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169, n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177, n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185, n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193, n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201, n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209, n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217, n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225, n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233, n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241, n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249, n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257, n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265, n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273, n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281, n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289, n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297, n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305, n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313, n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321, n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329, n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337, n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345, n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353, n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361, n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369, n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377, n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385, n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393, n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409, n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417, n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425, n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433, n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441, n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449, n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457, n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465, n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473, n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481, n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489, n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497, n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505, n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513, n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521, n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537, n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545, n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553, n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561, n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569, n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577, n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585, n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593, n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601, n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609, n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617, n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625, n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633, n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641, n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649, n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657, n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665, n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673, n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681, n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689, n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697, n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705, n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713, n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721, n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729, n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737, n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745, n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753, n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761, n29762, n29763, n29764, n29765, n29766, n29767, n29768, n29769, n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777, n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785, n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793, n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801, n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809, n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817, n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825, n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833, n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841, n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849, n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857, n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865, n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873, n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881, n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889, n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897, n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905, n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913, n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921, n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929, n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937, n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945, n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953, n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961, n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969, n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977, n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985, n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993, n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001, n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009, n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017, n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025, n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033, n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041, n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049, n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057, n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065, n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073, n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081, n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089, n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097, n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105, n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113, n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121, n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129, n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137, n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145, n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153, n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161, n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169, n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177, n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193, n30194, n30195, n30196, n30197, n30198, n30199, n30200, n30201, n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209, n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217, n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225, n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233, n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241, n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249, n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257, n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265, n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273, n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281, n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289, n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297, n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305, n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313, n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321, n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329, n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337, n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345, n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353, n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361, n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369, n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377, n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385, n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393, n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401, n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409, n30410, n30411, n30412, n30413, n30414, n30415, n30416, n30417, n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425, n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433, n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441, n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449, n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457, n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465, n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473, n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481, n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489, n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497, n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505, n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513, n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521, n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529, n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537, n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545, n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553, n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561, n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569, n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577, n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585, n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593, n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601, n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609, n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617, n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625, n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633, n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641, n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649, n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657, n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665, n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673, n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681, n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689, n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697, n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705, n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713, n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721, n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729, n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737, n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745, n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753, n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761, n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769, n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777, n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785, n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793, n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801, n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809, n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817, n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825, n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833, n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841, n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849, n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857, n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865, n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873, n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881, n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889, n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897, n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905, n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913, n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921, n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929, n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937, n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945, n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953, n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961, n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969, n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977, n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985, n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993, n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001, n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009, n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017, n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025, n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033, n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041, n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049, n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057, n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065, n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073, n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081, n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089, n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097, n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105, n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113, n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121, n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129, n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137, n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145, n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153, n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161, n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169, n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177, n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185, n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193, n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201, n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209, n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217, n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225, n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233, n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241, n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249, n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257, n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265, n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273, n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281, n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289, n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297, n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305, n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313, n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321, n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329, n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337, n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345, n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353, n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361, n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369, n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377, n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385, n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393, n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401, n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409, n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417, n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425, n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433, n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441, n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449, n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457, n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465, n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473, n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481, n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489, n31490, n31491, n31492, n31493, n31494, n31495, n31496, n31497, n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505, n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513, n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521, n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529, n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537, n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545, n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553, n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561, n31562, n31563, n31564, n31565, n31566, n31567, n31568, n31569, n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577, n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585, n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593, n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601, n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609, n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617, n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625, n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633, n31634, n31635, n31636, n31637, n31638, n31639, n31640, n31641, n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649, n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657, n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665, n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673, n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681, n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689, n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697, n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705, n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713, n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721, n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729, n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737, n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745, n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753, n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761, n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769, n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777, n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785, n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793, n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801, n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809, n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817, n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825, n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833, n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841, n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849, n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857, n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865, n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873, n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881, n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889, n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897, n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905, n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913, n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921, n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929, n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937, n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945, n31946, n31947, n31948, n31949, n31950, n31951, n31952, n31953, n31954, n31955, n31956, n31957, n31958, n31959, n31960, n31961, n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969, n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977, n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985, n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993, n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001, n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009, n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017, n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025, n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033, n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041, n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049, n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057, n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065, n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073, n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081, n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089, n32090, n32091, n32092, n32093, n32094, n32095, n32096, n32097, n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105, n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113, n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121, n32122, n32123, n32124, n32125, n32126, n32127, n32128, n32129, n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137, n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145, n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153, n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161, n32162, n32163, n32164, n32165, n32166, n32167, n32168, n32169, n32170, n32171, n32172, n32173, n32174, n32175, n32176, n32177, n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185, n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193, n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201, n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209, n32210, n32211, n32212, n32213, n32214, n32215, n32216, n32217, n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225, n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233, n32234, n32235, n32236, n32237, n32238, n32239, n32240, n32241, n32242, n32243, n32244, n32245, n32246, n32247, n32248, n32249, n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257, n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265, n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273, n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281, n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289, n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297, n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305, n32306, n32307, n32308, n32309, n32310, n32311, n32312, n32313, n32314, n32315, n32316, n32317, n32318, n32319, n32320, n32321, n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329, n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337, n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345, n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353, n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361, n32362, n32363, n32364, n32365, n32366, n32367, n32368, n32369, n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377, n32378, n32379, n32380, n32381, n32382, n32383, n32384, n32385, n32386, n32387, n32388, n32389, n32390, n32391, n32392, n32393, n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401, n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409, n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417, n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425, n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32433, n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32441, n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449, n32450, n32451, n32452, n32453, n32454, n32455, n32456, n32457, n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465, n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473, n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481, n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489, n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497, n32498, n32499, n32500, n32501, n32502, n32503, n32504, n32505, n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513, n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521, n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529, n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537, n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545, n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553, n32554, n32555, n32556, n32557, n32558, n32559, n32560, n32561, n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569, n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577, n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585, n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593, n32594, n32595, n32596, n32597, n32598, n32599, n32600, n32601, n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609, n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617, n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625, n32626, n32627, n32628, n32629, n32630, n32631, n32632, n32633, n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641, n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649, n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657, n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665, n32666, n32667, n32668, n32669, n32670, n32671, n32672, n32673, n32674, n32675, n32676, n32677, n32678, n32679, n32680, n32681, n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689, n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697, n32698, n32699, n32700, n32701, n32702, n32703, n32704, n32705, n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713, n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721, n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729, n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737, n32738, n32739, n32740, n32741, n32742, n32743, n32744, n32745, n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753, n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761, n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769, n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777, n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785, n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793, n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801, n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809, n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817, n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825, n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833, n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841, n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849, n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857, n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865, n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873, n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881, n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889, n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897, n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905, n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913, n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921, n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929, n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937, n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945, n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953, n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961, n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969, n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977, n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985, n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993, n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001, n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009, n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017, n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025, n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033, n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041, n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049, n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057, n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065, n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073, n33074, n33075, n33076, n33077, n33078, n33079, n33080, n33081, n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089, n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097, n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105, n33106, n33107, n33108, n33109, n33110, n33111, n33112, n33113, n33114, n33115, n33116, n33117, n33118, n33119, n33120, n33121, n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129, n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137, n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145, n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153, n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161, n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169, n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177, n33178, n33179, n33180, n33181, n33182, n33183, n33184, n33185, n33186, n33187, n33188, n33189, n33190, n33191, n33192, n33193, n33194, n33195, n33196, n33197, n33198, n33199, n33200, n33201, n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209, n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217, n33218, n33219, n33220, n33221, n33222, n33223, n33224, n33225, n33226, n33227, n33228, n33229, n33230, n33231, n33232, n33233, n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241, n33242, n33243, n33244, n33245, n33246, n33247, n33248, n33249, n33250, n33251, n33252, n33253, n33254, n33255, n33256, n33257, n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265, n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273, n33274, n33275, n33276, n33277, n33278, n33279, n33280, n33281, n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289, n33290, n33291, n33292, n33293, n33294, n33295, n33296, n33297, n33298, n33299, n33300, n33301, n33302, n33303, n33304, n33305, n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313, n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321, n33322, n33323, n33324, n33325, n33326, n33327, n33328, n33329, n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337, n33338, n33339, n33340, n33341, n33342, n33343, n33344, n33345, n33346, n33347, n33348, n33349, n33350, n33351, n33352, n33353, n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361, n33362, n33363, n33364, n33365, n33366, n33367, n33368, n33369, n33370, n33371, n33372, n33373, n33374, n33375, n33376, n33377, n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385, n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393, n33394, n33395, n33396, n33397, n33398, n33399, n33400, n33401, n33402, n33403, n33404, n33405, n33406, n33407, n33408, n33409, n33410, n33411, n33412, n33413, n33414, n33415, n33416, n33417, n33418, n33419, n33420, n33421, n33422, n33423, n33424, n33425, n33426, n33427, n33428, n33429, n33430, n33431, n33432, n33433, n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441, n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449, n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457, n33458, n33459, n33460, n33461, n33462, n33463, n33464, n33465, n33466, n33467, n33468, n33469, n33470, n33471, n33472, n33473, n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481, n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489, n33490, n33491, n33492, n33493, n33494, n33495, n33496, n33497, n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505, n33506, n33507, n33508, n33509, n33510, n33511, n33512, n33513, n33514, n33515, n33516, n33517, n33518, n33519, n33520, n33521, n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529, n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537, n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545, n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553, n33554, n33555, n33556, n33557, n33558, n33559, n33560, n33561, n33562, n33563, n33564, n33565, n33566, n33567, n33568, n33569, n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577, n33578, n33579, n33580, n33581, n33582, n33583, n33584, n33585, n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593, n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601, n33602, n33603, n33604, n33605, n33606, n33607, n33608, n33609, n33610, n33611, n33612, n33613, n33614, n33615, n33616, n33617, n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625, n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633, n33634, n33635, n33636, n33637, n33638, n33639, n33640, n33641, n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649, n33650, n33651, n33652, n33653, n33654, n33655, n33656, n33657, n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665, n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673, n33674, n33675, n33676, n33677, n33678, n33679, n33680, n33681, n33682, n33683, n33684, n33685, n33686, n33687, n33688, n33689, n33690, n33691, n33692, n33693, n33694, n33695, n33696, n33697, n33698, n33699, n33700, n33701, n33702, n33703, n33704, n33705, n33706, n33707, n33708, n33709, n33710, n33711, n33712, n33713, n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721, n33722, n33723, n33724, n33725, n33726, n33727, n33728, n33729, n33730, n33731, n33732, n33733, n33734, n33735, n33736, n33737, n33738, n33739, n33740, n33741, n33742, n33743, n33744, n33745, n33746, n33747, n33748, n33749, n33750, n33751, n33752, n33753, n33754, n33755, n33756, n33757, n33758, n33759, n33760, n33761, n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769, n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777, n33778, n33779, n33780, n33781, n33782, n33783, n33784, n33785, n33786, n33787, n33788, n33789, n33790, n33791, n33792, n33793, n33794, n33795, n33796, n33797, n33798, n33799, n33800, n33801, n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809, n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817, n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825, n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833, n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841, n33842, n33843, n33844, n33845, n33846, n33847, n33848, n33849, n33850, n33851, n33852, n33853, n33854, n33855, n33856, n33857, n33858, n33859, n33860, n33861, n33862, n33863, n33864, n33865, n33866, n33867, n33868, n33869, n33870, n33871, n33872, n33873, n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881, n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889, n33890, n33891, n33892, n33893, n33894, n33895, n33896, n33897, n33898, n33899, n33900, n33901, n33902, n33903, n33904, n33905, n33906, n33907, n33908, n33909, n33910, n33911, n33912, n33913, n33914, n33915, n33916, n33917, n33918, n33919, n33920, n33921, n33922, n33923, n33924, n33925, n33926, n33927, n33928, n33929, n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937, n33938, n33939, n33940, n33941, n33942, n33943, n33944, n33945, n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953, n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961, n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969, n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977, n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985, n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993, n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001, n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009, n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017, n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025, n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033, n34034, n34035, n34036, n34037, n34038, n34039, n34040, n34041, n34042, n34043, n34044, n34045, n34046, n34047, n34048, n34049, n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057, n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065, n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073, n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081, n34082, n34083, n34084, n34085, n34086, n34087, n34088, n34089, n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097, n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105, n34106, n34107, n34108, n34109, n34110, n34111, n34112, n34113, n34114, n34115, n34116, n34117, n34118, n34119, n34120, n34121, n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129, n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137, n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145, n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153, n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161, n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169, n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177, n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185, n34186, n34187, n34188, n34189, n34190, n34191, n34192, n34193, n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201, n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209, n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217, n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225, n34226, n34227, n34228, n34229, n34230, n34231, n34232, n34233, n34234, n34235, n34236, n34237, n34238, n34239, n34240, n34241, n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249, n34250, n34251, n34252, n34253, n34254, n34255, n34256, n34257, n34258, n34259, n34260, n34261, n34262, n34263, n34264, n34265, n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273, n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281, n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289, n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297, n34298, n34299, n34300, n34301, n34302, n34303, n34304, n34305, n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313, n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321, n34322, n34323, n34324, n34325, n34326, n34327, n34328, n34329, n34330, n34331, n34332, n34333, n34334, n34335, n34336, n34337, n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345, n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353, n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361, n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369, n34370, n34371, n34372, n34373, n34374, n34375, n34376, n34377, n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385, n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393, n34394, n34395, n34396, n34397, n34398, n34399, n34400, n34401, n34402, n34403, n34404, n34405, n34406, n34407, n34408, n34409, n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417, n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425, n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433, n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441, n34442, n34443, n34444, n34445, n34446, n34447, n34448, n34449, n34450, n34451, n34452, n34453, n34454, n34455, n34456, n34457, n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465, n34466, n34467, n34468, n34469, n34470, n34471, n34472, n34473, n34474, n34475, n34476, n34477, n34478, n34479, n34480, n34481, n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489, n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497, n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505, n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513, n34514, n34515, n34516, n34517, n34518, n34519, n34520, n34521, n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529, n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537, n34538, n34539, n34540, n34541, n34542, n34543, n34544, n34545, n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553, n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561, n34562, n34563, n34564, n34565, n34566, n34567, n34568, n34569, n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577, n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585, n34586, n34587, n34588, n34589, n34590, n34591, n34592, n34593, n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601, n34602, n34603, n34604, n34605, n34606, n34607, n34608, n34609, n34610, n34611, n34612, n34613, n34614, n34615, n34616, n34617, n34618, n34619, n34620, n34621, n34622, n34623, n34624, n34625, n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633, n34634, n34635, n34636, n34637, n34638, n34639, n34640, n34641, n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649, n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657, n34658, n34659, n34660, n34661, n34662, n34663, n34664, n34665, n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673, n34674, n34675, n34676, n34677, n34678, n34679, n34680, n34681, n34682, n34683, n34684, n34685, n34686, n34687, n34688, n34689, n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697, n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705, n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713, n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721, n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729, n34730, n34731, n34732, n34733, n34734, n34735, n34736, n34737, n34738, n34739, n34740, n34741, n34742, n34743, n34744, n34745, n34746, n34747, n34748, n34749, n34750, n34751, n34752, n34753, n34754, n34755, n34756, n34757, n34758, n34759, n34760, n34761, n34762, n34763, n34764, n34765, n34766, n34767, n34768, n34769, n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777, n34778, n34779, n34780, n34781, n34782, n34783, n34784, n34785, n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793, n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801, n34802, n34803, n34804, n34805, n34806, n34807, n34808, n34809, n34810, n34811, n34812, n34813, n34814, n34815, n34816, n34817, n34818, n34819, n34820, n34821, n34822, n34823, n34824, n34825, n34826, n34827, n34828, n34829, n34830, n34831, n34832, n34833, n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841, n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849, n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857, n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865, n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873, n34874, n34875, n34876, n34877, n34878, n34879, n34880, n34881, n34882, n34883, n34884, n34885, n34886, n34887, n34888, n34889, n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897, n34898, n34899, n34900, n34901, n34902, n34903, n34904, n34905, n34906, n34907, n34908, n34909, n34910, n34911, n34912, n34913, n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921, n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929, n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937, n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945, n34946, n34947, n34948, n34949, n34950, n34951, n34952, n34953, n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961, n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969, n34970, n34971, n34972, n34973, n34974, n34975, n34976, n34977, n34978, n34979, n34980, n34981, n34982, n34983, n34984, n34985, n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993, n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001, n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009, n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017, n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35025, n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033, n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041, n35042, n35043, n35044, n35045, n35046, n35047, n35048, n35049, n35050, n35051, n35052, n35053, n35054, n35055, n35056, n35057, n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065, n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073, n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081, n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089, n35090, n35091, n35092, n35093, n35094, n35095, n35096, n35097, n35098, n35099, n35100, n35101, n35102, n35103, n35104, n35105, n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113, n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121, n35122, n35123, n35124, n35125, n35126, n35127, n35128, n35129, n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137, n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145, n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153, n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161, n35162, n35163, n35164, n35165, n35166, n35167, n35168, n35169, n35170, n35171, n35172, n35173, n35174, n35175, n35176, n35177, n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185, n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35193, n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201, n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209, n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217, n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225, n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233, n35234, n35235, n35236, n35237, n35238, n35239, n35240, n35241, n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249, n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257, n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265, n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273, n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281, n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289, n35290, n35291, n35292, n35293, n35294, n35295, n35296, n35297, n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305, n35306, n35307, n35308, n35309, n35310, n35311, n35312, n35313, n35314, n35315, n35316, n35317, n35318, n35319, n35320, n35321, n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329, n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337, n35338, n35339, n35340, n35341, n35342, n35343, n35344, n35345, n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353, n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361, n35362, n35363, n35364, n35365, n35366, n35367, n35368, n35369, n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377, n35378, n35379, n35380, n35381, n35382, n35383, n35384, n35385, n35386, n35387, n35388, n35389, n35390, n35391, n35392, n35393, n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401, n35402, n35403, n35404, n35405, n35406, n35407, n35408, n35409, n35410, n35411, n35412, n35413, n35414, n35415, n35416, n35417, n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425, n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433, n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441, n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449, n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457, n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465, n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473, n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481, n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489, n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497, n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505, n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513, n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521, n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529, n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537, n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545, n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553, n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561, n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569, n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577, n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585, n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593, n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601, n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609, n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617, n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625, n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633, n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641, n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649, n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657, n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665, n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673, n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681, n35682, n35683, n35684, n35685, n35686, n35687, n35688, n35689, n35690, n35691, n35692, n35693, n35694, n35695, n35696, n35697, n35698, n35699, n35700, n35701, n35702, n35703, n35704, n35705, n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713, n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721, n35722, n35723, n35724, n35725, n35726, n35727, n35728, n35729, n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737, n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745, n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753, n35754, n35755, n35756, n35757, n35758, n35759, n35760, n35761, n35762, n35763, n35764, n35765, n35766, n35767, n35768, n35769, n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777, n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785, n35786, n35787, n35788, n35789, n35790, n35791, n35792, n35793, n35794, n35795, n35796, n35797, n35798, n35799, n35800, n35801, n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809, n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35817, n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825, n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833, n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841, n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849, n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857, n35858, n35859, n35860, n35861, n35862, n35863, n35864, n35865, n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873, n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881, n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889, n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897, n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905, n35906, n35907, n35908, n35909, n35910, n35911, n35912, n35913, n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921, n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929, n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937, n35938, n35939, n35940, n35941, n35942, n35943, n35944, n35945, n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953, n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961, n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969, n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977, n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985, n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993, n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001, n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009, n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017, n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025, n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033, n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041, n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049, n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057, n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065, n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073, n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081, n36082, n36083, n36084, n36085, n36086, n36087, n36088, n36089, n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097, n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105, n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113, n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121, n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129, n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137, n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145, n36146, n36147, n36148, n36149, n36150, n36151, n36152, n36153, n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161, n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169, n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177, n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185, n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193, n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201, n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209, n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217, n36218, n36219, n36220, n36221, n36222, n36223, n36224, n36225, n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233, n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241, n36242, n36243, n36244, n36245, n36246, n36247, n36248, n36249, n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257, n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265, n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273, n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281, n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289, n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297, n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305, n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313, n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321, n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329, n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337, n36338, n36339, n36340, n36341, n36342, n36343, n36344, n36345, n36346, n36347, n36348, n36349, n36350, n36351, n36352, n36353, n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361, n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369, n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377, n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385, n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393, n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401, n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409, n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417, n36418, n36419, n36420, n36421, n36422, n36423, n36424, n36425, n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433, n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441, n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449, n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457, n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465, n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473, n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481, n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489, n36490, n36491, n36492, n36493, n36494, n36495, n36496, n36497, n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505, n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513, n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521, n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529, n36530, n36531, n36532, n36533, n36534, n36535, n36536, n36537, n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545, n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553, n36554, n36555, n36556, n36557, n36558, n36559, n36560, n36561, n36562, n36563, n36564, n36565, n36566, n36567, n36568, n36569, n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577, n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585, n36586, n36587, n36588, n36589, n36590, n36591, n36592, n36593, n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601, n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609, n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617, n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625, n36626, n36627, n36628, n36629, n36630, n36631, n36632, n36633, n36634, n36635, n36636, n36637, n36638, n36639, n36640, n36641, n36642, n36643, n36644, n36645, n36646, n36647, n36648, n36649, n36650, n36651, n36652, n36653, n36654, n36655, n36656, n36657, n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665, n36666, n36667, n36668, n36669, n36670, n36671, n36672, n36673, n36674, n36675, n36676, n36677, n36678, n36679, n36680, n36681, n36682, n36683, n36684, n36685, n36686, n36687, n36688, n36689, n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697, n36698, n36699, n36700, n36701, n36702, n36703, n36704, n36705, n36706, n36707, n36708, n36709, n36710, n36711, n36712, n36713, n36714, n36715, n36716, n36717, n36718, n36719, n36720, n36721, n36722, n36723, n36724, n36725, n36726, n36727, n36728, n36729, n36730, n36731, n36732, n36733, n36734, n36735, n36736, n36737, n36738, n36739, n36740, n36741, n36742, n36743, n36744, n36745, n36746, n36747, n36748, n36749, n36750, n36751, n36752, n36753, n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761, n36762, n36763, n36764, n36765, n36766, n36767, n36768, n36769, n36770, n36771, n36772, n36773, n36774, n36775, n36776, n36777, n36778, n36779, n36780, n36781, n36782, n36783, n36784, n36785, n36786, n36787, n36788, n36789, n36790, n36791, n36792, n36793, n36794, n36795, n36796, n36797, n36798, n36799, n36800, n36801, n36802, n36803, n36804, n36805, n36806, n36807, n36808, n36809, n36810, n36811, n36812, n36813, n36814, n36815, n36816, n36817, n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825, n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833, n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841, n36842, n36843, n36844, n36845, n36846, n36847, n36848, n36849, n36850, n36851, n36852, n36853, n36854, n36855, n36856, n36857, n36858, n36859, n36860, n36861, n36862, n36863, n36864, n36865, n36866, n36867, n36868, n36869, n36870, n36871, n36872, n36873, n36874, n36875, n36876, n36877, n36878, n36879, n36880, n36881, n36882, n36883, n36884, n36885, n36886, n36887, n36888, n36889, n36890, n36891, n36892, n36893, n36894, n36895, n36896, n36897, n36898, n36899, n36900, n36901, n36902, n36903, n36904, n36905, n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913, n36914, n36915, n36916, n36917, n36918, n36919, n36920, n36921, n36922, n36923, n36924, n36925, n36926, n36927, n36928, n36929, n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937, n36938, n36939, n36940, n36941, n36942, n36943, n36944, n36945, n36946, n36947, n36948, n36949, n36950, n36951, n36952, n36953, n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961, n36962, n36963, n36964, n36965, n36966, n36967, n36968, n36969, n36970, n36971, n36972, n36973, n36974, n36975, n36976, n36977, n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985, n36986, n36987, n36988, n36989, n36990, n36991, n36992, n36993, n36994, n36995, n36996, n36997, n36998, n36999, n37000, n37001, n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009, n37010, n37011, n37012, n37013, n37014, n37015, n37016, n37017, n37018, n37019, n37020, n37021, n37022, n37023, n37024, n37025, n37026, n37027, n37028, n37029, n37030, n37031, n37032, n37033, n37034, n37035, n37036, n37037, n37038, n37039, n37040, n37041, n37042, n37043, n37044, n37045, n37046, n37047, n37048, n37049, n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057, n37058, n37059, n37060, n37061, n37062, n37063, n37064, n37065, n37066, n37067, n37068, n37069, n37070, n37071, n37072, n37073, n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081, n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089, n37090, n37091, n37092, n37093, n37094, n37095, n37096, n37097, n37098, n37099, n37100, n37101, n37102, n37103, n37104, n37105, n37106, n37107, n37108, n37109, n37110, n37111, n37112, n37113, n37114, n37115, n37116, n37117, n37118, n37119, n37120, n37121, n37122, n37123, n37124, n37125, n37126, n37127, n37128, n37129, n37130, n37131, n37132, n37133, n37134, n37135, n37136, n37137, n37138, n37139, n37140, n37141, n37142, n37143, n37144, n37145, n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153, n37154, n37155, n37156, n37157, n37158, n37159, n37160, n37161, n37162, n37163, n37164, n37165, n37166, n37167, n37168, n37169, n37170, n37171, n37172, n37173, n37174, n37175, n37176, n37177, n37178, n37179, n37180, n37181, n37182, n37183, n37184, n37185, n37186, n37187, n37188, n37189, n37190, n37191, n37192, n37193, n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201, n37202, n37203, n37204, n37205, n37206, n37207, n37208, n37209, n37210, n37211, n37212, n37213, n37214, n37215, n37216, n37217, n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225, n37226, n37227, n37228, n37229, n37230, n37231, n37232, n37233, n37234, n37235, n37236, n37237, n37238, n37239, n37240, n37241, n37242, n37243, n37244, n37245, n37246, n37247, n37248, n37249, n37250, n37251, n37252, n37253, n37254, n37255, n37256, n37257, n37258, n37259, n37260, n37261, n37262, n37263, n37264, n37265, n37266, n37267, n37268, n37269, n37270, n37271, n37272, n37273, n37274, n37275, n37276, n37277, n37278, n37279, n37280, n37281, n37282, n37283, n37284, n37285, n37286, n37287, n37288, n37289, n37290, n37291, n37292, n37293, n37294, n37295, n37296, n37297, n37298, n37299, n37300, n37301, n37302, n37303, n37304, n37305, n37306, n37307, n37308, n37309, n37310, n37311, n37312, n37313, n37314, n37315, n37316, n37317, n37318, n37319, n37320, n37321, n37322, n37323, n37324, n37325, n37326, n37327, n37328, n37329, n37330, n37331, n37332, n37333, n37334, n37335, n37336, n37337, n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345, n37346, n37347, n37348, n37349, n37350, n37351, n37352, n37353, n37354, n37355, n37356, n37357, n37358, n37359, n37360, n37361, n37362, n37363, n37364, n37365, n37366, n37367, n37368, n37369, n37370, n37371, n37372, n37373, n37374, n37375, n37376, n37377, n37378, n37379, n37380, n37381, n37382, n37383, n37384, n37385, n37386, n37387, n37388, n37389, n37390, n37391, n37392, n37393, n37394, n37395, n37396, n37397, n37398, n37399, n37400, n37401, n37402, n37403, n37404, n37405, n37406, n37407, n37408, n37409, n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417, n37418, n37419, n37420, n37421, n37422, n37423, n37424, n37425, n37426, n37427, n37428, n37429, n37430, n37431, n37432, n37433, n37434, n37435, n37436, n37437, n37438, n37439, n37440, n37441, n37442, n37443, n37444, n37445, n37446, n37447, n37448, n37449, n37450, n37451, n37452, n37453, n37454, n37455, n37456, n37457, n37458, n37459, n37460, n37461, n37462, n37463, n37464, n37465, n37466, n37467, n37468, n37469, n37470, n37471, n37472, n37473, n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481, n37482, n37483, n37484, n37485, n37486, n37487, n37488, n37489, n37490, n37491, n37492, n37493, n37494, n37495, n37496, n37497, n37498, n37499, n37500, n37501, n37502, n37503, n37504, n37505, n37506, n37507, n37508, n37509, n37510, n37511, n37512, n37513, n37514, n37515, n37516, n37517, n37518, n37519, n37520, n37521, n37522, n37523, n37524, n37525, n37526, n37527, n37528, n37529, n37530, n37531, n37532, n37533, n37534, n37535, n37536, n37537, n37538, n37539, n37540, n37541, n37542, n37543, n37544, n37545, n37546, n37547, n37548, n37549, n37550, n37551, n37552, n37553, n37554, n37555, n37556, n37557, n37558, n37559, n37560, n37561, n37562, n37563, n37564, n37565, n37566, n37567, n37568, n37569, n37570, n37571, n37572, n37573, n37574, n37575, n37576, n37577, n37578, n37579, n37580, n37581, n37582, n37583, n37584, n37585, n37586, n37587, n37588, n37589, n37590, n37591, n37592, n37593, n37594, n37595, n37596, n37597, n37598, n37599, n37600, n37601, n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609, n37610, n37611, n37612, n37613, n37614, n37615, n37616, n37617, n37618, n37619, n37620, n37621, n37622, n37623, n37624, n37625, n37626, n37627, n37628, n37629, n37630, n37631, n37632, n37633, n37634, n37635, n37636, n37637, n37638, n37639, n37640, n37641, n37642, n37643, n37644, n37645, n37646, n37647, n37648, n37649, n37650, n37651, n37652, n37653, n37654, n37655, n37656, n37657, n37658, n37659, n37660, n37661, n37662, n37663, n37664, n37665, n37666, n37667, n37668, n37669, n37670, n37671, n37672, n37673, n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681, n37682, n37683, n37684, n37685, n37686, n37687, n37688, n37689, n37690, n37691, n37692, n37693, n37694, n37695, n37696, n37697, n37698, n37699, n37700, n37701, n37702, n37703, n37704, n37705, n37706, n37707, n37708, n37709, n37710, n37711, n37712, n37713, n37714, n37715, n37716, n37717, n37718, n37719, n37720, n37721, n37722, n37723, n37724, n37725, n37726, n37727, n37728, n37729, n37730, n37731, n37732, n37733, n37734, n37735, n37736, n37737, n37738, n37739, n37740, n37741, n37742, n37743, n37744, n37745, n37746, n37747, n37748, n37749, n37750, n37751, n37752, n37753, n37754, n37755, n37756, n37757, n37758, n37759, n37760, n37761, n37762, n37763, n37764, n37765, n37766, n37767, n37768, n37769, n37770, n37771, n37772, n37773, n37774, n37775, n37776, n37777, n37778, n37779, n37780, n37781, n37782, n37783, n37784, n37785, n37786, n37787, n37788, n37789, n37790, n37791, n37792, n37793, n37794, n37795, n37796, n37797, n37798, n37799, n37800, n37801, n37802, n37803, n37804, n37805, n37806, n37807, n37808, n37809, n37810, n37811, n37812, n37813, n37814, n37815, n37816, n37817, n37818, n37819, n37820, n37821, n37822, n37823, n37824, n37825, n37826, n37827, n37828, n37829, n37830, n37831, n37832, n37833, n37834, n37835, n37836, n37837, n37838, n37839, n37840, n37841, n37842, n37843, n37844, n37845, n37846, n37847, n37848, n37849, n37850, n37851, n37852, n37853, n37854, n37855, n37856, n37857, n37858, n37859, n37860, n37861, n37862, n37863, n37864, n37865, n37866, n37867, n37868, n37869, n37870, n37871, n37872, n37873, n37874, n37875, n37876, n37877, n37878, n37879, n37880, n37881, n37882, n37883, n37884, n37885, n37886, n37887, n37888, n37889, n37890, n37891, n37892, n37893, n37894, n37895, n37896, n37897, n37898, n37899, n37900, n37901, n37902, n37903, n37904, n37905, n37906, n37907, n37908, n37909, n37910, n37911, n37912, n37913, n37914, n37915, n37916, n37917, n37918, n37919, n37920, n37921, n37922, n37923, n37924, n37925, n37926, n37927, n37928, n37929, n37930, n37931, n37932, n37933, n37934, n37935, n37936, n37937, n37938, n37939, n37940, n37941, n37942, n37943, n37944, n37945, n37946, n37947, n37948, n37949, n37950, n37951, n37952, n37953, n37954, n37955, n37956, n37957, n37958, n37959, n37960, n37961, n37962, n37963, n37964, n37965, n37966, n37967, n37968, n37969, n37970, n37971, n37972, n37973, n37974, n37975, n37976, n37977, n37978, n37979, n37980, n37981, n37982, n37983, n37984, n37985, n37986, n37987, n37988, n37989, n37990, n37991, n37992, n37993, n37994, n37995, n37996, n37997, n37998, n37999, n38000, n38001, n38002, n38003, n38004, n38005, n38006, n38007, n38008, n38009, n38010, n38011, n38012, n38013, n38014, n38015, n38016, n38017, n38018, n38019, n38020, n38021, n38022, n38023, n38024, n38025, n38026, n38027, n38028, n38029, n38030, n38031, n38032, n38033, n38034, n38035, n38036, n38037, n38038, n38039, n38040, n38041, n38042, n38043, n38044, n38045, n38046, n38047, n38048, n38049, n38050, n38051, n38052, n38053, n38054, n38055, n38056, n38057, n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065, n38066, n38067, n38068, n38069, n38070, n38071, n38072, n38073, n38074, n38075, n38076, n38077, n38078, n38079, n38080, n38081, n38082, n38083, n38084, n38085, n38086, n38087, n38088, n38089, n38090, n38091, n38092, n38093, n38094, n38095, n38096, n38097, n38098, n38099, n38100, n38101, n38102, n38103, n38104, n38105, n38106, n38107, n38108, n38109, n38110, n38111, n38112, n38113, n38114, n38115, n38116, n38117, n38118, n38119, n38120, n38121, n38122, n38123, n38124, n38125, n38126, n38127, n38128, n38129, n38130, n38131, n38132, n38133, n38134, n38135, n38136, n38137, n38138, n38139, n38140, n38141, n38142, n38143, n38144, n38145, n38146, n38147, n38148, n38149, n38150, n38151, n38152, n38153, n38154, n38155, n38156, n38157, n38158, n38159, n38160, n38161, n38162, n38163, n38164, n38165, n38166, n38167, n38168, n38169, n38170, n38171, n38172, n38173, n38174, n38175, n38176, n38177, n38178, n38179, n38180, n38181, n38182, n38183, n38184, n38185, n38186, n38187, n38188, n38189, n38190, n38191, n38192, n38193, n38194, n38195, n38196, n38197, n38198, n38199, n38200, n38201, n38202, n38203, n38204, n38205, n38206, n38207, n38208, n38209, n38210, n38211, n38212, n38213, n38214, n38215, n38216, n38217, n38218, n38219, n38220, n38221, n38222, n38223, n38224, n38225, n38226, n38227, n38228, n38229, n38230, n38231, n38232, n38233, n38234, n38235, n38236, n38237, n38238, n38239, n38240, n38241, n38242, n38243, n38244, n38245, n38246, n38247, n38248, n38249, n38250, n38251, n38252, n38253, n38254, n38255, n38256, n38257, n38258, n38259, n38260, n38261, n38262, n38263, n38264, n38265, n38266, n38267, n38268, n38269, n38270, n38271, n38272, n38273, n38274, n38275, n38276, n38277, n38278, n38279, n38280, n38281, n38282, n38283, n38284, n38285, n38286, n38287, n38288, n38289, n38290, n38291, n38292, n38293, n38294, n38295, n38296, n38297, n38298, n38299, n38300, n38301, n38302, n38303, n38304, n38305, n38306, n38307, n38308, n38309, n38310, n38311, n38312, n38313, n38314, n38315, n38316, n38317, n38318, n38319, n38320, n38321, n38322, n38323, n38324, n38325, n38326, n38327, n38328, n38329, n38330, n38331, n38332, n38333, n38334, n38335, n38336, n38337, n38338, n38339, n38340, n38341, n38342, n38343, n38344, n38345, n38346, n38347, n38348, n38349, n38350, n38351, n38352, n38353, n38354, n38355, n38356, n38357, n38358, n38359, n38360, n38361, n38362, n38363, n38364, n38365, n38366, n38367, n38368, n38369, n38370, n38371, n38372, n38373, n38374, n38375, n38376, n38377, n38378, n38379, n38380, n38381, n38382, n38383, n38384, n38385, n38386, n38387, n38388, n38389, n38390, n38391, n38392, n38393, n38394, n38395, n38396, n38397, n38398, n38399, n38400, n38401, n38402, n38403, n38404, n38405, n38406, n38407, n38408, n38409, n38410, n38411, n38412, n38413, n38414, n38415, n38416, n38417, n38418, n38419, n38420, n38421, n38422, n38423, n38424, n38425, n38426, n38427, n38428, n38429, n38430, n38431, n38432, n38433, n38434, n38435, n38436, n38437, n38438, n38439, n38440, n38441, n38442, n38443, n38444, n38445, n38446, n38447, n38448, n38449, n38450, n38451, n38452, n38453, n38454, n38455, n38456, n38457, n38458, n38459, n38460, n38461, n38462, n38463, n38464, n38465, n38466, n38467, n38468, n38469, n38470, n38471, n38472, n38473, n38474, n38475, n38476, n38477, n38478, n38479, n38480, n38481, n38482, n38483, n38484, n38485, n38486, n38487, n38488, n38489, n38490, n38491, n38492, n38493, n38494, n38495, n38496, n38497, n38498, n38499, n38500, n38501, n38502, n38503, n38504, n38505, n38506, n38507, n38508, n38509, n38510, n38511, n38512, n38513, n38514, n38515, n38516, n38517, n38518, n38519, n38520, n38521, n38522, n38523, n38524, n38525, n38526, n38527, n38528, n38529, n38530, n38531, n38532, n38533, n38534, n38535, n38536, n38537, n38538, n38539, n38540, n38541, n38542, n38543, n38544, n38545, n38546, n38547, n38548, n38549, n38550, n38551, n38552, n38553, n38554, n38555, n38556, n38557, n38558, n38559, n38560, n38561, n38562, n38563, n38564, n38565, n38566, n38567, n38568, n38569, n38570, n38571, n38572, n38573, n38574, n38575, n38576, n38577, n38578, n38579, n38580, n38581, n38582, n38583, n38584, n38585, n38586, n38587, n38588, n38589, n38590, n38591, n38592, n38593, n38594, n38595, n38596, n38597, n38598, n38599, n38600, n38601, n38602, n38603, n38604, n38605, n38606, n38607, n38608, n38609, n38610, n38611, n38612, n38613, n38614, n38615, n38616, n38617, n38618, n38619, n38620, n38621, n38622, n38623, n38624, n38625, n38626, n38627, n38628, n38629, n38630, n38631, n38632, n38633, n38634, n38635, n38636, n38637, n38638, n38639, n38640, n38641, n38642, n38643, n38644, n38645, n38646, n38647, n38648, n38649, n38650, n38651, n38652, n38653, n38654, n38655, n38656, n38657, n38658, n38659, n38660, n38661, n38662, n38663, n38664, n38665, n38666, n38667, n38668, n38669, n38670, n38671, n38672, n38673, n38674, n38675, n38676, n38677, n38678, n38679, n38680, n38681, n38682, n38683, n38684, n38685, n38686, n38687, n38688, n38689, n38690, n38691, n38692, n38693, n38694, n38695, n38696, n38697, n38698, n38699, n38700, n38701, n38702, n38703, n38704, n38705, n38706, n38707, n38708, n38709, n38710, n38711, n38712, n38713, n38714, n38715, n38716, n38717, n38718, n38719, n38720, n38721, n38722, n38723, n38724, n38725, n38726, n38727, n38728, n38729, n38730, n38731, n38732, n38733, n38734, n38735, n38736, n38737, n38738, n38739, n38740, n38741, n38742, n38743, n38744, n38745, n38746, n38747, n38748, n38749, n38750, n38751, n38752, n38753, n38754, n38755, n38756, n38757, n38758, n38759, n38760, n38761, n38762, n38763, n38764, n38765, n38766, n38767, n38768, n38769, n38770, n38771, n38772, n38773, n38774, n38775, n38776, n38777, n38778, n38779, n38780, n38781, n38782, n38783, n38784, n38785, n38786, n38787, n38788, n38789, n38790, n38791, n38792, n38793, n38794, n38795, n38796, n38797, n38798, n38799, n38800, n38801, n38802, n38803, n38804, n38805, n38806, n38807, n38808, n38809, n38810, n38811, n38812, n38813, n38814, n38815, n38816, n38817, n38818, n38819, n38820, n38821, n38822, n38823, n38824, n38825, n38826, n38827, n38828, n38829, n38830, n38831, n38832, n38833, n38834, n38835, n38836, n38837, n38838, n38839, n38840, n38841, n38842, n38843, n38844, n38845, n38846, n38847, n38848, n38849, n38850, n38851, n38852, n38853, n38854, n38855, n38856, n38857, n38858, n38859, n38860, n38861, n38862, n38863, n38864, n38865, n38866, n38867, n38868, n38869, n38870, n38871, n38872, n38873, n38874, n38875, n38876, n38877, n38878, n38879, n38880, n38881, n38882, n38883, n38884, n38885, n38886, n38887, n38888, n38889, n38890, n38891, n38892, n38893, n38894, n38895, n38896, n38897, n38898, n38899, n38900, n38901, n38902, n38903, n38904, n38905, n38906, n38907, n38908, n38909, n38910, n38911, n38912, n38913, n38914, n38915, n38916, n38917, n38918, n38919, n38920, n38921, n38922, n38923, n38924, n38925, n38926, n38927, n38928, n38929, n38930, n38931, n38932, n38933, n38934, n38935, n38936, n38937, n38938, n38939, n38940, n38941, n38942, n38943, n38944, n38945, n38946, n38947, n38948, n38949, n38950, n38951, n38952, n38953, n38954, n38955, n38956, n38957, n38958, n38959, n38960, n38961, n38962, n38963, n38964, n38965, n38966, n38967, n38968, n38969, n38970, n38971, n38972, n38973, n38974, n38975, n38976, n38977, n38978, n38979, n38980, n38981, n38982, n38983, n38984, n38985, n38986, n38987, n38988, n38989, n38990, n38991, n38992, n38993, n38994, n38995, n38996, n38997, n38998, n38999, n39000, n39001, n39002, n39003, n39004, n39005, n39006, n39007, n39008, n39009, n39010, n39011, n39012, n39013, n39014, n39015, n39016, n39017, n39018, n39019, n39020, n39021, n39022, n39023, n39024, n39025, n39026, n39027, n39028, n39029, n39030, n39031, n39032, n39033, n39034, n39035, n39036, n39037, n39038, n39039, n39040, n39041, n39042, n39043, n39044, n39045, n39046, n39047, n39048, n39049, n39050, n39051, n39052, n39053, n39054, n39055, n39056, n39057, n39058, n39059, n39060, n39061, n39062, n39063, n39064, n39065, n39066, n39067, n39068, n39069, n39070, n39071, n39072, n39073, n39074, n39075, n39076, n39077, n39078, n39079, n39080, n39081, n39082, n39083, n39084, n39085, n39086, n39087, n39088, n39089, n39090, n39091, n39092, n39093, n39094, n39095, n39096, n39097, n39098, n39099, n39100, n39101, n39102, n39103, n39104, n39105, n39106, n39107, n39108, n39109, n39110, n39111, n39112, n39113, n39114, n39115, n39116, n39117, n39118, n39119, n39120, n39121, n39122, n39123, n39124, n39125, n39126, n39127, n39128, n39129, n39130, n39131, n39132, n39133, n39134, n39135, n39136, n39137, n39138, n39139, n39140, n39141, n39142, n39143, n39144, n39145, n39146, n39147, n39148, n39149, n39150, n39151, n39152, n39153, n39154, n39155, n39156, n39157, n39158, n39159, n39160, n39161, n39162, n39163, n39164, n39165, n39166, n39167, n39168, n39169, n39170, n39171, n39172, n39173, n39174, n39175, n39176, n39177, n39178, n39179, n39180, n39181, n39182, n39183, n39184, n39185, n39186, n39187, n39188, n39189, n39190, n39191, n39192, n39193, n39194, n39195, n39196, n39197, n39198, n39199, n39200, n39201, n39202, n39203, n39204, n39205, n39206, n39207, n39208, n39209, n39210, n39211, n39212, n39213, n39214, n39215, n39216, n39217, n39218, n39219, n39220, n39221, n39222, n39223, n39224, n39225, n39226, n39227, n39228, n39229, n39230, n39231, n39232, n39233, n39234, n39235, n39236, n39237, n39238, n39239, n39240, n39241, n39242, n39243, n39244, n39245, n39246, n39247, n39248, n39249, n39250, n39251, n39252, n39253, n39254, n39255, n39256, n39257, n39258, n39259, n39260, n39261, n39262, n39263, n39264, n39265, n39266, n39267, n39268, n39269, n39270, n39271, n39272, n39273, n39274, n39275, n39276, n39277, n39278, n39279, n39280, n39281, n39282, n39283, n39284, n39285, n39286, n39287, n39288, n39289, n39290, n39291, n39292, n39293, n39294, n39295, n39296, n39297, n39298, n39299, n39300, n39301, n39302, n39303, n39304, n39305, n39306, n39307, n39308, n39309, n39310, n39311, n39312, n39313, n39314, n39315, n39316, n39317, n39318, n39319, n39320, n39321, n39322, n39323, n39324, n39325, n39326, n39327, n39328, n39329, n39330, n39331, n39332, n39333, n39334, n39335, n39336, n39337, n39338, n39339, n39340, n39341, n39342, n39343, n39344, n39345, n39346, n39347, n39348, n39349, n39350, n39351, n39352, n39353, n39354, n39355, n39356, n39357, n39358, n39359, n39360, n39361, n39362, n39363, n39364, n39365, n39366, n39367, n39368, n39369, n39370, n39371, n39372, n39373, n39374, n39375, n39376, n39377, n39378, n39379, n39380, n39381, n39382, n39383, n39384, n39385, n39386, n39387, n39388, n39389, n39390, n39391, n39392, n39393, n39394, n39395, n39396, n39397, n39398, n39399, n39400, n39401, n39402, n39403, n39404, n39405, n39406, n39407, n39408, n39409, n39410, n39411, n39412, n39413, n39414, n39415, n39416, n39417, n39418, n39419, n39420, n39421, n39422, n39423, n39424, n39425, n39426, n39427, n39428, n39429, n39430, n39431, n39432, n39433, n39434, n39435, n39436, n39437, n39438, n39439, n39440, n39441, n39442, n39443, n39444, n39445, n39446, n39447, n39448, n39449, n39450, n39451, n39452, n39453, n39454, n39455, n39456, n39457, n39458, n39459, n39460, n39461, n39462, n39463, n39464, n39465, n39466, n39467, n39468, n39469, n39470, n39471, n39472, n39473, n39474, n39475, n39476, n39477, n39478, n39479, n39480, n39481, n39482, n39483, n39484, n39485, n39486, n39487, n39488, n39489, n39490, n39491, n39492, n39493, n39494, n39495, n39496, n39497, n39498, n39499, n39500, n39501, n39502, n39503, n39504, n39505, n39506, n39507, n39508, n39509, n39510, n39511, n39512, n39513, n39514, n39515, n39516, n39517, n39518, n39519, n39520, n39521, n39522, n39523, n39524, n39525, n39526, n39527, n39528, n39529, n39530, n39531, n39532, n39533, n39534, n39535, n39536, n39537, n39538, n39539, n39540, n39541, n39542, n39543, n39544, n39545, n39546, n39547, n39548, n39549, n39550, n39551, n39552, n39553, n39554, n39555, n39556, n39557, n39558, n39559, n39560, n39561, n39562, n39563, n39564, n39565, n39566, n39567, n39568, n39569, n39570, n39571, n39572, n39573, n39574, n39575, n39576, n39577, n39578, n39579, n39580, n39581, n39582, n39583, n39584, n39585, n39586, n39587, n39588, n39589, n39590, n39591, n39592, n39593, n39594, n39595, n39596, n39597, n39598, n39599, n39600, n39601, n39602, n39603, n39604, n39605, n39606, n39607, n39608, n39609, n39610, n39611, n39612, n39613, n39614, n39615, n39616, n39617, n39618, n39619, n39620, n39621, n39622, n39623, n39624, n39625, n39626, n39627, n39628, n39629, n39630, n39631, n39632, n39633, n39634, n39635, n39636, n39637, n39638, n39639, n39640, n39641, n39642, n39643, n39644, n39645, n39646, n39647, n39648, n39649, n39650, n39651, n39652, n39653, n39654, n39655, n39656, n39657, n39658, n39659, n39660, n39661, n39662, n39663, n39664, n39665, n39666, n39667, n39668, n39669, n39670, n39671, n39672, n39673, n39674, n39675, n39676, n39677, n39678, n39679, n39680, n39681, n39682, n39683, n39684, n39685, n39686, n39687, n39688, n39689, n39690, n39691, n39692, n39693, n39694, n39695, n39696, n39697, n39698, n39699, n39700, n39701, n39702, n39703, n39704, n39705, n39706, n39707, n39708, n39709, n39710, n39711, n39712, n39713, n39714, n39715, n39716, n39717, n39718, n39719, n39720, n39721, n39722, n39723, n39724, n39725, n39726, n39727, n39728, n39729, n39730, n39731, n39732, n39733, n39734, n39735, n39736, n39737, n39738, n39739, n39740, n39741, n39742, n39743, n39744, n39745, n39746, n39747, n39748, n39749, n39750, n39751, n39752, n39753, n39754, n39755, n39756, n39757, n39758, n39759, n39760, n39761, n39762, n39763, n39764, n39765, n39766, n39767, n39768, n39769, n39770, n39771, n39772, n39773, n39774, n39775, n39776, n39777, n39778, n39779, n39780, n39781, n39782, n39783, n39784, n39785, n39786, n39787, n39788, n39789, n39790, n39791, n39792, n39793, n39794, n39795, n39796, n39797, n39798, n39799, n39800, n39801, n39802, n39803, n39804, n39805, n39806, n39807, n39808, n39809, n39810, n39811, n39812, n39813, n39814, n39815, n39816, n39817, n39818, n39819, n39820, n39821, n39822, n39823, n39824, n39825, n39826, n39827, n39828, n39829, n39830, n39831, n39832, n39833, n39834, n39835, n39836, n39837, n39838, n39839, n39840, n39841, n39842, n39843, n39844, n39845, n39846, n39847, n39848, n39849, n39850, n39851, n39852, n39853, n39854, n39855, n39856, n39857, n39858, n39859, n39860, n39861, n39862, n39863, n39864, n39865, n39866, n39867, n39868, n39869, n39870, n39871, n39872, n39873, n39874, n39875, n39876, n39877, n39878, n39879, n39880, n39881, n39882, n39883, n39884, n39885, n39886, n39887, n39888, n39889, n39890, n39891, n39892, n39893, n39894, n39895, n39896, n39897, n39898, n39899, n39900, n39901, n39902, n39903, n39904, n39905, n39906, n39907, n39908, n39909, n39910, n39911, n39912, n39913, n39914, n39915, n39916, n39917, n39918, n39919, n39920, n39921, n39922, n39923, n39924, n39925, n39926, n39927, n39928, n39929, n39930, n39931, n39932, n39933, n39934, n39935, n39936, n39937, n39938, n39939, n39940, n39941, n39942, n39943, n39944, n39945, n39946, n39947, n39948, n39949, n39950, n39951, n39952, n39953, n39954, n39955, n39956, n39957, n39958, n39959, n39960, n39961, n39962, n39963, n39964, n39965, n39966, n39967, n39968, n39969, n39970, n39971, n39972, n39973, n39974, n39975, n39976, n39977, n39978, n39979, n39980, n39981, n39982, n39983, n39984, n39985, n39986, n39987, n39988, n39989, n39990, n39991, n39992, n39993, n39994, n39995, n39996, n39997, n39998, n39999, n40000, n40001, n40002, n40003, n40004, n40005, n40006, n40007, n40008, n40009, n40010, n40011, n40012, n40013, n40014, n40015, n40016, n40017, n40018, n40019, n40020, n40021, n40022, n40023, n40024, n40025, n40026, n40027, n40028, n40029, n40030, n40031, n40032, n40033, n40034, n40035, n40036, n40037, n40038, n40039, n40040, n40041, n40042, n40043, n40044, n40045, n40046, n40047, n40048, n40049, n40050, n40051, n40052, n40053, n40054, n40055, n40056, n40057, n40058, n40059, n40060, n40061, n40062, n40063, n40064, n40065, n40066, n40067, n40068, n40069, n40070, n40071, n40072, n40073, n40074, n40075, n40076, n40077, n40078, n40079, n40080, n40081, n40082, n40083, n40084, n40085, n40086, n40087, n40088, n40089, n40090, n40091, n40092, n40093, n40094, n40095, n40096, n40097, n40098, n40099, n40100, n40101, n40102, n40103, n40104, n40105, n40106, n40107, n40108, n40109, n40110, n40111, n40112, n40113, n40114, n40115, n40116, n40117, n40118, n40119, n40120, n40121, n40122, n40123, n40124, n40125, n40126, n40127, n40128, n40129, n40130, n40131, n40132, n40133, n40134, n40135, n40136, n40137, n40138, n40139, n40140, n40141, n40142, n40143, n40144, n40145, n40146, n40147, n40148, n40149, n40150, n40151, n40152, n40153, n40154, n40155, n40156, n40157, n40158, n40159, n40160, n40161, n40162, n40163, n40164, n40165, n40166, n40167, n40168, n40169, n40170, n40171, n40172, n40173, n40174, n40175, n40176, n40177, n40178, n40179, n40180, n40181, n40182, n40183, n40184, n40185, n40186, n40187, n40188, n40189, n40190, n40191, n40192, n40193, n40194, n40195, n40196, n40197, n40198, n40199, n40200, n40201, n40202, n40203, n40204, n40205, n40206, n40207, n40208, n40209, n40210, n40211, n40212, n40213, n40214, n40215, n40216, n40217, n40218, n40219, n40220, n40221, n40222, n40223, n40224, n40225, n40226, n40227, n40228, n40229, n40230, n40231, n40232, n40233, n40234, n40235, n40236, n40237, n40238, n40239, n40240, n40241, n40242, n40243, n40244, n40245, n40246, n40247, n40248, n40249, n40250, n40251, n40252, n40253, n40254, n40255, n40256, n40257, n40258, n40259, n40260, n40261, n40262, n40263, n40264, n40265, n40266, n40267, n40268, n40269, n40270, n40271, n40272, n40273, n40274, n40275, n40276, n40277, n40278, n40279, n40280, n40281, n40282, n40283, n40284, n40285, n40286, n40287, n40288, n40289, n40290, n40291, n40292, n40293, n40294, n40295, n40296, n40297, n40298, n40299, n40300, n40301, n40302, n40303, n40304, n40305, n40306, n40307, n40308, n40309, n40310, n40311, n40312, n40313, n40314, n40315, n40316, n40317, n40318, n40319, n40320, n40321, n40322, n40323, n40324, n40325, n40326, n40327, n40328, n40329, n40330, n40331, n40332, n40333, n40334, n40335, n40336, n40337, n40338, n40339, n40340, n40341, n40342, n40343, n40344, n40345, n40346, n40347, n40348, n40349, n40350, n40351, n40352, n40353, n40354, n40355, n40356, n40357, n40358, n40359, n40360, n40361, n40362, n40363, n40364, n40365, n40366, n40367, n40368, n40369, n40370, n40371, n40372, n40373, n40374, n40375, n40376, n40377, n40378, n40379, n40380, n40381, n40382, n40383, n40384, n40385, n40386, n40387, n40388, n40389, n40390, n40391, n40392, n40393, n40394, n40395, n40396, n40397, n40398, n40399, n40400, n40401, n40402, n40403, n40404, n40405, n40406, n40407, n40408, n40409, n40410, n40411, n40412, n40413, n40414, n40415, n40416, n40417, n40418, n40419, n40420, n40421, n40422, n40423, n40424, n40425, n40426, n40427, n40428, n40429, n40430, n40431, n40432, n40433, n40434, n40435, n40436, n40437, n40438, n40439, n40440, n40441, n40442, n40443, n40444, n40445, n40446, n40447, n40448, n40449, n40450, n40451, n40452, n40453, n40454, n40455, n40456, n40457, n40458, n40459, n40460, n40461, n40462, n40463, n40464, n40465, n40466, n40467, n40468, n40469, n40470, n40471, n40472, n40473, n40474, n40475, n40476, n40477, n40478, n40479, n40480, n40481, n40482, n40483, n40484, n40485, n40486, n40487, n40488, n40489, n40490, n40491, n40492, n40493, n40494, n40495, n40496, n40497, n40498, n40499, n40500, n40501, n40502, n40503, n40504, n40505, n40506, n40507, n40508, n40509, n40510, n40511, n40512, n40513, n40514, n40515, n40516, n40517, n40518, n40519, n40520, n40521, n40522, n40523, n40524, n40525, n40526, n40527, n40528, n40529, n40530, n40531, n40532, n40533, n40534, n40535, n40536, n40537, n40538, n40539, n40540, n40541, n40542, n40543, n40544, n40545, n40546, n40547, n40548, n40549, n40550, n40551, n40552, n40553, n40554, n40555, n40556, n40557, n40558, n40559, n40560, n40561, n40562, n40563, n40564, n40565, n40566, n40567, n40568, n40569, n40570, n40571, n40572, n40573, n40574, n40575, n40576, n40577, n40578, n40579, n40580, n40581, n40582, n40583, n40584, n40585, n40586, n40587, n40588, n40589, n40590, n40591, n40592, n40593, n40594, n40595, n40596, n40597, n40598, n40599, n40600, n40601, n40602, n40603, n40604, n40605, n40606, n40607, n40608, n40609, n40610, n40611, n40612, n40613, n40614, n40615, n40616, n40617, n40618, n40619, n40620, n40621, n40622, n40623, n40624, n40625, n40626, n40627, n40628, n40629, n40630, n40631, n40632, n40633, n40634, n40635, n40636, n40637, n40638, n40639, n40640, n40641, n40642, n40643, n40644, n40645, n40646, n40647, n40648, n40649, n40650, n40651, n40652, n40653, n40654, n40655, n40656, n40657, n40658, n40659, n40660, n40661, n40662, n40663, n40664, n40665, n40666, n40667, n40668, n40669, n40670, n40671, n40672, n40673, n40674, n40675, n40676, n40677, n40678, n40679, n40680, n40681, n40682, n40683, n40684, n40685, n40686, n40687, n40688, n40689, n40690, n40691, n40692, n40693, n40694, n40695, n40696, n40697, n40698, n40699, n40700, n40701, n40702, n40703, n40704, n40705, n40706, n40707, n40708, n40709, n40710, n40711, n40712, n40713, n40714, n40715, n40716, n40717, n40718, n40719, n40720, n40721, n40722, n40723, n40724, n40725, n40726, n40727, n40728, n40729, n40730, n40731, n40732, n40733, n40734, n40735, n40736, n40737, n40738, n40739, n40740, n40741, n40742, n40743, n40744, n40745, n40746, n40747, n40748, n40749, n40750, n40751, n40752, n40753, n40754, n40755, n40756, n40757, n40758, n40759, n40760, n40761, n40762, n40763, n40764, n40765, n40766, n40767, n40768, n40769, n40770, n40771, n40772, n40773, n40774, n40775, n40776, n40777, n40778, n40779, n40780, n40781, n40782, n40783, n40784, n40785, n40786, n40787, n40788, n40789, n40790, n40791, n40792, n40793, n40794, n40795, n40796, n40797, n40798, n40799, n40800, n40801, n40802, n40803, n40804, n40805, n40806, n40807, n40808, n40809, n40810, n40811, n40812, n40813, n40814, n40815, n40816, n40817, n40818, n40819, n40820, n40821, n40822, n40823, n40824, n40825, n40826, n40827, n40828, n40829, n40830, n40831, n40832, n40833, n40834, n40835, n40836, n40837, n40838, n40839, n40840, n40841, n40842, n40843, n40844, n40845, n40846, n40847, n40848, n40849, n40850, n40851, n40852, n40853, n40854, n40855, n40856, n40857, n40858, n40859, n40860, n40861, n40862, n40863, n40864, n40865, n40866, n40867, n40868, n40869, n40870, n40871, n40872, n40873, n40874, n40875, n40876, n40877, n40878, n40879, n40880, n40881, n40882, n40883, n40884, n40885, n40886, n40887, n40888, n40889, n40890, n40891, n40892, n40893, n40894, n40895, n40896, n40897, n40898, n40899, n40900, n40901, n40902, n40903, n40904, n40905, n40906, n40907, n40908, n40909, n40910, n40911, n40912, n40913, n40914, n40915, n40916, n40917, n40918, n40919, n40920, n40921, n40922, n40923, n40924, n40925, n40926, n40927, n40928, n40929, n40930, n40931, n40932, n40933, n40934, n40935, n40936, n40937, n40938, n40939, n40940, n40941, n40942, n40943, n40944, n40945, n40946, n40947, n40948, n40949, n40950, n40951, n40952, n40953, n40954, n40955, n40956, n40957, n40958, n40959, n40960, n40961, n40962, n40963, n40964, n40965, n40966, n40967, n40968, n40969, n40970, n40971, n40972, n40973, n40974, n40975, n40976, n40977, n40978, n40979, n40980, n40981, n40982, n40983, n40984, n40985, n40986, n40987, n40988, n40989, n40990, n40991, n40992, n40993, n40994, n40995, n40996, n40997, n40998, n40999, n41000, n41001, n41002, n41003, n41004, n41005, n41006, n41007, n41008, n41009, n41010, n41011, n41012, n41013, n41014, n41015, n41016, n41017, n41018, n41019, n41020, n41021, n41022, n41023, n41024, n41025, n41026, n41027, n41028, n41029, n41030, n41031, n41032, n41033, n41034, n41035, n41036, n41037, n41038, n41039, n41040, n41041, n41042, n41043, n41044, n41045, n41046, n41047, n41048, n41049, n41050, n41051, n41052, n41053, n41054, n41055, n41056, n41057, n41058, n41059, n41060, n41061, n41062, n41063, n41064, n41065, n41066, n41067, n41068, n41069, n41070, n41071, n41072, n41073, n41074, n41075, n41076, n41077, n41078, n41079, n41080, n41081, n41082, n41083, n41084, n41085, n41086, n41087, n41088, n41089, n41090, n41091, n41092, n41093, n41094, n41095, n41096, n41097, n41098, n41099, n41100, n41101, n41102, n41103, n41104, n41105, n41106, n41107, n41108, n41109, n41110, n41111, n41112, n41113, n41114, n41115, n41116, n41117, n41118, n41119, n41120, n41121, n41122, n41123, n41124, n41125, n41126, n41127, n41128, n41129, n41130, n41131, n41132, n41133, n41134, n41135, n41136, n41137, n41138, n41139, n41140, n41141, n41142, n41143, n41144, n41145, n41146, n41147, n41148, n41149, n41150, n41151, n41152, n41153, n41154, n41155, n41156, n41157, n41158, n41159, n41160, n41161, n41162, n41163, n41164, n41165, n41166, n41167, n41168, n41169, n41170, n41171, n41172, n41173, n41174, n41175, n41176, n41177, n41178, n41179, n41180, n41181, n41182, n41183, n41184, n41185, n41186, n41187, n41188, n41189, n41190, n41191, n41192, n41193, n41194, n41195, n41196, n41197, n41198, n41199, n41200, n41201, n41202, n41203, n41204, n41205, n41206, n41207, n41208, n41209, n41210, n41211, n41212, n41213, n41214, n41215, n41216, n41217, n41218, n41219, n41220, n41221, n41222, n41223, n41224, n41225, n41226, n41227, n41228, n41229, n41230, n41231, n41232, n41233, n41234, n41235, n41236, n41237, n41238, n41239, n41240, n41241, n41242, n41243, n41244, n41245, n41246, n41247, n41248, n41249, n41250, n41251, n41252, n41253, n41254, n41255, n41256, n41257, n41258, n41259, n41260, n41261, n41262, n41263, n41264, n41265, n41266, n41267, n41268, n41269, n41270, n41271, n41272, n41273, n41274, n41275, n41276, n41277, n41278, n41279, n41280, n41281, n41282, n41283, n41284, n41285, n41286, n41287, n41288, n41289, n41290, n41291, n41292, n41293, n41294, n41295, n41296, n41297, n41298, n41299, n41300, n41301, n41302, n41303, n41304, n41305, n41306, n41307, n41308, n41309, n41310, n41311, n41312, n41313, n41314, n41315, n41316, n41317, n41318, n41319, n41320, n41321, n41322, n41323, n41324, n41325, n41326, n41327, n41328, n41329, n41330, n41331, n41332, n41333, n41334, n41335, n41336, n41337, n41338, n41339, n41340, n41341, n41342, n41343, n41344, n41345, n41346, n41347, n41348, n41349, n41350, n41351, n41352, n41353, n41354, n41355, n41356, n41357, n41358, n41359, n41360, n41361, n41362, n41363, n41364, n41365, n41366, n41367, n41368, n41369, n41370, n41371, n41372, n41373, n41374, n41375, n41376, n41377, n41378, n41379, n41380, n41381, n41382, n41383, n41384, n41385, n41386, n41387, n41388, n41389, n41390, n41391, n41392, n41393, n41394, n41395, n41396, n41397, n41398, n41399, n41400, n41401, n41402, n41403, n41404, n41405, n41406, n41407, n41408, n41409, n41410, n41411, n41412, n41413, n41414, n41415, n41416, n41417, n41418, n41419, n41420, n41421, n41422, n41423, n41424, n41425, n41426, n41427, n41428, n41429, n41430, n41431, n41432, n41433, n41434, n41435, n41436, n41437, n41438, n41439, n41440, n41441, n41442, n41443, n41444, n41445, n41446, n41447, n41448, n41449, n41450, n41451, n41452, n41453, n41454, n41455, n41456, n41457, n41458, n41459, n41460, n41461, n41462, n41463, n41464, n41465, n41466, n41467, n41468, n41469, n41470, n41471, n41472, n41473, n41474, n41475, n41476, n41477, n41478, n41479, n41480, n41481, n41482, n41483, n41484, n41485, n41486, n41487, n41488, n41489, n41490, n41491, n41492, n41493, n41494, n41495, n41496, n41497, n41498, n41499, n41500, n41501, n41502, n41503, n41504, n41505, n41506, n41507, n41508, n41509, n41510, n41511, n41512, n41513, n41514, n41515, n41516, n41517, n41518, n41519, n41520, n41521, n41522, n41523, n41524, n41525, n41526, n41527, n41528, n41529, n41530, n41531, n41532, n41533, n41534, n41535, n41536, n41537, n41538, n41539, n41540, n41541, n41542, n41543, n41544, n41545, n41546, n41547, n41548, n41549, n41550, n41551, n41552, n41553, n41554, n41555, n41556, n41557, n41558, n41559, n41560, n41561, n41562, n41563, n41564, n41565, n41566, n41567, n41568, n41569, n41570, n41571, n41572, n41573, n41574, n41575, n41576, n41577, n41578, n41579, n41580, n41581, n41582, n41583, n41584, n41585, n41586, n41587, n41588, n41589, n41590, n41591, n41592, n41593, n41594, n41595, n41596, n41597, n41598, n41599, n41600, n41601, n41602, n41603, n41604, n41605, n41606, n41607, n41608, n41609, n41610, n41611, n41612, n41613, n41614, n41615, n41616, n41617, n41618, n41619, n41620, n41621, n41622, n41623, n41624, n41625, n41626, n41627, n41628, n41629, n41630, n41631, n41632, n41633, n41634, n41635, n41636, n41637, n41638, n41639, n41640, n41641, n41642, n41643, n41644, n41645, n41646, n41647, n41648, n41649, n41650, n41651, n41652, n41653, n41654, n41655, n41656, n41657, n41658, n41659, n41660, n41661, n41662, n41663, n41664, n41665, n41666, n41667, n41668, n41669, n41670, n41671, n41672, n41673, n41674, n41675, n41676, n41677, n41678, n41679, n41680, n41681, n41682, n41683, n41684, n41685, n41686, n41687, n41688, n41689, n41690, n41691, n41692, n41693, n41694, n41695, n41696, n41697, n41698, n41699, n41700, n41701, n41702, n41703, n41704, n41705, n41706, n41707, n41708, n41709, n41710, n41711, n41712, n41713, n41714, n41715, n41716, n41717, n41718, n41719, n41720, n41721, n41722, n41723, n41724, n41725, n41726, n41727, n41728, n41729, n41730, n41731, n41732, n41733, n41734, n41735, n41736, n41737, n41738, n41739, n41740, n41741, n41742, n41743, n41744, n41745, n41746, n41747, n41748, n41749, n41750, n41751, n41752, n41753, n41754, n41755, n41756, n41757, n41758, n41759, n41760, n41761, n41762, n41763, n41764, n41765, n41766, n41767, n41768, n41769, n41770, n41771, n41772, n41773, n41774, n41775, n41776, n41777, n41778, n41779, n41780, n41781, n41782, n41783, n41784, n41785, n41786, n41787, n41788, n41789, n41790, n41791, n41792, n41793, n41794, n41795, n41796, n41797, n41798, n41799, n41800, n41801, n41802, n41803, n41804, n41805, n41806, n41807, n41808, n41809, n41810, n41811, n41812, n41813, n41814, n41815, n41816, n41817, n41818, n41819, n41820, n41821, n41822, n41823, n41824, n41825, n41826, n41827, n41828, n41829, n41830, n41831, n41832, n41833, n41834, n41835, n41836, n41837, n41838, n41839, n41840, n41841, n41842, n41843, n41844, n41845, n41846, n41847, n41848, n41849, n41850, n41851, n41852, n41853, n41854, n41855, n41856, n41857, n41858, n41859, n41860, n41861, n41862, n41863, n41864, n41865, n41866, n41867, n41868, n41869, n41870, n41871, n41872, n41873, n41874, n41875, n41876, n41877, n41878, n41879, n41880, n41881, n41882, n41883, n41884, n41885, n41886, n41887, n41888, n41889, n41890, n41891, n41892, n41893, n41894, n41895, n41896, n41897, n41898, n41899, n41900, n41901, n41902, n41903, n41904, n41905, n41906, n41907, n41908, n41909, n41910, n41911, n41912, n41913, n41914, n41915, n41916, n41917, n41918, n41919, n41920, n41921, n41922, n41923, n41924, n41925, n41926, n41927, n41928, n41929, n41930, n41931, n41932, n41933, n41934, n41935, n41936, n41937, n41938, n41939, n41940, n41941, n41942, n41943, n41944, n41945, n41946, n41947, n41948, n41949, n41950, n41951, n41952, n41953, n41954, n41955, n41956, n41957, n41958, n41959, n41960, n41961, n41962, n41963, n41964, n41965, n41966, n41967, n41968, n41969, n41970, n41971, n41972, n41973, n41974, n41975, n41976, n41977, n41978, n41979, n41980, n41981, n41982, n41983, n41984, n41985, n41986, n41987, n41988, n41989, n41990, n41991, n41992, n41993, n41994, n41995, n41996, n41997, n41998, n41999, n42000, n42001, n42002, n42003, n42004, n42005, n42006, n42007, n42008, n42009, n42010, n42011, n42012, n42013, n42014, n42015, n42016, n42017, n42018, n42019, n42020, n42021, n42022, n42023, n42024, n42025, n42026, n42027, n42028, n42029, n42030, n42031, n42032, n42033, n42034, n42035, n42036, n42037, n42038, n42039, n42040, n42041, n42042, n42043, n42044, n42045, n42046, n42047, n42048, n42049, n42050, n42051, n42052, n42053, n42054, n42055, n42056, n42057, n42058, n42059, n42060, n42061, n42062, n42063, n42064, n42065, n42066, n42067, n42068, n42069, n42070, n42071, n42072, n42073, n42074, n42075, n42076, n42077, n42078, n42079, n42080, n42081, n42082, n42083, n42084, n42085, n42086, n42087, n42088, n42089, n42090, n42091, n42092, n42093, n42094, n42095, n42096, n42097, n42098, n42099, n42100, n42101, n42102, n42103, n42104, n42105, n42106, n42107, n42108, n42109, n42110, n42111, n42112, n42113, n42114, n42115, n42116, n42117, n42118, n42119, n42120, n42121, n42122, n42123, n42124, n42125, n42126, n42127, n42128, n42129, n42130, n42131, n42132, n42133, n42134, n42135, n42136, n42137, n42138, n42139, n42140, n42141, n42142, n42143, n42144, n42145, n42146, n42147, n42148, n42149, n42150, n42151, n42152, n42153, n42154, n42155, n42156, n42157, n42158, n42159, n42160, n42161, n42162, n42163, n42164, n42165, n42166, n42167, n42168, n42169, n42170, n42171, n42172, n42173, n42174, n42175, n42176, n42177, n42178, n42179, n42180, n42181, n42182, n42183, n42184, n42185, n42186, n42187, n42188, n42189, n42190, n42191, n42192, n42193, n42194, n42195, n42196, n42197, n42198, n42199, n42200, n42201, n42202, n42203, n42204, n42205, n42206, n42207, n42208, n42209, n42210, n42211, n42212, n42213, n42214, n42215, n42216, n42217, n42218, n42219, n42220, n42221, n42222, n42223, n42224, n42225, n42226, n42227, n42228, n42229, n42230, n42231, n42232, n42233, n42234, n42235, n42236, n42237, n42238, n42239, n42240, n42241, n42242, n42243, n42244, n42245, n42246, n42247, n42248, n42249, n42250, n42251, n42252, n42253, n42254, n42255, n42256, n42257, n42258, n42259, n42260, n42261, n42262, n42263, n42264, n42265, n42266, n42267, n42268, n42269, n42270, n42271, n42272, n42273, n42274, n42275, n42276, n42277, n42278, n42279, n42280, n42281, n42282, n42283, n42284, n42285, n42286, n42287, n42288, n42289, n42290, n42291, n42292, n42293, n42294, n42295, n42296, n42297, n42298, n42299, n42300, n42301, n42302, n42303, n42304, n42305, n42306, n42307, n42308, n42309, n42310, n42311, n42312, n42313, n42314, n42315, n42316, n42317, n42318, n42319, n42320, n42321, n42322, n42323, n42324, n42325, n42326, n42327, n42328, n42329, n42330, n42331, n42332, n42333, n42334, n42335, n42336, n42337, n42338, n42339, n42340, n42341, n42342, n42343, n42344, n42345, n42346, n42347, n42348, n42349, n42350, n42351, n42352, n42353, n42354, n42355, n42356, n42357, n42358, n42359, n42360, n42361, n42362, n42363, n42364, n42365, n42366, n42367, n42368, n42369, n42370, n42371, n42372, n42373, n42374, n42375, n42376, n42377, n42378, n42379, n42380, n42381, n42382, n42383, n42384, n42385, n42386, n42387, n42388, n42389, n42390, n42391, n42392, n42393, n42394, n42395, n42396, n42397, n42398, n42399, n42400, n42401, n42402, n42403, n42404, n42405, n42406, n42407, n42408, n42409, n42410, n42411, n42412, n42413, n42414, n42415, n42416, n42417, n42418, n42419, n42420, n42421, n42422, n42423, n42424, n42425, n42426, n42427, n42428, n42429, n42430, n42431, n42432, n42433, n42434, n42435, n42436, n42437, n42438, n42439, n42440, n42441, n42442, n42443, n42444, n42445, n42446, n42447, n42448, n42449, n42450, n42451, n42452, n42453, n42454, n42455, n42456, n42457, n42458, n42459, n42460, n42461, n42462, n42463, n42464, n42465, n42466, n42467, n42468, n42469, n42470, n42471, n42472, n42473, n42474, n42475, n42476, n42477, n42478, n42479, n42480, n42481, n42482, n42483, n42484, n42485, n42486, n42487, n42488, n42489, n42490, n42491, n42492, n42493, n42494, n42495, n42496, n42497, n42498, n42499, n42500, n42501, n42502, n42503, n42504, n42505, n42506, n42507, n42508, n42509, n42510, n42511, n42512, n42513, n42514, n42515, n42516, n42517, n42518, n42519, n42520, n42521, n42522, n42523, n42524, n42525, n42526, n42527, n42528, n42529, n42530, n42531, n42532, n42533, n42534, n42535, n42536, n42537, n42538, n42539, n42540, n42541, n42542, n42543, n42544, n42545, n42546, n42547, n42548, n42549, n42550, n42551, n42552, n42553, n42554, n42555, n42556, n42557, n42558, n42559, n42560, n42561, n42562, n42563, n42564, n42565, n42566, n42567, n42568, n42569, n42570, n42571, n42572, n42573, n42574, n42575, n42576, n42577, n42578, n42579, n42580, n42581, n42582, n42583, n42584, n42585, n42586, n42587, n42588, n42589, n42590, n42591, n42592, n42593, n42594, n42595, n42596, n42597, n42598, n42599, n42600, n42601, n42602, n42603, n42604, n42605, n42606, n42607, n42608, n42609, n42610, n42611, n42612, n42613, n42614, n42615, n42616, n42617, n42618, n42619, n42620, n42621, n42622, n42623, n42624, n42625, n42626, n42627, n42628, n42629, n42630, n42631, n42632, n42633, n42634, n42635, n42636, n42637, n42638, n42639, n42640, n42641, n42642, n42643, n42644, n42645, n42646, n42647, n42648, n42649, n42650, n42651, n42652, n42653, n42654, n42655, n42656, n42657, n42658, n42659, n42660, n42661, n42662, n42663, n42664, n42665, n42666, n42667, n42668, n42669, n42670, n42671, n42672, n42673, n42674, n42675, n42676, n42677, n42678, n42679, n42680, n42681, n42682, n42683, n42684, n42685, n42686, n42687, n42688, n42689, n42690, n42691, n42692, n42693, n42694, n42695, n42696, n42697, n42698, n42699, n42700, n42701, n42702, n42703, n42704, n42705, n42706, n42707, n42708, n42709, n42710, n42711, n42712, n42713, n42714, n42715, n42716, n42717, n42718, n42719, n42720, n42721, n42722, n42723, n42724, n42725, n42726, n42727, n42728, n42729, n42730, n42731, n42732, n42733, n42734, n42735, n42736, n42737, n42738, n42739, n42740, n42741, n42742, n42743, n42744, n42745, n42746, n42747, n42748, n42749, n42750, n42751, n42752, n42753, n42754, n42755, n42756, n42757, n42758, n42759, n42760, n42761, n42762, n42763, n42764, n42765, n42766, n42767, n42768, n42769, n42770, n42771, n42772, n42773, n42774, n42775, n42776, n42777, n42778, n42779, n42780, n42781, n42782, n42783, n42784, n42785, n42786, n42787, n42788, n42789, n42790, n42791, n42792, n42793, n42794, n42795, n42796, n42797, n42798, n42799, n42800, n42801, n42802, n42803, n42804, n42805, n42806, n42807, n42808, n42809, n42810, n42811, n42812, n42813, n42814, n42815, n42816, n42817, n42818, n42819, n42820, n42821, n42822, n42823, n42824, n42825, n42826, n42827, n42828, n42829, n42830, n42831, n42832, n42833, n42834, n42835, n42836, n42837, n42838, n42839, n42840, n42841, n42842, n42843, n42844, n42845, n42846, n42847, n42848, n42849, n42850, n42851, n42852, n42853, n42854, n42855, n42856, n42857, n42858, n42859, n42860, n42861, n42862, n42863, n42864, n42865, n42866, n42867, n42868, n42869, n42870, n42871, n42872, n42873, n42874, n42875, n42876, n42877, n42878, n42879, n42880, n42881, n42882, n42883, n42884, n42885, n42886, n42887, n42888, n42889, n42890, n42891, n42892, n42893, n42894, n42895, n42896, n42897, n42898, n42899, n42900, n42901, n42902, n42903, n42904, n42905, n42906, n42907, n42908, n42909, n42910, n42911, n42912, n42913, n42914, n42915, n42916, n42917, n42918, n42919, n42920, n42921, n42922, n42923, n42924, n42925, n42926, n42927, n42928, n42929, n42930, n42931, n42932, n42933, n42934, n42935, n42936, n42937, n42938, n42939, n42940, n42941, n42942, n42943, n42944, n42945, n42946, n42947, n42948, n42949, n42950, n42951, n42952, n42953, n42954, n42955, n42956, n42957, n42958, n42959, n42960, n42961, n42962, n42963, n42964, n42965, n42966, n42967, n42968, n42969, n42970, n42971, n42972, n42973, n42974, n42975, n42976, n42977, n42978, n42979, n42980, n42981, n42982, n42983, n42984, n42985, n42986, n42987, n42988, n42989, n42990, n42991, n42992, n42993, n42994, n42995, n42996, n42997, n42998, n42999, n43000, n43001, n43002, n43003, n43004, n43005, n43006, n43007, n43008, n43009, n43010, n43011, n43012, n43013, n43014, n43015, n43016, n43017, n43018, n43019, n43020, n43021, n43022, n43023, n43024, n43025, n43026, n43027, n43028, n43029, n43030, n43031, n43032, n43033, n43034, n43035, n43036, n43037, n43038, n43039, n43040, n43041, n43042, n43043, n43044, n43045, n43046, n43047, n43048, n43049, n43050, n43051, n43052, n43053, n43054, n43055, n43056, n43057, n43058, n43059, n43060, n43061, n43062, n43063, n43064, n43065, n43066, n43067, n43068, n43069, n43070, n43071, n43072, n43073, n43074, n43075, n43076, n43077, n43078, n43079, n43080, n43081, n43082, n43083, n43084, n43085, n43086, n43087, n43088, n43089, n43090, n43091, n43092, n43093, n43094, n43095, n43096, n43097, n43098, n43099, n43100, n43101, n43102, n43103, n43104, n43105, n43106, n43107, n43108, n43109, n43110, n43111, n43112, n43113, n43114, n43115, n43116, n43117, n43118, n43119, n43120, n43121, n43122, n43123, n43124, n43125, n43126, n43127, n43128, n43129, n43130, n43131, n43132, n43133, n43134, n43135, n43136, n43137, n43138, n43139, n43140, n43141, n43142, n43143, n43144, n43145, n43146, n43147, n43148, n43149, n43150, n43151, n43152, n43153, n43154, n43155, n43156, n43157, n43158, n43159, n43160, n43161, n43162, n43163, n43164, n43165, n43166, n43167, n43168, n43169, n43170, n43171, n43172, n43173, n43174, n43175, n43176, n43177, n43178, n43179, n43180, n43181, n43182, n43183, n43184, n43185, n43186, n43187, n43188, n43189, n43190, n43191, n43192, n43193, n43194, n43195, n43196, n43197, n43198, n43199, n43200, n43201, n43202, n43203, n43204, n43205, n43206, n43207, n43208, n43209, n43210, n43211, n43212, n43213, n43214, n43215, n43216, n43217, n43218, n43219, n43220, n43221, n43222, n43223, n43224, n43225, n43226, n43227, n43228, n43229, n43230, n43231, n43232, n43233, n43234, n43235, n43236, n43237, n43238, n43239, n43240, n43241, n43242, n43243, n43244, n43245, n43246, n43247, n43248, n43249, n43250, n43251, n43252, n43253, n43254, n43255, n43256, n43257, n43258, n43259, n43260, n43261, n43262, n43263, n43264, n43265, n43266, n43267, n43268, n43269, n43270, n43271, n43272, n43273, n43274, n43275, n43276, n43277, n43278, n43279, n43280, n43281, n43282, n43283, n43284, n43285, n43286, n43287, n43288, n43289, n43290, n43291, n43292, n43293, n43294, n43295, n43296, n43297, n43298, n43299, n43300, n43301, n43302, n43303, n43304, n43305, n43306, n43307, n43308, n43309, n43310, n43311, n43312, n43313, n43314, n43315, n43316, n43317, n43318, n43319, n43320, n43321, n43322, n43323, n43324, n43325, n43326, n43327, n43328, n43329, n43330, n43331, n43332, n43333, n43334, n43335, n43336, n43337, n43338, n43339, n43340, n43341, n43342, n43343, n43344, n43345, n43346, n43347, n43348, n43349, n43350, n43351, n43352, n43353, n43354, n43355, n43356, n43357, n43358, n43359, n43360, n43361, n43362, n43363, n43364, n43365, n43366, n43367, n43368, n43369, n43370, n43371, n43372, n43373, n43374, n43375, n43376, n43377, n43378, n43379, n43380, n43381, n43382, n43383, n43384, n43385, n43386, n43387, n43388, n43389, n43390, n43391, n43392, n43393, n43394, n43395, n43396, n43397, n43398, n43399, n43400, n43401, n43402, n43403, n43404, n43405, n43406, n43407, n43408, n43409, n43410, n43411, n43412, n43413, n43414, n43415, n43416, n43417, n43418, n43419, n43420, n43421, n43422, n43423, n43424, n43425, n43426, n43427, n43428, n43429, n43430, n43431, n43432, n43433, n43434, n43435, n43436, n43437, n43438, n43439, n43440, n43441, n43442, n43443, n43444, n43445, n43446, n43447, n43448, n43449, n43450, n43451, n43452, n43453, n43454, n43455, n43456, n43457, n43458, n43459, n43460, n43461, n43462, n43463, n43464, n43465, n43466, n43467, n43468, n43469, n43470, n43471, n43472, n43473, n43474, n43475, n43476, n43477, n43478, n43479, n43480, n43481, n43482, n43483, n43484, n43485, n43486, n43487, n43488, n43489, n43490, n43491, n43492, n43493, n43494, n43495, n43496, n43497, n43498, n43499, n43500, n43501, n43502, n43503, n43504, n43505, n43506, n43507, n43508, n43509, n43510, n43511, n43512, n43513, n43514, n43515, n43516, n43517, n43518, n43519, n43520, n43521, n43522, n43523, n43524, n43525, n43526, n43527, n43528, n43529, n43530, n43531, n43532, n43533, n43534, n43535, n43536, n43537, n43538, n43539, n43540, n43541, n43542, n43543, n43544, n43545, n43546, n43547, n43548, n43549, n43550, n43551, n43552, n43553, n43554, n43555, n43556, n43557, n43558, n43559, n43560, n43561, n43562, n43563, n43564, n43565, n43566, n43567, n43568, n43569, n43570, n43571, n43572, n43573, n43574, n43575, n43576, n43577, n43578, n43579, n43580, n43581, n43582, n43583, n43584, n43585, n43586, n43587, n43588, n43589, n43590, n43591, n43592, n43593, n43594, n43595, n43596, n43597, n43598, n43599, n43600, n43601, n43602, n43603, n43604, n43605, n43606, n43607, n43608, n43609, n43610, n43611, n43612, n43613, n43614, n43615, n43616, n43617, n43618, n43619, n43620, n43621, n43622, n43623, n43624, n43625, n43626, n43627, n43628, n43629, n43630, n43631, n43632, n43633, n43634, n43635, n43636, n43637, n43638, n43639, n43640, n43641, n43642, n43643, n43644, n43645, n43646, n43647, n43648, n43649, n43650, n43651, n43652, n43653, n43654, n43655, n43656, n43657, n43658, n43659, n43660, n43661, n43662, n43663, n43664, n43665, n43666, n43667, n43668, n43669, n43670, n43671, n43672, n43673, n43674, n43675, n43676, n43677, n43678, n43679, n43680, n43681, n43682, n43683, n43684, n43685, n43686, n43687, n43688, n43689, n43690, n43691, n43692, n43693, n43694, n43695, n43696, n43697, n43698, n43699, n43700, n43701, n43702, n43703, n43704, n43705, n43706, n43707, n43708, n43709, n43710, n43711, n43712, n43713, n43714, n43715, n43716, n43717, n43718, n43719, n43720, n43721, n43722, n43723, n43724, n43725, n43726, n43727, n43728, n43729, n43730, n43731, n43732, n43733, n43734, n43735, n43736, n43737, n43738, n43739, n43740, n43741, n43742, n43743, n43744, n43745, n43746, n43747, n43748, n43749, n43750, n43751, n43752, n43753, n43754, n43755, n43756, n43757, n43758, n43759, n43760, n43761, n43762, n43763, n43764, n43765, n43766, n43767, n43768, n43769, n43770, n43771, n43772, n43773, n43774, n43775, n43776, n43777, n43778, n43779, n43780, n43781, n43782, n43783, n43784, n43785, n43786, n43787, n43788, n43789, n43790, n43791, n43792, n43793, n43794, n43795, n43796, n43797, n43798, n43799, n43800, n43801, n43802, n43803, n43804, n43805, n43806, n43807, n43808, n43809, n43810, n43811, n43812, n43813, n43814, n43815, n43816, n43817, n43818, n43819, n43820, n43821, n43822, n43823, n43824, n43825, n43826, n43827, n43828, n43829, n43830, n43831, n43832, n43833, n43834, n43835, n43836, n43837, n43838, n43839, n43840, n43841, n43842, n43843, n43844, n43845, n43846, n43847, n43848, n43849, n43850, n43851, n43852, n43853, n43854, n43855, n43856, n43857, n43858, n43859, n43860, n43861, n43862, n43863, n43864, n43865, n43866, n43867, n43868, n43869, n43870, n43871, n43872, n43873, n43874, n43875, n43876, n43877, n43878, n43879, n43880, n43881, n43882, n43883, n43884, n43885, n43886, n43887, n43888, n43889, n43890, n43891, n43892, n43893, n43894, n43895, n43896, n43897, n43898, n43899, n43900, n43901, n43902, n43903, n43904, n43905, n43906, n43907, n43908, n43909, n43910, n43911, n43912, n43913, n43914, n43915, n43916, n43917, n43918, n43919, n43920, n43921, n43922, n43923, n43924, n43925, n43926, n43927, n43928, n43929, n43930, n43931, n43932, n43933, n43934, n43935, n43936, n43937, n43938, n43939, n43940, n43941, n43942, n43943, n43944, n43945, n43946, n43947, n43948, n43949, n43950, n43951, n43952, n43953, n43954, n43955, n43956, n43957, n43958, n43959, n43960, n43961, n43962, n43963, n43964, n43965, n43966, n43967, n43968, n43969, n43970, n43971, n43972, n43973, n43974, n43975, n43976, n43977, n43978, n43979, n43980, n43981, n43982, n43983, n43984, n43985, n43986, n43987, n43988, n43989, n43990, n43991, n43992, n43993, n43994, n43995, n43996, n43997, n43998, n43999, n44000, n44001, n44002, n44003, n44004, n44005, n44006, n44007, n44008, n44009, n44010, n44011, n44012, n44013, n44014, n44015, n44016, n44017, n44018, n44019, n44020, n44021, n44022, n44023, n44024, n44025, n44026, n44027, n44028, n44029, n44030, n44031, n44032, n44033, n44034, n44035, n44036, n44037, n44038, n44039, n44040, n44041, n44042, n44043, n44044, n44045, n44046, n44047, n44048, n44049, n44050, n44051, n44052, n44053, n44054, n44055, n44056, n44057, n44058, n44059, n44060, n44061, n44062, n44063, n44064, n44065, n44066, n44067, n44068, n44069, n44070, n44071, n44072, n44073, n44074, n44075, n44076, n44077, n44078, n44079, n44080, n44081, n44082, n44083, n44084, n44085, n44086, n44087, n44088, n44089, n44090, n44091, n44092, n44093, n44094, n44095, n44096, n44097, n44098, n44099, n44100, n44101, n44102, n44103, n44104, n44105, n44106, n44107, n44108, n44109, n44110, n44111, n44112, n44113, n44114, n44115, n44116, n44117, n44118, n44119, n44120, n44121, n44122, n44123, n44124, n44125, n44126, n44127, n44128, n44129, n44130, n44131, n44132, n44133, n44134, n44135, n44136, n44137, n44138, n44139, n44140, n44141, n44142, n44143, n44144, n44145, n44146, n44147, n44148, n44149, n44150, n44151, n44152, n44153, n44154, n44155, n44156, n44157, n44158, n44159, n44160, n44161, n44162, n44163, n44164, n44165, n44166, n44167, n44168, n44169, n44170, n44171, n44172, n44173, n44174, n44175, n44176, n44177, n44178, n44179, n44180, n44181, n44182, n44183, n44184, n44185, n44186, n44187, n44188, n44189, n44190, n44191, n44192, n44193, n44194, n44195, n44196, n44197, n44198, n44199, n44200, n44201, n44202, n44203, n44204, n44205, n44206, n44207, n44208, n44209, n44210, n44211, n44212, n44213, n44214, n44215, n44216, n44217, n44218, n44219, n44220, n44221, n44222, n44223, n44224, n44225, n44226, n44227, n44228, n44229, n44230, n44231, n44232, n44233, n44234, n44235, n44236, n44237, n44238, n44239, n44240, n44241, n44242, n44243, n44244, n44245, n44246, n44247, n44248, n44249, n44250, n44251, n44252, n44253, n44254, n44255, n44256, n44257, n44258, n44259, n44260, n44261, n44262, n44263, n44264, n44265, n44266, n44267, n44268, n44269, n44270, n44271, n44272, n44273, n44274, n44275, n44276, n44277, n44278, n44279, n44280, n44281, n44282, n44283, n44284, n44285, n44286, n44287, n44288, n44289, n44290, n44291, n44292, n44293, n44294, n44295, n44296, n44297, n44298, n44299, n44300, n44301, n44302, n44303, n44304, n44305, n44306, n44307, n44308, n44309, n44310, n44311, n44312, n44313, n44314, n44315, n44316, n44317, n44318, n44319, n44320, n44321, n44322, n44323, n44324, n44325, n44326, n44327, n44328, n44329, n44330, n44331, n44332, n44333, n44334, n44335, n44336, n44337, n44338, n44339, n44340, n44341, n44342, n44343, n44344, n44345, n44346, n44347, n44348, n44349, n44350, n44351, n44352, n44353, n44354, n44355, n44356, n44357, n44358, n44359, n44360, n44361, n44362, n44363, n44364, n44365, n44366, n44367, n44368, n44369, n44370, n44371, n44372, n44373, n44374, n44375, n44376, n44377, n44378, n44379, n44380, n44381, n44382, n44383, n44384, n44385, n44386, n44387, n44388, n44389, n44390, n44391, n44392, n44393, n44394, n44395, n44396, n44397, n44398, n44399, n44400, n44401, n44402, n44403, n44404, n44405, n44406, n44407, n44408, n44409, n44410, n44411, n44412, n44413, n44414, n44415, n44416, n44417, n44418, n44419, n44420, n44421, n44422, n44423, n44424, n44425, n44426, n44427, n44428, n44429, n44430, n44431, n44432, n44433, n44434, n44435, n44436, n44437, n44438, n44439, n44440, n44441, n44442, n44443, n44444, n44445, n44446, n44447, n44448, n44449, n44450, n44451, n44452, n44453, n44454, n44455, n44456, n44457, n44458, n44459, n44460, n44461, n44462, n44463, n44464, n44465, n44466, n44467, n44468, n44469, n44470, n44471, n44472, n44473, n44474, n44475, n44476, n44477, n44478, n44479, n44480, n44481, n44482, n44483, n44484, n44485, n44486, n44487, n44488, n44489, n44490, n44491, n44492, n44493, n44494, n44495, n44496, n44497, n44498, n44499, n44500, n44501, n44502, n44503, n44504, n44505, n44506, n44507, n44508, n44509, n44510, n44511, n44512, n44513, n44514, n44515, n44516, n44517, n44518, n44519, n44520, n44521, n44522, n44523, n44524, n44525, n44526, n44527, n44528, n44529, n44530, n44531, n44532, n44533, n44534, n44535, n44536, n44537, n44538, n44539, n44540, n44541, n44542, n44543, n44544, n44545, n44546, n44547, n44548, n44549, n44550, n44551, n44552, n44553, n44554, n44555, n44556, n44557, n44558, n44559, n44560, n44561, n44562, n44563, n44564, n44565, n44566, n44567, n44568, n44569, n44570, n44571, n44572, n44573, n44574, n44575, n44576, n44577, n44578, n44579, n44580, n44581, n44582, n44583, n44584, n44585, n44586, n44587, n44588, n44589, n44590, n44591, n44592, n44593, n44594, n44595, n44596, n44597, n44598, n44599, n44600, n44601, n44602, n44603, n44604, n44605, n44606, n44607, n44608, n44609, n44610, n44611, n44612, n44613, n44614, n44615, n44616, n44617, n44618, n44619, n44620, n44621, n44622, n44623, n44624, n44625, n44626, n44627, n44628, n44629, n44630, n44631, n44632, n44633, n44634, n44635, n44636, n44637, n44638, n44639, n44640, n44641, n44642, n44643, n44644, n44645, n44646, n44647, n44648, n44649, n44650, n44651, n44652, n44653, n44654, n44655, n44656, n44657, n44658, n44659, n44660, n44661, n44662, n44663, n44664, n44665, n44666, n44667, n44668, n44669, n44670, n44671, n44672, n44673, n44674, n44675, n44676, n44677, n44678, n44679, n44680, n44681, n44682, n44683, n44684, n44685, n44686, n44687, n44688, n44689, n44690, n44691, n44692, n44693, n44694, n44695, n44696, n44697, n44698, n44699, n44700, n44701, n44702, n44703, n44704, n44705, n44706, n44707, n44708, n44709, n44710, n44711, n44712, n44713, n44714, n44715, n44716, n44717, n44718, n44719, n44720, n44721, n44722, n44723, n44724, n44725, n44726, n44727, n44728, n44729, n44730, n44731, n44732, n44733, n44734, n44735, n44736, n44737, n44738, n44739, n44740, n44741, n44742, n44743, n44744, n44745, n44746, n44747, n44748, n44749, n44750, n44751, n44752, n44753, n44754, n44755, n44756, n44757, n44758, n44759, n44760, n44761, n44762, n44763, n44764, n44765, n44766, n44767, n44768, n44769, n44770, n44771, n44772, n44773, n44774, n44775, n44776, n44777, n44778, n44779, n44780, n44781, n44782, n44783, n44784, n44785, n44786, n44787, n44788, n44789, n44790, n44791, n44792, n44793, n44794, n44795, n44796, n44797, n44798, n44799, n44800, n44801, n44802, n44803, n44804, n44805, n44806, n44807, n44808, n44809, n44810, n44811, n44812, n44813, n44814, n44815, n44816, n44817, n44818, n44819, n44820, n44821, n44822, n44823, n44824, n44825, n44826, n44827, n44828, n44829, n44830, n44831, n44832, n44833, n44834, n44835, n44836, n44837, n44838, n44839, n44840, n44841, n44842, n44843, n44844, n44845, n44846, n44847, n44848, n44849, n44850, n44851, n44852, n44853, n44854, n44855, n44856, n44857, n44858, n44859, n44860, n44861, n44862, n44863, n44864, n44865, n44866, n44867, n44868, n44869, n44870, n44871, n44872, n44873, n44874, n44875, n44876, n44877, n44878, n44879, n44880, n44881, n44882, n44883, n44884, n44885, n44886, n44887, n44888, n44889, n44890, n44891, n44892, n44893, n44894, n44895, n44896, n44897, n44898, n44899, n44900, n44901, n44902, n44903, n44904, n44905, n44906, n44907, n44908, n44909, n44910, n44911, n44912, n44913, n44914, n44915, n44916, n44917, n44918, n44919, n44920, n44921, n44922, n44923, n44924, n44925, n44926, n44927, n44928, n44929, n44930, n44931, n44932, n44933, n44934, n44935, n44936, n44937, n44938, n44939, n44940, n44941, n44942, n44943, n44944, n44945, n44946, n44947, n44948, n44949, n44950, n44951, n44952, n44953, n44954, n44955, n44956, n44957, n44958, n44959, n44960, n44961, n44962, n44963, n44964, n44965, n44966, n44967, n44968, n44969, n44970, n44971, n44972, n44973, n44974, n44975, n44976, n44977, n44978, n44979, n44980, n44981, n44982, n44983, n44984, n44985, n44986, n44987, n44988, n44989, n44990, n44991, n44992, n44993, n44994, n44995, n44996, n44997, n44998, n44999, n45000, n45001, n45002, n45003, n45004, n45005, n45006, n45007, n45008, n45009, n45010, n45011, n45012, n45013, n45014, n45015, n45016, n45017, n45018, n45019, n45020, n45021, n45022, n45023, n45024, n45025, n45026, n45027, n45028, n45029, n45030, n45031, n45032, n45033, n45034, n45035, n45036, n45037, n45038, n45039, n45040, n45041, n45042, n45043, n45044, n45045, n45046, n45047, n45048, n45049, n45050, n45051, n45052, n45053, n45054, n45055, n45056, n45057, n45058, n45059, n45060, n45061, n45062, n45063, n45064, n45065, n45066, n45067, n45068, n45069, n45070, n45071, n45072, n45073, n45074, n45075, n45076, n45077, n45078, n45079, n45080, n45081, n45082, n45083, n45084, n45085, n45086, n45087, n45088, n45089, n45090, n45091, n45092, n45093, n45094, n45095, n45096, n45097, n45098, n45099, n45100, n45101, n45102, n45103, n45104, n45105, n45106, n45107, n45108, n45109, n45110, n45111, n45112, n45113, n45114, n45115, n45116, n45117, n45118, n45119, n45120, n45121, n45122, n45123, n45124, n45125, n45126, n45127, n45128, n45129, n45130, n45131, n45132, n45133, n45134, n45135, n45136, n45137, n45138, n45139, n45140, n45141, n45142, n45143, n45144, n45145, n45146, n45147, n45148, n45149, n45150, n45151, n45152, n45153, n45154, n45155, n45156, n45157, n45158, n45159, n45160, n45161, n45162, n45163, n45164, n45165, n45166, n45167, n45168, n45169, n45170, n45171, n45172, n45173, n45174, n45175, n45176, n45177, n45178, n45179, n45180, n45181, n45182, n45183, n45184, n45185, n45186, n45187, n45188, n45189, n45190, n45191, n45192, n45193, n45194, n45195, n45196, n45197, n45198, n45199, n45200, n45201, n45202, n45203, n45204, n45205, n45206, n45207, n45208, n45209, n45210, n45211, n45212, n45213, n45214, n45215, n45216, n45217, n45218, n45219, n45220, n45221, n45222, n45223, n45224, n45225, n45226, n45227, n45228, n45229, n45230, n45231, n45232, n45233, n45234, n45235, n45236, n45237, n45238, n45239, n45240, n45241, n45242, n45243, n45244, n45245, n45246, n45247, n45248, n45249, n45250, n45251, n45252, n45253, n45254, n45255, n45256, n45257, n45258, n45259, n45260, n45261, n45262, n45263, n45264, n45265, n45266, n45267, n45268, n45269, n45270, n45271, n45272, n45273, n45274, n45275, n45276, n45277, n45278, n45279, n45280, n45281, n45282, n45283, n45284, n45285, n45286, n45287, n45288, n45289, n45290, n45291, n45292, n45293, n45294, n45295, n45296, n45297, n45298, n45299, n45300, n45301, n45302, n45303, n45304, n45305, n45306, n45307, n45308, n45309, n45310, n45311, n45312, n45313, n45314, n45315, n45316, n45317, n45318, n45319, n45320, n45321, n45322, n45323, n45324, n45325, n45326, n45327, n45328, n45329, n45330, n45331, n45332, n45333, n45334, n45335, n45336, n45337, n45338, n45339, n45340, n45341, n45342, n45343, n45344, n45345, n45346, n45347, n45348, n45349, n45350, n45351, n45352, n45353, n45354, n45355, n45356, n45357, n45358, n45359, n45360, n45361, n45362, n45363, n45364, n45365, n45366, n45367, n45368, n45369, n45370, n45371, n45372, n45373, n45374, n45375, n45376, n45377, n45378, n45379, n45380, n45381, n45382, n45383, n45384, n45385, n45386, n45387, n45388, n45389, n45390, n45391, n45392, n45393, n45394, n45395, n45396, n45397, n45398, n45399, n45400, n45401, n45402, n45403, n45404, n45405, n45406, n45407, n45408, n45409, n45410, n45411, n45412, n45413, n45414, n45415, n45416, n45417, n45418, n45419, n45420, n45421, n45422, n45423, n45424, n45425, n45426, n45427, n45428, n45429, n45430, n45431, n45432, n45433, n45434, n45435, n45436, n45437, n45438, n45439, n45440, n45441, n45442, n45443, n45444, n45445, n45446, n45447, n45448, n45449, n45450, n45451, n45452, n45453, n45454, n45455, n45456, n45457, n45458, n45459, n45460, n45461, n45462, n45463, n45464, n45465, n45466, n45467, n45468, n45469, n45470, n45471, n45472, n45473, n45474, n45475, n45476, n45477, n45478, n45479, n45480, n45481, n45482, n45483, n45484, n45485, n45486, n45487, n45488, n45489, n45490, n45491, n45492, n45493, n45494, n45495, n45496, n45497, n45498, n45499, n45500, n45501, n45502, n45503, n45504, n45505, n45506, n45507, n45508, n45509, n45510, n45511, n45512, n45513, n45514, n45515, n45516, n45517, n45518, n45519, n45520, n45521, n45522, n45523, n45524, n45525, n45526, n45527, n45528, n45529, n45530, n45531, n45532, n45533, n45534, n45535, n45536, n45537, n45538, n45539, n45540, n45541, n45542, n45543, n45544, n45545, n45546, n45547, n45548, n45549, n45550, n45551, n45552, n45553, n45554, n45555, n45556, n45557, n45558, n45559, n45560, n45561, n45562, n45563, n45564, n45565, n45566, n45567, n45568, n45569, n45570, n45571, n45572, n45573, n45574, n45575, n45576, n45577, n45578, n45579, n45580, n45581, n45582, n45583, n45584, n45585, n45586, n45587, n45588, n45589, n45590, n45591, n45592, n45593, n45594, n45595, n45596, n45597, n45598, n45599, n45600, n45601, n45602, n45603, n45604, n45605, n45606, n45607, n45608, n45609, n45610, n45611, n45612, n45613, n45614, n45615, n45616, n45617, n45618, n45619, n45620, n45621, n45622, n45623, n45624, n45625, n45626, n45627, n45628, n45629, n45630, n45631, n45632, n45633, n45634, n45635, n45636, n45637, n45638, n45639, n45640, n45641, n45642, n45643, n45644, n45645, n45646, n45647, n45648, n45649, n45650, n45651, n45652, n45653, n45654, n45655, n45656, n45657, n45658, n45659, n45660, n45661, n45662, n45663, n45664, n45665, n45666, n45667, n45668, n45669, n45670, n45671, n45672, n45673, n45674, n45675, n45676, n45677, n45678, n45679, n45680, n45681, n45682, n45683, n45684, n45685, n45686, n45687, n45688, n45689, n45690, n45691, n45692, n45693, n45694, n45695, n45696, n45697, n45698, n45699, n45700, n45701, n45702, n45703, n45704, n45705, n45706, n45707, n45708, n45709, n45710, n45711, n45712, n45713, n45714, n45715, n45716, n45717, n45718, n45719, n45720, n45721, n45722, n45723, n45724, n45725, n45726, n45727, n45728, n45729, n45730, n45731, n45732, n45733, n45734, n45735, n45736, n45737, n45738, n45739, n45740, n45741, n45742, n45743, n45744, n45745, n45746, n45747, n45748, n45749, n45750, n45751, n45752, n45753, n45754, n45755, n45756, n45757, n45758, n45759, n45760, n45761, n45762, n45763, n45764, n45765, n45766, n45767, n45768, n45769, n45770, n45771, n45772, n45773, n45774, n45775, n45776, n45777, n45778, n45779, n45780, n45781, n45782, n45783, n45784, n45785, n45786, n45787, n45788, n45789, n45790, n45791, n45792, n45793, n45794, n45795, n45796, n45797, n45798, n45799, n45800, n45801, n45802, n45803, n45804, n45805, n45806, n45807, n45808, n45809, n45810, n45811, n45812, n45813, n45814, n45815, n45816, n45817, n45818, n45819, n45820, n45821, n45822, n45823, n45824, n45825, n45826, n45827, n45828, n45829, n45830, n45831, n45832, n45833, n45834, n45835, n45836, n45837, n45838, n45839, n45840, n45841, n45842, n45843, n45844, n45845, n45846, n45847, n45848, n45849, n45850, n45851, n45852, n45853, n45854, n45855, n45856, n45857, n45858, n45859, n45860, n45861, n45862, n45863, n45864, n45865, n45866, n45867, n45868, n45869, n45870, n45871, n45872, n45873, n45874, n45875, n45876, n45877, n45878, n45879, n45880, n45881, n45882, n45883, n45884, n45885, n45886, n45887, n45888, n45889, n45890, n45891, n45892, n45893, n45894, n45895, n45896, n45897, n45898, n45899, n45900, n45901, n45902, n45903, n45904, n45905, n45906, n45907, n45908, n45909, n45910, n45911, n45912, n45913, n45914, n45915, n45916, n45917, n45918, n45919, n45920, n45921, n45922, n45923, n45924, n45925, n45926, n45927, n45928, n45929, n45930, n45931, n45932, n45933, n45934, n45935, n45936, n45937, n45938, n45939, n45940, n45941, n45942, n45943, n45944, n45945, n45946, n45947, n45948, n45949, n45950, n45951, n45952, n45953, n45954, n45955, n45956, n45957, n45958, n45959, n45960, n45961, n45962, n45963, n45964, n45965, n45966, n45967, n45968, n45969, n45970, n45971, n45972, n45973, n45974, n45975, n45976, n45977, n45978, n45979, n45980, n45981, n45982, n45983, n45984, n45985, n45986, n45987, n45988, n45989, n45990, n45991, n45992, n45993, n45994, n45995, n45996, n45997, n45998, n45999, n46000, n46001, n46002, n46003, n46004, n46005, n46006, n46007, n46008, n46009, n46010, n46011, n46012, n46013, n46014, n46015, n46016, n46017, n46018, n46019, n46020, n46021, n46022, n46023, n46024, n46025, n46026, n46027, n46028, n46029, n46030, n46031, n46032, n46033, n46034, n46035, n46036, n46037, n46038, n46039, n46040, n46041, n46042, n46043, n46044, n46045, n46046, n46047, n46048, n46049, n46050, n46051, n46052, n46053, n46054, n46055, n46056, n46057, n46058, n46059, n46060, n46061, n46062, n46063, n46064, n46065, n46066, n46067, n46068, n46069, n46070, n46071, n46072, n46073, n46074, n46075, n46076, n46077, n46078, n46079, n46080, n46081, n46082, n46083, n46084, n46085, n46086, n46087, n46088, n46089, n46090, n46091, n46092, n46093, n46094, n46095, n46096, n46097, n46098, n46099, n46100, n46101, n46102, n46103, n46104, n46105, n46106, n46107, n46108, n46109, n46110, n46111, n46112, n46113, n46114, n46115, n46116, n46117, n46118, n46119, n46120, n46121, n46122, n46123, n46124, n46125, n46126, n46127, n46128, n46129, n46130, n46131, n46132, n46133, n46134, n46135, n46136, n46137, n46138, n46139, n46140, n46141, n46142, n46143, n46144, n46145, n46146, n46147, n46148, n46149, n46150, n46151, n46152, n46153, n46154, n46155, n46156, n46157, n46158, n46159, n46160, n46161, n46162, n46163, n46164, n46165, n46166, n46167, n46168, n46169, n46170, n46171, n46172, n46173, n46174, n46175, n46176, n46177, n46178, n46179, n46180, n46181, n46182, n46183, n46184, n46185, n46186, n46187, n46188, n46189, n46190, n46191, n46192, n46193, n46194, n46195, n46196, n46197, n46198, n46199, n46200, n46201, n46202, n46203, n46204, n46205, n46206, n46207, n46208, n46209, n46210, n46211, n46212, n46213, n46214, n46215, n46216, n46217, n46218, n46219, n46220, n46221, n46222, n46223, n46224, n46225, n46226, n46227, n46228, n46229, n46230, n46231, n46232, n46233, n46234, n46235, n46236, n46237, n46238, n46239, n46240, n46241, n46242, n46243, n46244, n46245, n46246, n46247, n46248, n46249, n46250, n46251, n46252, n46253, n46254, n46255, n46256, n46257, n46258, n46259, n46260, n46261, n46262, n46263, n46264, n46265, n46266, n46267, n46268, n46269, n46270, n46271, n46272, n46273, n46274, n46275, n46276, n46277, n46278, n46279, n46280, n46281, n46282, n46283, n46284, n46285, n46286, n46287, n46288, n46289, n46290, n46291, n46292, n46293, n46294, n46295, n46296, n46297, n46298, n46299, n46300, n46301, n46302, n46303, n46304, n46305, n46306, n46307, n46308, n46309, n46310, n46311, n46312, n46313, n46314, n46315, n46316, n46317, n46318, n46319, n46320, n46321, n46322, n46323, n46324, n46325, n46326, n46327, n46328, n46329, n46330, n46331, n46332, n46333, n46334, n46335, n46336, n46337, n46338, n46339, n46340, n46341, n46342, n46343, n46344, n46345, n46346, n46347, n46348, n46349, n46350, n46351, n46352, n46353, n46354, n46355, n46356, n46357, n46358, n46359, n46360, n46361, n46362, n46363, n46364, n46365, n46366, n46367, n46368, n46369, n46370, n46371, n46372, n46373, n46374, n46375, n46376, n46377, n46378, n46379, n46380, n46381, n46382, n46383, n46384, n46385, n46386, n46387, n46388, n46389, n46390, n46391, n46392, n46393, n46394, n46395, n46396, n46397, n46398, n46399, n46400, n46401, n46402, n46403, n46404, n46405, n46406, n46407, n46408, n46409, n46410, n46411, n46412, n46413, n46414, n46415, n46416, n46417, n46418, n46419, n46420, n46421, n46422, n46423, n46424, n46425, n46426, n46427, n46428, n46429, n46430, n46431, n46432, n46433, n46434, n46435, n46436, n46437, n46438, n46439, n46440, n46441, n46442, n46443, n46444, n46445, n46446, n46447, n46448, n46449, n46450, n46451, n46452, n46453, n46454, n46455, n46456, n46457, n46458, n46459, n46460, n46461, n46462, n46463, n46464, n46465, n46466, n46467, n46468, n46469, n46470, n46471, n46472, n46473, n46474, n46475, n46476, n46477, n46478, n46479, n46480, n46481, n46482, n46483, n46484, n46485, n46486, n46487, n46488, n46489, n46490, n46491, n46492, n46493, n46494, n46495, n46496, n46497, n46498, n46499, n46500, n46501, n46502, n46503, n46504, n46505, n46506, n46507, n46508, n46509, n46510, n46511, n46512, n46513, n46514, n46515, n46516, n46517, n46518, n46519, n46520, n46521, n46522, n46523, n46524, n46525, n46526, n46527, n46528, n46529, n46530, n46531, n46532, n46533, n46534, n46535, n46536, n46537, n46538, n46539, n46540, n46541, n46542, n46543, n46544, n46545, n46546, n46547, n46548, n46549, n46550, n46551, n46552, n46553, n46554, n46555, n46556, n46557, n46558, n46559, n46560, n46561, n46562, n46563, n46564, n46565, n46566, n46567, n46568, n46569, n46570, n46571, n46572, n46573, n46574, n46575, n46576, n46577, n46578, n46579, n46580, n46581, n46582, n46583, n46584, n46585, n46586, n46587, n46588, n46589, n46590, n46591, n46592, n46593, n46594, n46595, n46596, n46597, n46598, n46599, n46600, n46601, n46602, n46603, n46604, n46605, n46606, n46607, n46608, n46609, n46610, n46611, n46612, n46613, n46614, n46615, n46616, n46617, n46618, n46619, n46620, n46621, n46622, n46623, n46624, n46625, n46626, n46627, n46628, n46629, n46630, n46631, n46632, n46633, n46634, n46635, n46636, n46637, n46638, n46639, n46640, n46641, n46642, n46643, n46644, n46645, n46646, n46647, n46648, n46649, n46650, n46651, n46652, n46653, n46654, n46655, n46656, n46657, n46658, n46659, n46660, n46661, n46662, n46663, n46664, n46665, n46666, n46667, n46668, n46669, n46670, n46671, n46672, n46673, n46674, n46675, n46676, n46677, n46678, n46679, n46680, n46681, n46682, n46683, n46684, n46685, n46686, n46687, n46688, n46689, n46690, n46691, n46692, n46693, n46694, n46695, n46696, n46697, n46698, n46699, n46700, n46701, n46702, n46703, n46704, n46705, n46706, n46707, n46708, n46709, n46710, n46711, n46712, n46713, n46714, n46715, n46716, n46717, n46718, n46719, n46720, n46721, n46722, n46723, n46724, n46725, n46726, n46727, n46728, n46729, n46730, n46731, n46732, n46733, n46734, n46735, n46736, n46737, n46738, n46739, n46740, n46741, n46742, n46743, n46744, n46745, n46746, n46747, n46748, n46749, n46750, n46751, n46752, n46753, n46754, n46755, n46756, n46757, n46758, n46759, n46760, n46761, n46762, n46763, n46764, n46765, n46766, n46767, n46768, n46769, n46770, n46771, n46772, n46773, n46774, n46775, n46776, n46777, n46778, n46779, n46780, n46781, n46782, n46783, n46784, n46785, n46786, n46787, n46788, n46789, n46790, n46791, n46792, n46793, n46794, n46795, n46796, n46797, n46798, n46799, n46800, n46801, n46802, n46803, n46804, n46805, n46806, n46807, n46808, n46809, n46810, n46811, n46812, n46813, n46814, n46815, n46816, n46817, n46818, n46819, n46820, n46821, n46822, n46823, n46824, n46825, n46826, n46827, n46828, n46829, n46830, n46831, n46832, n46833, n46834, n46835, n46836, n46837, n46838, n46839, n46840, n46841, n46842, n46843, n46844, n46845, n46846, n46847, n46848, n46849, n46850, n46851, n46852, n46853, n46854, n46855, n46856, n46857, n46858, n46859, n46860, n46861, n46862, n46863, n46864, n46865, n46866, n46867, n46868, n46869, n46870, n46871, n46872, n46873, n46874, n46875, n46876, n46877, n46878, n46879, n46880, n46881, n46882, n46883, n46884, n46885, n46886, n46887, n46888, n46889, n46890, n46891, n46892, n46893, n46894, n46895, n46896, n46897, n46898, n46899, n46900, n46901, n46902, n46903, n46904, n46905, n46906, n46907, n46908, n46909, n46910, n46911, n46912, n46913, n46914, n46915, n46916, n46917, n46918, n46919, n46920, n46921, n46922, n46923, n46924, n46925, n46926, n46927, n46928, n46929, n46930, n46931, n46932, n46933, n46934, n46935, n46936, n46937, n46938, n46939, n46940, n46941, n46942, n46943, n46944, n46945, n46946, n46947, n46948, n46949, n46950, n46951, n46952, n46953, n46954, n46955, n46956, n46957, n46958, n46959, n46960, n46961, n46962, n46963, n46964, n46965, n46966, n46967, n46968, n46969, n46970, n46971, n46972, n46973, n46974, n46975, n46976, n46977, n46978, n46979, n46980, n46981, n46982, n46983, n46984, n46985, n46986, n46987, n46988, n46989, n46990, n46991, n46992, n46993, n46994, n46995, n46996, n46997, n46998, n46999, n47000, n47001, n47002, n47003, n47004, n47005, n47006, n47007, n47008, n47009, n47010, n47011, n47012, n47013, n47014, n47015, n47016, n47017, n47018, n47019, n47020, n47021, n47022, n47023, n47024, n47025, n47026, n47027, n47028, n47029, n47030, n47031, n47032, n47033, n47034, n47035, n47036, n47037, n47038, n47039, n47040, n47041, n47042, n47043, n47044, n47045, n47046, n47047, n47048, n47049, n47050, n47051, n47052, n47053, n47054, n47055, n47056, n47057, n47058, n47059, n47060, n47061, n47062, n47063, n47064, n47065, n47066, n47067, n47068, n47069, n47070, n47071, n47072, n47073, n47074, n47075, n47076, n47077, n47078, n47079, n47080, n47081, n47082, n47083, n47084, n47085, n47086, n47087, n47088, n47089, n47090, n47091, n47092, n47093, n47094, n47095, n47096, n47097, n47098, n47099, n47100, n47101, n47102, n47103, n47104, n47105, n47106, n47107, n47108, n47109, n47110, n47111, n47112, n47113, n47114, n47115, n47116, n47117, n47118, n47119, n47120, n47121, n47122, n47123, n47124, n47125, n47126, n47127, n47128, n47129, n47130, n47131, n47132, n47133, n47134, n47135, n47136, n47137, n47138, n47139, n47140, n47141, n47142, n47143, n47144, n47145, n47146, n47147, n47148, n47149, n47150, n47151, n47152, n47153, n47154, n47155, n47156, n47157, n47158, n47159, n47160, n47161, n47162, n47163, n47164, n47165, n47166, n47167, n47168, n47169, n47170, n47171, n47172, n47173, n47174, n47175, n47176, n47177, n47178, n47179, n47180, n47181, n47182, n47183, n47184, n47185, n47186, n47187, n47188, n47189, n47190, n47191, n47192, n47193, n47194, n47195, n47196, n47197, n47198, n47199, n47200, n47201, n47202, n47203, n47204, n47205, n47206, n47207, n47208, n47209, n47210, n47211, n47212, n47213, n47214, n47215, n47216, n47217, n47218, n47219, n47220, n47221, n47222, n47223, n47224, n47225, n47226, n47227, n47228, n47229, n47230, n47231, n47232, n47233, n47234, n47235, n47236, n47237, n47238, n47239, n47240, n47241, n47242, n47243, n47244, n47245, n47246, n47247, n47248, n47249, n47250, n47251, n47252, n47253, n47254, n47255, n47256, n47257, n47258, n47259, n47260, n47261, n47262, n47263, n47264, n47265, n47266, n47267, n47268, n47269, n47270, n47271, n47272, n47273, n47274, n47275, n47276, n47277, n47278, n47279, n47280, n47281, n47282, n47283, n47284, n47285, n47286, n47287, n47288, n47289, n47290, n47291, n47292, n47293, n47294, n47295, n47296, n47297, n47298, n47299, n47300, n47301, n47302, n47303, n47304, n47305, n47306, n47307, n47308, n47309, n47310, n47311, n47312, n47313, n47314, n47315, n47316, n47317, n47318, n47319, n47320, n47321, n47322, n47323, n47324, n47325, n47326, n47327, n47328, n47329, n47330, n47331, n47332, n47333, n47334, n47335, n47336, n47337, n47338, n47339, n47340, n47341, n47342, n47343, n47344, n47345, n47346, n47347, n47348, n47349, n47350, n47351, n47352, n47353, n47354, n47355, n47356, n47357, n47358, n47359, n47360, n47361, n47362, n47363, n47364, n47365, n47366, n47367, n47368, n47369, n47370, n47371, n47372, n47373, n47374, n47375, n47376, n47377, n47378, n47379, n47380, n47381, n47382, n47383, n47384, n47385, n47386, n47387, n47388, n47389, n47390, n47391, n47392, n47393, n47394, n47395, n47396, n47397, n47398, n47399, n47400, n47401, n47402, n47403, n47404, n47405, n47406, n47407, n47408, n47409, n47410, n47411, n47412, n47413, n47414, n47415, n47416, n47417, n47418, n47419, n47420, n47421, n47422, n47423, n47424, n47425, n47426, n47427, n47428, n47429, n47430, n47431, n47432, n47433, n47434, n47435, n47436, n47437, n47438, n47439, n47440, n47441, n47442, n47443, n47444, n47445, n47446, n47447, n47448, n47449, n47450, n47451, n47452, n47453, n47454, n47455, n47456, n47457, n47458, n47459, n47460, n47461, n47462, n47463, n47464, n47465, n47466, n47467, n47468, n47469, n47470, n47471, n47472, n47473, n47474, n47475, n47476, n47477, n47478, n47479, n47480, n47481, n47482, n47483, n47484, n47485, n47486, n47487, n47488, n47489, n47490, n47491, n47492, n47493, n47494, n47495, n47496, n47497, n47498, n47499, n47500, n47501, n47502, n47503, n47504, n47505, n47506, n47507, n47508, n47509, n47510, n47511, n47512, n47513, n47514, n47515, n47516, n47517, n47518, n47519, n47520, n47521, n47522, n47523, n47524, n47525, n47526, n47527, n47528, n47529, n47530, n47531, n47532, n47533, n47534, n47535, n47536, n47537, n47538, n47539, n47540, n47541, n47542, n47543, n47544, n47545, n47546, n47547, n47548, n47549, n47550, n47551, n47552, n47553, n47554, n47555, n47556, n47557, n47558, n47559, n47560, n47561, n47562, n47563, n47564, n47565, n47566, n47567, n47568, n47569, n47570, n47571, n47572, n47573, n47574, n47575, n47576, n47577, n47578, n47579, n47580, n47581, n47582, n47583, n47584, n47585, n47586, n47587, n47588, n47589, n47590, n47591, n47592, n47593, n47594, n47595, n47596, n47597, n47598, n47599, n47600, n47601, n47602, n47603, n47604, n47605, n47606, n47607, n47608, n47609, n47610, n47611, n47612, n47613, n47614, n47615, n47616, n47617, n47618, n47619, n47620, n47621, n47622, n47623, n47624, n47625, n47626, n47627, n47628, n47629, n47630, n47631, n47632, n47633, n47634, n47635, n47636, n47637, n47638, n47639, n47640, n47641, n47642, n47643, n47644, n47645, n47646, n47647, n47648, n47649, n47650, n47651, n47652, n47653, n47654, n47655, n47656, n47657, n47658, n47659, n47660, n47661, n47662, n47663, n47664, n47665, n47666, n47667, n47668, n47669, n47670, n47671, n47672, n47673, n47674, n47675, n47676, n47677, n47678, n47679, n47680, n47681, n47682, n47683, n47684, n47685, n47686, n47687, n47688, n47689, n47690, n47691, n47692, n47693, n47694, n47695, n47696, n47697, n47698, n47699, n47700, n47701, n47702, n47703, n47704, n47705, n47706, n47707, n47708, n47709, n47710, n47711, n47712, n47713, n47714, n47715, n47716, n47717, n47718, n47719, n47720, n47721, n47722, n47723, n47724, n47725, n47726, n47727, n47728, n47729, n47730, n47731, n47732, n47733, n47734, n47735, n47736, n47737, n47738, n47739, n47740, n47741, n47742, n47743, n47744, n47745, n47746, n47747, n47748, n47749, n47750, n47751, n47752, n47753, n47754, n47755, n47756, n47757, n47758, n47759, n47760, n47761, n47762, n47763, n47764, n47765, n47766, n47767, n47768, n47769, n47770, n47771, n47772, n47773, n47774, n47775, n47776, n47777, n47778, n47779, n47780, n47781, n47782, n47783, n47784, n47785, n47786, n47787, n47788, n47789, n47790, n47791, n47792, n47793, n47794, n47795, n47796, n47797, n47798, n47799, n47800, n47801, n47802, n47803, n47804, n47805, n47806, n47807, n47808, n47809, n47810, n47811, n47812, n47813, n47814, n47815, n47816, n47817, n47818, n47819, n47820, n47821, n47822, n47823, n47824, n47825, n47826, n47827, n47828, n47829, n47830, n47831, n47832, n47833, n47834, n47835, n47836, n47837, n47838, n47839, n47840, n47841, n47842, n47843, n47844, n47845, n47846, n47847, n47848, n47849, n47850, n47851, n47852, n47853, n47854, n47855, n47856, n47857, n47858, n47859, n47860, n47861, n47862, n47863, n47864, n47865, n47866, n47867, n47868, n47869, n47870, n47871, n47872, n47873, n47874, n47875, n47876, n47877, n47878, n47879, n47880, n47881, n47882, n47883, n47884, n47885, n47886, n47887, n47888, n47889, n47890, n47891, n47892, n47893, n47894, n47895, n47896, n47897, n47898, n47899, n47900, n47901, n47902, n47903, n47904, n47905, n47906, n47907, n47908, n47909, n47910, n47911, n47912, n47913, n47914, n47915, n47916, n47917, n47918, n47919, n47920, n47921, n47922, n47923, n47924, n47925, n47926, n47927, n47928, n47929, n47930, n47931, n47932, n47933, n47934, n47935, n47936, n47937, n47938, n47939, n47940, n47941, n47942, n47943, n47944, n47945, n47946, n47947, n47948, n47949, n47950, n47951, n47952, n47953, n47954, n47955, n47956, n47957, n47958, n47959, n47960, n47961, n47962, n47963, n47964, n47965, n47966, n47967, n47968, n47969, n47970, n47971, n47972, n47973, n47974, n47975, n47976, n47977, n47978, n47979, n47980, n47981, n47982, n47983, n47984, n47985, n47986, n47987, n47988, n47989, n47990, n47991, n47992, n47993, n47994, n47995, n47996, n47997, n47998, n47999, n48000, n48001, n48002, n48003, n48004, n48005, n48006, n48007, n48008, n48009, n48010, n48011, n48012, n48013, n48014, n48015, n48016, n48017, n48018, n48019, n48020, n48021, n48022, n48023, n48024, n48025, n48026, n48027, n48028, n48029, n48030, n48031, n48032, n48033, n48034, n48035, n48036, n48037, n48038, n48039, n48040, n48041, n48042, n48043, n48044, n48045, n48046, n48047, n48048, n48049, n48050, n48051, n48052, n48053, n48054, n48055, n48056, n48057, n48058, n48059, n48060, n48061, n48062, n48063, n48064, n48065, n48066, n48067, n48068, n48069, n48070, n48071, n48072, n48073, n48074, n48075, n48076, n48077, n48078, n48079, n48080, n48081, n48082, n48083, n48084, n48085, n48086, n48087, n48088, n48089, n48090, n48091, n48092, n48093, n48094, n48095, n48096, n48097, n48098, n48099, n48100, n48101, n48102, n48103, n48104, n48105, n48106, n48107, n48108, n48109, n48110, n48111, n48112, n48113, n48114, n48115, n48116, n48117, n48118, n48119, n48120, n48121, n48122, n48123, n48124, n48125, n48126, n48127, n48128, n48129, n48130, n48131, n48132, n48133, n48134, n48135, n48136, n48137, n48138, n48139, n48140, n48141, n48142, n48143, n48144, n48145, n48146, n48147, n48148, n48149, n48150, n48151, n48152, n48153, n48154, n48155, n48156, n48157, n48158, n48159, n48160, n48161, n48162, n48163, n48164, n48165, n48166, n48167, n48168, n48169, n48170, n48171, n48172, n48173, n48174, n48175, n48176, n48177, n48178, n48179, n48180, n48181, n48182, n48183, n48184, n48185, n48186, n48187, n48188, n48189, n48190, n48191, n48192, n48193, n48194, n48195, n48196, n48197, n48198, n48199, n48200, n48201, n48202, n48203, n48204, n48205, n48206, n48207, n48208, n48209, n48210, n48211, n48212, n48213, n48214, n48215, n48216, n48217, n48218, n48219, n48220, n48221, n48222, n48223, n48224, n48225, n48226, n48227, n48228, n48229, n48230, n48231, n48232, n48233, n48234, n48235, n48236, n48237, n48238, n48239, n48240, n48241, n48242, n48243, n48244, n48245, n48246, n48247, n48248, n48249, n48250, n48251, n48252, n48253, n48254, n48255, n48256, n48257, n48258, n48259, n48260, n48261, n48262, n48263, n48264, n48265, n48266, n48267, n48268, n48269, n48270, n48271, n48272, n48273, n48274, n48275, n48276, n48277, n48278, n48279, n48280, n48281, n48282, n48283, n48284, n48285, n48286, n48287, n48288, n48289, n48290, n48291, n48292, n48293, n48294, n48295, n48296, n48297, n48298, n48299, n48300, n48301, n48302, n48303, n48304, n48305, n48306, n48307, n48308, n48309, n48310, n48311, n48312, n48313, n48314, n48315, n48316, n48317, n48318, n48319, n48320, n48321, n48322, n48323, n48324, n48325, n48326, n48327, n48328, n48329, n48330, n48331, n48332, n48333, n48334, n48335, n48336, n48337, n48338, n48339, n48340, n48341, n48342, n48343, n48344, n48345, n48346, n48347, n48348, n48349, n48350, n48351, n48352, n48353, n48354, n48355, n48356, n48357, n48358, n48359, n48360, n48361, n48362, n48363, n48364, n48365, n48366, n48367, n48368, n48369, n48370, n48371, n48372, n48373, n48374, n48375, n48376, n48377, n48378, n48379, n48380, n48381, n48382, n48383, n48384, n48385, n48386, n48387, n48388, n48389, n48390, n48391, n48392, n48393, n48394, n48395, n48396, n48397, n48398, n48399, n48400, n48401, n48402, n48403, n48404, n48405, n48406, n48407, n48408, n48409, n48410, n48411, n48412, n48413, n48414, n48415, n48416, n48417, n48418, n48419, n48420, n48421, n48422, n48423, n48424, n48425, n48426, n48427, n48428, n48429, n48430, n48431, n48432, n48433, n48434, n48435, n48436, n48437, n48438, n48439, n48440, n48441, n48442, n48443, n48444, n48445, n48446, n48447, n48448, n48449, n48450, n48451, n48452, n48453, n48454, n48455, n48456, n48457, n48458, n48459, n48460, n48461, n48462, n48463, n48464, n48465, n48466, n48467, n48468, n48469, n48470, n48471, n48472, n48473, n48474, n48475, n48476, n48477, n48478, n48479, n48480, n48481, n48482, n48483, n48484, n48485, n48486, n48487, n48488, n48489, n48490, n48491, n48492, n48493, n48494, n48495, n48496, n48497, n48498, n48499, n48500, n48501, n48502, n48503, n48504, n48505, n48506, n48507, n48508, n48509, n48510, n48511, n48512, n48513, n48514, n48515, n48516, n48517, n48518, n48519, n48520, n48521, n48522, n48523, n48524, n48525, n48526, n48527, n48528, n48529, n48530, n48531, n48532, n48533, n48534, n48535, n48536, n48537, n48538, n48539, n48540, n48541, n48542, n48543, n48544, n48545, n48546, n48547, n48548, n48549, n48550, n48551, n48552, n48553, n48554, n48555, n48556, n48557, n48558, n48559, n48560, n48561, n48562, n48563, n48564, n48565, n48566, n48567, n48568, n48569, n48570, n48571, n48572, n48573, n48574, n48575, n48576, n48577, n48578, n48579, n48580, n48581, n48582, n48583, n48584, n48585, n48586, n48587, n48588, n48589, n48590, n48591, n48592, n48593, n48594, n48595, n48596, n48597, n48598, n48599, n48600, n48601, n48602, n48603, n48604, n48605, n48606, n48607, n48608, n48609, n48610, n48611, n48612, n48613, n48614, n48615, n48616, n48617, n48618, n48619, n48620, n48621, n48622, n48623, n48624, n48625, n48626, n48627, n48628, n48629, n48630, n48631, n48632, n48633, n48634, n48635, n48636, n48637, n48638, n48639, n48640, n48641, n48642, n48643, n48644, n48645, n48646, n48647, n48648, n48649, n48650, n48651, n48652, n48653, n48654, n48655, n48656, n48657, n48658, n48659, n48660, n48661, n48662, n48663, n48664, n48665, n48666, n48667, n48668, n48669, n48670, n48671, n48672, n48673, n48674, n48675, n48676, n48677, n48678, n48679, n48680, n48681, n48682, n48683, n48684, n48685, n48686, n48687, n48688, n48689, n48690, n48691, n48692, n48693, n48694, n48695, n48696, n48697, n48698, n48699, n48700, n48701, n48702, n48703, n48704, n48705, n48706, n48707, n48708, n48709, n48710, n48711, n48712, n48713, n48714, n48715, n48716, n48717, n48718, n48719, n48720, n48721, n48722, n48723, n48724, n48725, n48726, n48727, n48728, n48729, n48730, n48731, n48732, n48733, n48734, n48735, n48736, n48737, n48738, n48739, n48740, n48741, n48742, n48743, n48744, n48745, n48746, n48747, n48748, n48749, n48750, n48751, n48752, n48753, n48754, n48755, n48756, n48757, n48758, n48759, n48760, n48761, n48762, n48763, n48764, n48765, n48766, n48767, n48768, n48769, n48770, n48771, n48772, n48773, n48774, n48775, n48776, n48777, n48778, n48779, n48780, n48781, n48782, n48783, n48784, n48785, n48786, n48787, n48788, n48789, n48790, n48791, n48792, n48793, n48794, n48795, n48796, n48797, n48798, n48799, n48800, n48801, n48802, n48803, n48804, n48805, n48806, n48807, n48808, n48809, n48810, n48811, n48812, n48813, n48814, n48815, n48816, n48817, n48818, n48819, n48820, n48821, n48822, n48823, n48824, n48825, n48826, n48827, n48828, n48829, n48830, n48831, n48832, n48833, n48834, n48835, n48836, n48837, n48838, n48839, n48840, n48841, n48842, n48843, n48844, n48845, n48846, n48847, n48848, n48849, n48850, n48851, n48852, n48853, n48854, n48855, n48856, n48857, n48858, n48859, n48860, n48861, n48862, n48863, n48864, n48865, n48866, n48867, n48868, n48869, n48870, n48871, n48872, n48873, n48874, n48875, n48876, n48877, n48878, n48879, n48880, n48881, n48882, n48883, n48884, n48885, n48886, n48887, n48888, n48889, n48890, n48891, n48892, n48893, n48894, n48895, n48896, n48897, n48898, n48899, n48900, n48901, n48902, n48903, n48904, n48905, n48906, n48907, n48908, n48909, n48910, n48911, n48912, n48913, n48914, n48915, n48916, n48917, n48918, n48919, n48920, n48921, n48922, n48923, n48924, n48925, n48926, n48927, n48928, n48929, n48930, n48931, n48932, n48933, n48934, n48935, n48936, n48937, n48938, n48939, n48940, n48941, n48942, n48943, n48944, n48945, n48946, n48947, n48948, n48949, n48950, n48951, n48952, n48953, n48954, n48955, n48956, n48957, n48958, n48959, n48960, n48961, n48962, n48963, n48964, n48965, n48966, n48967, n48968, n48969, n48970, n48971, n48972, n48973, n48974, n48975, n48976, n48977, n48978, n48979, n48980, n48981, n48982, n48983, n48984, n48985, n48986, n48987, n48988, n48989, n48990, n48991, n48992, n48993, n48994, n48995, n48996, n48997, n48998, n48999, n49000, n49001, n49002, n49003, n49004, n49005, n49006, n49007, n49008, n49009, n49010, n49011, n49012, n49013, n49014, n49015, n49016, n49017, n49018, n49019, n49020, n49021, n49022, n49023, n49024, n49025, n49026, n49027, n49028, n49029, n49030, n49031, n49032, n49033, n49034, n49035, n49036, n49037, n49038, n49039, n49040, n49041, n49042, n49043, n49044, n49045, n49046, n49047, n49048, n49049, n49050, n49051, n49052, n49053, n49054, n49055, n49056, n49057, n49058, n49059, n49060, n49061, n49062, n49063, n49064, n49065, n49066, n49067, n49068, n49069, n49070, n49071, n49072, n49073, n49074, n49075, n49076, n49077, n49078, n49079, n49080, n49081, n49082, n49083, n49084, n49085, n49086, n49087, n49088, n49089, n49090, n49091, n49092, n49093, n49094, n49095, n49096, n49097, n49098, n49099, n49100, n49101, n49102, n49103, n49104, n49105, n49106, n49107, n49108, n49109, n49110, n49111, n49112, n49113, n49114, n49115, n49116, n49117, n49118, n49119, n49120, n49121, n49122, n49123, n49124, n49125, n49126, n49127, n49128, n49129, n49130, n49131, n49132, n49133, n49134, n49135, n49136, n49137, n49138, n49139, n49140, n49141, n49142, n49143, n49144, n49145, n49146, n49147, n49148, n49149, n49150, n49151, n49152, n49153, n49154, n49155, n49156, n49157, n49158, n49159, n49160, n49161, n49162, n49163, n49164, n49165, n49166, n49167, n49168, n49169, n49170, n49171, n49172, n49173, n49174, n49175, n49176, n49177, n49178, n49179, n49180, n49181, n49182, n49183, n49184, n49185, n49186, n49187, n49188, n49189, n49190, n49191, n49192, n49193, n49194, n49195, n49196, n49197, n49198, n49199, n49200, n49201, n49202, n49203, n49204, n49205, n49206, n49207, n49208, n49209, n49210, n49211, n49212, n49213, n49214, n49215, n49216, n49217, n49218, n49219, n49220, n49221, n49222, n49223, n49224, n49225, n49226, n49227, n49228, n49229, n49230, n49231, n49232, n49233, n49234, n49235, n49236, n49237, n49238, n49239, n49240, n49241, n49242, n49243, n49244, n49245, n49246, n49247, n49248, n49249, n49250, n49251, n49252, n49253, n49254, n49255, n49256, n49257, n49258, n49259, n49260, n49261, n49262, n49263, n49264, n49265, n49266, n49267, n49268, n49269, n49270, n49271, n49272, n49273, n49274, n49275, n49276, n49277, n49278, n49279, n49280, n49281, n49282, n49283, n49284, n49285, n49286, n49287, n49288, n49289, n49290, n49291, n49292, n49293, n49294, n49295, n49296, n49297, n49298, n49299, n49300, n49301, n49302, n49303, n49304, n49305, n49306, n49307, n49308, n49309, n49310, n49311, n49312, n49313, n49314, n49315, n49316, n49317, n49318, n49319, n49320, n49321, n49322, n49323, n49324, n49325, n49326, n49327, n49328, n49329, n49330, n49331, n49332, n49333, n49334, n49335, n49336, n49337, n49338, n49339, n49340, n49341, n49342, n49343, n49344, n49345, n49346, n49347, n49348, n49349, n49350, n49351, n49352, n49353, n49354, n49355, n49356, n49357, n49358, n49359, n49360, n49361, n49362, n49363, n49364, n49365, n49366, n49367, n49368, n49369, n49370, n49371, n49372, n49373, n49374, n49375, n49376, n49377, n49378, n49379, n49380, n49381, n49382, n49383, n49384, n49385, n49386, n49387, n49388, n49389, n49390, n49391, n49392, n49393, n49394, n49395, n49396, n49397, n49398, n49399, n49400, n49401, n49402, n49403, n49404, n49405, n49406, n49407, n49408, n49409, n49410, n49411, n49412, n49413, n49414, n49415, n49416, n49417, n49418, n49419, n49420, n49421, n49422, n49423, n49424, n49425, n49426, n49427, n49428, n49429, n49430, n49431, n49432, n49433, n49434, n49435, n49436, n49437, n49438, n49439, n49440, n49441, n49442, n49443, n49444, n49445, n49446, n49447, n49448, n49449, n49450, n49451, n49452, n49453, n49454, n49455, n49456, n49457, n49458, n49459, n49460, n49461, n49462, n49463, n49464, n49465, n49466, n49467, n49468, n49469, n49470, n49471, n49472, n49473, n49474, n49475, n49476, n49477, n49478, n49479, n49480, n49481, n49482, n49483, n49484, n49485, n49486, n49487, n49488, n49489, n49490, n49491, n49492, n49493, n49494, n49495, n49496, n49497, n49498, n49499, n49500, n49501, n49502, n49503, n49504, n49505, n49506, n49507, n49508, n49509, n49510, n49511, n49512, n49513, n49514, n49515, n49516, n49517, n49518, n49519, n49520, n49521, n49522, n49523, n49524, n49525, n49526, n49527, n49528, n49529, n49530, n49531, n49532, n49533, n49534, n49535, n49536, n49537, n49538, n49539, n49540, n49541, n49542, n49543, n49544, n49545, n49546, n49547, n49548, n49549, n49550, n49551, n49552, n49553, n49554, n49555, n49556, n49557, n49558, n49559, n49560, n49561, n49562, n49563, n49564, n49565, n49566, n49567, n49568, n49569, n49570, n49571, n49572, n49573, n49574, n49575, n49576, n49577, n49578, n49579, n49580, n49581, n49582, n49583, n49584, n49585, n49586, n49587, n49588, n49589, n49590, n49591, n49592, n49593, n49594, n49595, n49596, n49597, n49598, n49599, n49600, n49601, n49602, n49603, n49604, n49605, n49606, n49607, n49608, n49609, n49610, n49611, n49612, n49613, n49614, n49615, n49616, n49617, n49618, n49619, n49620, n49621, n49622, n49623, n49624, n49625, n49626, n49627, n49628, n49629, n49630, n49631, n49632, n49633, n49634, n49635, n49636, n49637, n49638, n49639, n49640, n49641, n49642, n49643, n49644, n49645, n49646, n49647, n49648, n49649, n49650, n49651, n49652, n49653, n49654, n49655, n49656, n49657, n49658, n49659, n49660, n49661, n49662, n49663, n49664, n49665, n49666, n49667, n49668, n49669, n49670, n49671, n49672, n49673, n49674, n49675, n49676, n49677, n49678, n49679, n49680, n49681, n49682, n49683, n49684, n49685, n49686, n49687, n49688, n49689, n49690, n49691, n49692, n49693, n49694, n49695, n49696, n49697, n49698, n49699, n49700, n49701, n49702, n49703, n49704, n49705, n49706, n49707, n49708, n49709, n49710, n49711, n49712, n49713, n49714, n49715, n49716, n49717, n49718, n49719, n49720, n49721, n49722, n49723, n49724, n49725, n49726, n49727, n49728, n49729, n49730, n49731, n49732, n49733, n49734, n49735, n49736, n49737, n49738, n49739, n49740, n49741, n49742, n49743, n49744, n49745, n49746, n49747, n49748, n49749, n49750, n49751, n49752, n49753, n49754, n49755, n49756, n49757, n49758, n49759, n49760, n49761, n49762, n49763, n49764, n49765, n49766, n49767, n49768, n49769, n49770, n49771, n49772, n49773, n49774, n49775, n49776, n49777, n49778, n49779, n49780, n49781, n49782, n49783, n49784, n49785, n49786, n49787, n49788, n49789, n49790, n49791, n49792, n49793, n49794, n49795, n49796, n49797, n49798, n49799, n49800, n49801, n49802, n49803, n49804, n49805, n49806, n49807, n49808, n49809, n49810, n49811, n49812, n49813, n49814, n49815, n49816, n49817, n49818, n49819, n49820, n49821, n49822, n49823, n49824, n49825, n49826, n49827, n49828, n49829, n49830, n49831, n49832, n49833, n49834, n49835, n49836, n49837, n49838, n49839, n49840, n49841, n49842, n49843, n49844, n49845, n49846, n49847, n49848, n49849, n49850, n49851, n49852, n49853, n49854, n49855, n49856, n49857, n49858, n49859, n49860, n49861, n49862, n49863, n49864, n49865, n49866, n49867, n49868, n49869, n49870, n49871, n49872, n49873, n49874, n49875, n49876, n49877, n49878, n49879, n49880, n49881, n49882, n49883, n49884, n49885, n49886, n49887, n49888, n49889, n49890, n49891, n49892, n49893, n49894, n49895, n49896, n49897, n49898, n49899, n49900, n49901, n49902, n49903, n49904, n49905, n49906, n49907, n49908, n49909, n49910, n49911, n49912, n49913, n49914, n49915, n49916, n49917, n49918, n49919, n49920, n49921, n49922, n49923, n49924, n49925, n49926, n49927, n49928, n49929, n49930, n49931, n49932, n49933, n49934, n49935, n49936, n49937, n49938, n49939, n49940, n49941, n49942, n49943, n49944, n49945, n49946, n49947, n49948, n49949, n49950, n49951, n49952, n49953, n49954, n49955, n49956, n49957, n49958, n49959, n49960, n49961, n49962, n49963, n49964, n49965, n49966, n49967, n49968, n49969, n49970, n49971, n49972, n49973, n49974, n49975, n49976, n49977, n49978, n49979, n49980, n49981, n49982, n49983, n49984, n49985, n49986, n49987, n49988, n49989, n49990, n49991, n49992, n49993, n49994, n49995, n49996, n49997, n49998, n49999, n50000, n50001, n50002, n50003, n50004, n50005, n50006, n50007, n50008, n50009, n50010, n50011, n50012, n50013, n50014, n50015, n50016, n50017, n50018, n50019, n50020, n50021, n50022, n50023, n50024, n50025, n50026, n50027, n50028, n50029, n50030, n50031, n50032, n50033, n50034, n50035, n50036, n50037, n50038, n50039, n50040, n50041, n50042, n50043, n50044, n50045, n50046, n50047, n50048, n50049, n50050, n50051, n50052, n50053, n50054, n50055, n50056, n50057, n50058, n50059, n50060, n50061, n50062, n50063, n50064, n50065, n50066, n50067, n50068, n50069, n50070, n50071, n50072, n50073, n50074, n50075, n50076, n50077, n50078, n50079, n50080, n50081, n50082, n50083, n50084, n50085, n50086, n50087, n50088, n50089, n50090, n50091, n50092, n50093, n50094, n50095, n50096, n50097, n50098, n50099, n50100, n50101, n50102, n50103, n50104, n50105, n50106, n50107, n50108, n50109, n50110, n50111, n50112, n50113, n50114, n50115, n50116, n50117, n50118, n50119, n50120, n50121, n50122, n50123, n50124, n50125, n50126, n50127, n50128, n50129, n50130, n50131, n50132, n50133, n50134, n50135, n50136, n50137, n50138, n50139, n50140, n50141, n50142, n50143, n50144, n50145, n50146, n50147, n50148, n50149, n50150, n50151, n50152, n50153, n50154, n50155, n50156, n50157, n50158, n50159, n50160, n50161, n50162, n50163, n50164, n50165, n50166, n50167, n50168, n50169, n50170, n50171, n50172, n50173, n50174, n50175, n50176, n50177, n50178, n50179, n50180, n50181, n50182, n50183, n50184, n50185, n50186, n50187, n50188, n50189, n50190, n50191, n50192, n50193, n50194, n50195, n50196, n50197, n50198, n50199, n50200, n50201, n50202, n50203, n50204, n50205, n50206, n50207, n50208, n50209, n50210, n50211, n50212, n50213, n50214, n50215, n50216, n50217, n50218, n50219, n50220, n50221, n50222, n50223, n50224, n50225, n50226, n50227, n50228, n50229, n50230, n50231, n50232, n50233, n50234, n50235, n50236, n50237, n50238, n50239, n50240, n50241, n50242, n50243, n50244, n50245, n50246, n50247, n50248, n50249, n50250, n50251, n50252, n50253, n50254, n50255, n50256, n50257, n50258, n50259, n50260, n50261, n50262, n50263, n50264, n50265, n50266, n50267, n50268, n50269, n50270, n50271, n50272, n50273, n50274, n50275, n50276, n50277, n50278, n50279, n50280, n50281, n50282, n50283, n50284, n50285, n50286, n50287, n50288, n50289, n50290, n50291, n50292, n50293, n50294, n50295, n50296, n50297, n50298, n50299, n50300, n50301, n50302, n50303, n50304, n50305, n50306, n50307, n50308, n50309, n50310, n50311, n50312, n50313, n50314, n50315, n50316, n50317, n50318, n50319, n50320, n50321, n50322, n50323, n50324, n50325, n50326, n50327, n50328, n50329, n50330, n50331, n50332, n50333, n50334, n50335, n50336, n50337, n50338, n50339, n50340, n50341, n50342, n50343, n50344, n50345, n50346, n50347, n50348, n50349, n50350, n50351, n50352, n50353, n50354, n50355, n50356, n50357, n50358, n50359, n50360, n50361, n50362, n50363, n50364, n50365, n50366, n50367, n50368, n50369, n50370, n50371, n50372, n50373, n50374, n50375, n50376, n50377, n50378, n50379, n50380, n50381, n50382, n50383, n50384, n50385, n50386, n50387, n50388, n50389, n50390, n50391, n50392, n50393, n50394, n50395, n50396, n50397, n50398, n50399, n50400, n50401, n50402, n50403, n50404, n50405, n50406, n50407, n50408, n50409, n50410, n50411, n50412, n50413, n50414, n50415, n50416, n50417, n50418, n50419, n50420, n50421, n50422, n50423, n50424, n50425, n50426, n50427, n50428, n50429, n50430, n50431, n50432, n50433, n50434, n50435, n50436, n50437, n50438, n50439, n50440, n50441, n50442, n50443, n50444, n50445, n50446, n50447, n50448, n50449, n50450, n50451, n50452, n50453, n50454, n50455, n50456, n50457, n50458, n50459, n50460, n50461, n50462, n50463, n50464, n50465, n50466, n50467, n50468, n50469, n50470, n50471, n50472, n50473, n50474, n50475, n50476, n50477, n50478, n50479, n50480, n50481, n50482, n50483, n50484, n50485, n50486, n50487, n50488, n50489, n50490, n50491, n50492, n50493, n50494, n50495, n50496, n50497, n50498, n50499, n50500, n50501, n50502, n50503, n50504, n50505, n50506, n50507, n50508, n50509, n50510, n50511, n50512, n50513, n50514, n50515, n50516, n50517, n50518, n50519, n50520, n50521, n50522, n50523, n50524, n50525, n50526, n50527, n50528, n50529, n50530, n50531, n50532, n50533, n50534, n50535, n50536, n50537, n50538, n50539, n50540, n50541, n50542, n50543, n50544, n50545, n50546, n50547, n50548, n50549, n50550, n50551, n50552, n50553, n50554, n50555, n50556, n50557, n50558, n50559, n50560, n50561, n50562, n50563, n50564, n50565, n50566, n50567, n50568, n50569, n50570, n50571, n50572, n50573, n50574, n50575, n50576, n50577, n50578, n50579, n50580, n50581, n50582, n50583, n50584, n50585, n50586, n50587, n50588, n50589, n50590, n50591, n50592, n50593, n50594, n50595, n50596, n50597, n50598, n50599, n50600, n50601, n50602, n50603, n50604, n50605, n50606, n50607, n50608, n50609, n50610, n50611, n50612, n50613, n50614, n50615, n50616, n50617, n50618, n50619, n50620, n50621, n50622, n50623, n50624, n50625, n50626, n50627, n50628, n50629, n50630, n50631, n50632, n50633, n50634, n50635, n50636, n50637, n50638, n50639, n50640, n50641, n50642, n50643, n50644, n50645, n50646, n50647, n50648, n50649, n50650, n50651, n50652, n50653, n50654, n50655, n50656, n50657, n50658, n50659, n50660, n50661, n50662, n50663, n50664, n50665, n50666, n50667, n50668, n50669, n50670, n50671, n50672, n50673, n50674, n50675, n50676, n50677, n50678, n50679, n50680, n50681, n50682, n50683, n50684, n50685, n50686, n50687, n50688, n50689, n50690, n50691, n50692, n50693, n50694, n50695, n50696, n50697, n50698, n50699, n50700, n50701, n50702, n50703, n50704, n50705, n50706, n50707, n50708, n50709, n50710, n50711, n50712, n50713, n50714, n50715, n50716, n50717, n50718, n50719, n50720, n50721, n50722, n50723, n50724, n50725, n50726, n50727, n50728, n50729, n50730, n50731, n50732, n50733, n50734, n50735, n50736, n50737, n50738, n50739, n50740, n50741, n50742, n50743, n50744, n50745, n50746, n50747, n50748, n50749, n50750, n50751, n50752, n50753, n50754, n50755, n50756, n50757, n50758, n50759, n50760, n50761, n50762, n50763, n50764, n50765, n50766, n50767, n50768, n50769, n50770, n50771, n50772, n50773, n50774, n50775, n50776, n50777, n50778, n50779, n50780, n50781, n50782, n50783, n50784, n50785, n50786, n50787, n50788, n50789, n50790, n50791, n50792, n50793, n50794, n50795, n50796, n50797, n50798, n50799, n50800, n50801, n50802, n50803, n50804, n50805, n50806, n50807, n50808, n50809, n50810, n50811, n50812, n50813, n50814, n50815, n50816, n50817, n50818, n50819, n50820, n50821, n50822, n50823, n50824, n50825, n50826, n50827, n50828, n50829, n50830, n50831, n50832, n50833, n50834, n50835, n50836, n50837, n50838, n50839, n50840, n50841, n50842, n50843, n50844, n50845, n50846, n50847, n50848, n50849, n50850, n50851, n50852, n50853, n50854, n50855, n50856, n50857, n50858, n50859, n50860, n50861, n50862, n50863, n50864, n50865, n50866, n50867, n50868, n50869, n50870, n50871, n50872, n50873, n50874, n50875, n50876, n50877, n50878, n50879, n50880, n50881, n50882, n50883, n50884, n50885, n50886, n50887, n50888, n50889, n50890, n50891, n50892, n50893, n50894, n50895, n50896, n50897, n50898, n50899, n50900, n50901, n50902, n50903, n50904, n50905, n50906, n50907, n50908, n50909, n50910, n50911, n50912, n50913, n50914, n50915, n50916, n50917, n50918, n50919, n50920, n50921, n50922, n50923, n50924, n50925, n50926, n50927, n50928, n50929, n50930, n50931, n50932, n50933, n50934, n50935, n50936, n50937, n50938, n50939, n50940, n50941, n50942, n50943, n50944, n50945, n50946, n50947, n50948, n50949, n50950, n50951, n50952, n50953, n50954, n50955, n50956, n50957, n50958, n50959, n50960, n50961, n50962, n50963, n50964, n50965, n50966, n50967, n50968, n50969, n50970, n50971, n50972, n50973, n50974, n50975, n50976, n50977, n50978, n50979, n50980, n50981, n50982, n50983, n50984, n50985, n50986, n50987, n50988, n50989, n50990, n50991, n50992, n50993, n50994, n50995, n50996, n50997, n50998, n50999, n51000, n51001, n51002, n51003, n51004, n51005, n51006, n51007, n51008, n51009, n51010, n51011, n51012, n51013, n51014, n51015, n51016, n51017, n51018, n51019, n51020, n51021, n51022, n51023, n51024, n51025, n51026, n51027, n51028, n51029, n51030, n51031, n51032, n51033, n51034, n51035, n51036, n51037, n51038, n51039, n51040, n51041, n51042, n51043, n51044, n51045, n51046, n51047, n51048, n51049, n51050, n51051, n51052, n51053, n51054, n51055, n51056, n51057, n51058, n51059, n51060, n51061, n51062, n51063, n51064, n51065, n51066, n51067, n51068, n51069, n51070, n51071, n51072, n51073, n51074, n51075, n51076, n51077, n51078, n51079, n51080, n51081, n51082, n51083, n51084, n51085, n51086, n51087, n51088, n51089, n51090, n51091, n51092, n51093, n51094, n51095, n51096, n51097, n51098, n51099, n51100, n51101, n51102, n51103, n51104, n51105, n51106, n51107, n51108, n51109, n51110, n51111, n51112, n51113, n51114, n51115, n51116, n51117, n51118, n51119, n51120, n51121, n51122, n51123, n51124, n51125, n51126, n51127, n51128, n51129, n51130, n51131, n51132, n51133, n51134, n51135, n51136, n51137, n51138, n51139, n51140, n51141, n51142, n51143, n51144, n51145, n51146, n51147, n51148, n51149, n51150, n51151, n51152, n51153, n51154, n51155, n51156, n51157, n51158, n51159, n51160, n51161, n51162, n51163, n51164, n51165, n51166, n51167, n51168, n51169, n51170, n51171, n51172, n51173, n51174, n51175, n51176, n51177, n51178, n51179, n51180, n51181, n51182, n51183, n51184, n51185, n51186, n51187, n51188, n51189, n51190, n51191, n51192, n51193, n51194, n51195, n51196, n51197, n51198, n51199, n51200, n51201, n51202, n51203, n51204, n51205, n51206, n51207, n51208, n51209, n51210, n51211, n51212, n51213, n51214, n51215, n51216, n51217, n51218, n51219, n51220, n51221, n51222, n51223, n51224, n51225, n51226, n51227, n51228, n51229, n51230, n51231, n51232, n51233, n51234, n51235, n51236, n51237, n51238, n51239, n51240, n51241, n51242, n51243, n51244, n51245, n51246, n51247, n51248, n51249, n51250, n51251, n51252, n51253, n51254, n51255, n51256, n51257, n51258, n51259, n51260, n51261, n51262, n51263, n51264, n51265, n51266, n51267, n51268, n51269, n51270, n51271, n51272, n51273, n51274, n51275, n51276, n51277, n51278, n51279, n51280, n51281, n51282, n51283, n51284, n51285, n51286, n51287, n51288, n51289, n51290, n51291, n51292, n51293, n51294, n51295, n51296, n51297, n51298, n51299, n51300, n51301, n51302, n51303, n51304, n51305, n51306, n51307, n51308, n51309, n51310, n51311, n51312, n51313, n51314, n51315, n51316, n51317, n51318, n51319, n51320, n51321, n51322, n51323, n51324, n51325, n51326, n51327, n51328, n51329, n51330, n51331, n51332, n51333, n51334, n51335, n51336, n51337, n51338, n51339, n51340, n51341, n51342, n51343, n51344, n51345, n51346, n51347, n51348, n51349, n51350, n51351, n51352, n51353, n51354, n51355, n51356, n51357, n51358, n51359, n51360, n51361, n51362, n51363, n51364, n51365, n51366, n51367, n51368, n51369, n51370, n51371, n51372, n51373, n51374, n51375, n51376, n51377, n51378, n51379, n51380, n51381, n51382, n51383, n51384, n51385, n51386, n51387, n51388, n51389, n51390, n51391, n51392, n51393, n51394, n51395, n51396, n51397, n51398, n51399, n51400, n51401, n51402, n51403, n51404, n51405, n51406, n51407, n51408, n51409, n51410, n51411, n51412, n51413, n51414, n51415, n51416, n51417, n51418, n51419, n51420, n51421, n51422, n51423, n51424, n51425, n51426, n51427, n51428, n51429, n51430, n51431, n51432, n51433, n51434, n51435, n51436, n51437, n51438, n51439, n51440, n51441, n51442, n51443, n51444, n51445, n51446, n51447, n51448, n51449, n51450, n51451, n51452, n51453, n51454, n51455, n51456, n51457, n51458, n51459, n51460, n51461, n51462, n51463, n51464, n51465, n51466, n51467, n51468, n51469, n51470, n51471, n51472, n51473, n51474, n51475, n51476, n51477, n51478, n51479, n51480, n51481, n51482, n51483, n51484, n51485, n51486, n51487, n51488, n51489, n51490, n51491, n51492, n51493, n51494, n51495, n51496, n51497, n51498, n51499, n51500, n51501, n51502, n51503, n51504, n51505, n51506, n51507, n51508, n51509, n51510, n51511, n51512, n51513, n51514, n51515, n51516, n51517, n51518, n51519, n51520, n51521, n51522, n51523, n51524, n51525, n51526, n51527, n51528, n51529, n51530, n51531, n51532, n51533, n51534, n51535, n51536, n51537, n51538, n51539, n51540, n51541, n51542, n51543, n51544, n51545, n51546, n51547, n51548, n51549, n51550, n51551, n51552, n51553, n51554, n51555, n51556, n51557, n51558, n51559, n51560, n51561, n51562, n51563, n51564, n51565, n51566, n51567, n51568, n51569, n51570, n51571, n51572, n51573, n51574, n51575, n51576, n51577, n51578, n51579, n51580, n51581, n51582, n51583, n51584, n51585, n51586, n51587, n51588, n51589, n51590, n51591, n51592, n51593, n51594, n51595, n51596, n51597, n51598, n51599, n51600, n51601, n51602, n51603, n51604, n51605, n51606, n51607, n51608, n51609, n51610, n51611, n51612, n51613, n51614, n51615, n51616, n51617, n51618, n51619, n51620, n51621, n51622, n51623, n51624, n51625, n51626, n51627, n51628, n51629, n51630, n51631, n51632, n51633, n51634, n51635, n51636, n51637, n51638, n51639, n51640, n51641, n51642, n51643, n51644, n51645, n51646, n51647, n51648, n51649, n51650, n51651, n51652, n51653, n51654, n51655, n51656, n51657, n51658, n51659, n51660, n51661, n51662, n51663, n51664, n51665, n51666, n51667, n51668, n51669, n51670, n51671, n51672, n51673, n51674, n51675, n51676, n51677, n51678, n51679, n51680, n51681, n51682, n51683, n51684, n51685, n51686, n51687, n51688, n51689, n51690, n51691, n51692, n51693, n51694, n51695, n51696, n51697, n51698, n51699, n51700, n51701, n51702, n51703, n51704, n51705, n51706, n51707, n51708, n51709, n51710, n51711, n51712, n51713, n51714, n51715, n51716, n51717, n51718, n51719, n51720, n51721, n51722, n51723, n51724, n51725, n51726, n51727, n51728, n51729, n51730, n51731, n51732, n51733, n51734, n51735, n51736, n51737, n51738, n51739, n51740, n51741, n51742, n51743, n51744, n51745, n51746, n51747, n51748, n51749, n51750, n51751, n51752, n51753, n51754, n51755, n51756, n51757, n51758, n51759, n51760, n51761, n51762, n51763, n51764, n51765, n51766, n51767, n51768, n51769, n51770, n51771, n51772, n51773, n51774, n51775, n51776, n51777, n51778, n51779, n51780, n51781, n51782, n51783, n51784, n51785, n51786, n51787, n51788, n51789, n51790, n51791, n51792, n51793, n51794, n51795, n51796, n51797, n51798, n51799, n51800, n51801, n51802, n51803, n51804, n51805, n51806, n51807, n51808, n51809, n51810, n51811, n51812, n51813, n51814, n51815, n51816, n51817, n51818, n51819, n51820, n51821, n51822, n51823, n51824, n51825, n51826, n51827, n51828, n51829, n51830, n51831, n51832, n51833, n51834, n51835, n51836, n51837, n51838, n51839, n51840, n51841, n51842, n51843, n51844, n51845, n51846, n51847, n51848, n51849, n51850, n51851, n51852, n51853, n51854, n51855, n51856, n51857, n51858, n51859, n51860, n51861, n51862, n51863, n51864, n51865, n51866, n51867, n51868, n51869, n51870, n51871, n51872, n51873, n51874, n51875, n51876, n51877, n51878, n51879, n51880, n51881, n51882, n51883, n51884, n51885, n51886, n51887, n51888, n51889, n51890, n51891, n51892, n51893, n51894, n51895, n51896, n51897, n51898, n51899, n51900, n51901, n51902, n51903, n51904, n51905, n51906, n51907, n51908, n51909, n51910, n51911, n51912, n51913, n51914, n51915, n51916, n51917, n51918, n51919, n51920, n51921, n51922, n51923, n51924, n51925, n51926, n51927, n51928, n51929, n51930, n51931, n51932, n51933, n51934, n51935, n51936, n51937, n51938, n51939, n51940, n51941, n51942, n51943, n51944, n51945, n51946, n51947, n51948, n51949, n51950, n51951, n51952, n51953, n51954, n51955, n51956, n51957, n51958, n51959, n51960, n51961, n51962, n51963, n51964, n51965, n51966, n51967, n51968, n51969, n51970, n51971, n51972, n51973, n51974, n51975, n51976, n51977, n51978, n51979, n51980, n51981, n51982, n51983, n51984, n51985, n51986, n51987, n51988, n51989, n51990, n51991, n51992, n51993, n51994, n51995, n51996, n51997, n51998, n51999, n52000, n52001, n52002, n52003, n52004, n52005, n52006, n52007, n52008, n52009, n52010, n52011, n52012, n52013, n52014, n52015, n52016, n52017, n52018, n52019, n52020, n52021, n52022, n52023, n52024, n52025, n52026, n52027, n52028, n52029, n52030, n52031, n52032, n52033, n52034, n52035, n52036, n52037, n52038, n52039, n52040, n52041, n52042, n52043, n52044, n52045, n52046, n52047, n52048, n52049, n52050, n52051, n52052, n52053, n52054, n52055, n52056, n52057, n52058, n52059, n52060, n52061, n52062, n52063, n52064, n52065, n52066, n52067, n52068, n52069, n52070, n52071, n52072, n52073, n52074, n52075, n52076, n52077, n52078, n52079, n52080, n52081, n52082, n52083, n52084, n52085, n52086, n52087, n52088, n52089, n52090, n52091, n52092, n52093, n52094, n52095, n52096, n52097, n52098, n52099, n52100, n52101, n52102, n52103, n52104, n52105, n52106, n52107, n52108, n52109, n52110, n52111, n52112, n52113, n52114, n52115, n52116, n52117, n52118, n52119, n52120, n52121, n52122, n52123, n52124, n52125, n52126, n52127, n52128, n52129, n52130, n52131, n52132, n52133, n52134, n52135, n52136, n52137, n52138, n52139, n52140, n52141, n52142, n52143, n52144, n52145, n52146, n52147, n52148, n52149, n52150, n52151, n52152, n52153, n52154, n52155, n52156, n52157, n52158, n52159, n52160, n52161, n52162, n52163, n52164, n52165, n52166, n52167, n52168, n52169, n52170, n52171, n52172, n52173, n52174, n52175, n52176, n52177, n52178, n52179, n52180, n52181, n52182, n52183, n52184, n52185, n52186, n52187, n52188, n52189, n52190, n52191, n52192, n52193, n52194, n52195, n52196, n52197, n52198, n52199, n52200, n52201, n52202, n52203, n52204, n52205, n52206, n52207, n52208, n52209, n52210, n52211, n52212, n52213, n52214, n52215, n52216, n52217, n52218, n52219, n52220, n52221, n52222, n52223, n52224, n52225, n52226, n52227, n52228, n52229, n52230, n52231, n52232, n52233, n52234, n52235, n52236, n52237, n52238, n52239, n52240, n52241, n52242, n52243, n52244, n52245, n52246, n52247, n52248, n52249, n52250, n52251, n52252, n52253, n52254, n52255, n52256, n52257, n52258, n52259, n52260, n52261, n52262, n52263, n52264, n52265, n52266, n52267, n52268, n52269, n52270, n52271, n52272, n52273, n52274, n52275, n52276, n52277, n52278, n52279, n52280, n52281, n52282, n52283, n52284, n52285, n52286, n52287, n52288, n52289, n52290, n52291, n52292, n52293, n52294, n52295, n52296, n52297, n52298, n52299, n52300, n52301, n52302, n52303, n52304, n52305, n52306, n52307, n52308, n52309, n52310, n52311, n52312, n52313, n52314, n52315, n52316, n52317, n52318, n52319, n52320, n52321, n52322, n52323, n52324, n52325, n52326, n52327, n52328, n52329, n52330, n52331, n52332, n52333, n52334, n52335, n52336, n52337, n52338, n52339, n52340, n52341, n52342, n52343, n52344, n52345, n52346, n52347, n52348, n52349, n52350, n52351, n52352, n52353, n52354, n52355, n52356, n52357, n52358, n52359, n52360, n52361, n52362, n52363, n52364, n52365, n52366, n52367, n52368, n52369, n52370, n52371, n52372, n52373, n52374, n52375, n52376, n52377, n52378, n52379, n52380, n52381, n52382, n52383, n52384, n52385, n52386, n52387, n52388, n52389, n52390, n52391, n52392, n52393, n52394, n52395, n52396, n52397, n52398, n52399, n52400, n52401, n52402, n52403, n52404, n52405, n52406, n52407, n52408, n52409, n52410, n52411, n52412, n52413, n52414, n52415, n52416, n52417, n52418, n52419, n52420, n52421, n52422, n52423, n52424, n52425, n52426, n52427, n52428, n52429, n52430, n52431, n52432, n52433, n52434, n52435, n52436, n52437, n52438, n52439, n52440, n52441, n52442, n52443, n52444, n52445, n52446, n52447, n52448, n52449, n52450, n52451, n52452, n52453, n52454, n52455, n52456, n52457, n52458, n52459, n52460, n52461, n52462, n52463, n52464, n52465, n52466, n52467, n52468, n52469, n52470, n52471, n52472, n52473, n52474, n52475, n52476, n52477, n52478, n52479, n52480, n52481, n52482, n52483, n52484, n52485, n52486, n52487, n52488, n52489, n52490, n52491, n52492, n52493, n52494, n52495, n52496, n52497, n52498, n52499, n52500, n52501, n52502, n52503, n52504, n52505, n52506, n52507, n52508, n52509, n52510, n52511, n52512, n52513, n52514, n52515, n52516, n52517, n52518, n52519, n52520, n52521, n52522, n52523, n52524, n52525, n52526, n52527, n52528, n52529, n52530, n52531, n52532, n52533, n52534, n52535, n52536, n52537, n52538, n52539, n52540, n52541, n52542, n52543, n52544, n52545, n52546, n52547, n52548, n52549, n52550, n52551, n52552, n52553, n52554, n52555, n52556, n52557, n52558, n52559, n52560, n52561, n52562, n52563, n52564, n52565, n52566, n52567, n52568, n52569, n52570, n52571, n52572, n52573, n52574, n52575, n52576, n52577, n52578, n52579, n52580, n52581, n52582, n52583, n52584, n52585, n52586, n52587, n52588, n52589, n52590, n52591, n52592, n52593, n52594, n52595, n52596, n52597, n52598, n52599, n52600, n52601, n52602, n52603, n52604, n52605, n52606, n52607, n52608, n52609, n52610, n52611, n52612, n52613, n52614, n52615, n52616, n52617, n52618, n52619, n52620, n52621, n52622, n52623, n52624, n52625, n52626, n52627, n52628, n52629, n52630, n52631, n52632, n52633, n52634, n52635, n52636, n52637, n52638, n52639, n52640, n52641, n52642, n52643, n52644, n52645, n52646, n52647, n52648, n52649, n52650, n52651, n52652, n52653, n52654, n52655, n52656, n52657, n52658, n52659, n52660, n52661, n52662, n52663, n52664, n52665, n52666, n52667, n52668, n52669, n52670, n52671, n52672, n52673, n52674, n52675, n52676, n52677, n52678, n52679, n52680, n52681, n52682, n52683, n52684, n52685, n52686, n52687, n52688, n52689, n52690, n52691, n52692, n52693, n52694, n52695, n52696, n52697, n52698, n52699, n52700, n52701, n52702, n52703, n52704, n52705, n52706, n52707, n52708, n52709, n52710, n52711, n52712, n52713, n52714, n52715, n52716, n52717, n52718, n52719, n52720, n52721, n52722, n52723, n52724, n52725, n52726, n52727, n52728, n52729, n52730, n52731, n52732, n52733, n52734, n52735, n52736, n52737, n52738, n52739, n52740, n52741, n52742, n52743, n52744, n52745, n52746, n52747, n52748, n52749, n52750, n52751, n52752, n52753, n52754, n52755, n52756, n52757, n52758, n52759, n52760, n52761, n52762, n52763, n52764, n52765, n52766, n52767, n52768, n52769, n52770, n52771, n52772, n52773, n52774, n52775, n52776, n52777, n52778, n52779, n52780, n52781, n52782, n52783, n52784, n52785, n52786, n52787, n52788, n52789, n52790, n52791, n52792, n52793, n52794, n52795, n52796, n52797, n52798, n52799, n52800, n52801, n52802, n52803, n52804, n52805, n52806, n52807, n52808, n52809, n52810, n52811, n52812, n52813, n52814, n52815, n52816, n52817, n52818, n52819, n52820, n52821, n52822, n52823, n52824, n52825, n52826, n52827, n52828, n52829, n52830, n52831, n52832, n52833, n52834, n52835, n52836, n52837, n52838, n52839, n52840, n52841, n52842, n52843, n52844, n52845, n52846, n52847, n52848, n52849, n52850, n52851, n52852, n52853, n52854, n52855, n52856, n52857, n52858, n52859, n52860, n52861, n52862, n52863, n52864, n52865, n52866, n52867, n52868, n52869, n52870, n52871, n52872, n52873, n52874, n52875, n52876, n52877, n52878, n52879, n52880, n52881, n52882, n52883, n52884, n52885, n52886, n52887, n52888, n52889, n52890, n52891, n52892, n52893, n52894, n52895, n52896, n52897, n52898, n52899, n52900, n52901, n52902, n52903, n52904, n52905, n52906, n52907, n52908, n52909, n52910, n52911, n52912, n52913, n52914, n52915, n52916, n52917, n52918, n52919, n52920, n52921, n52922, n52923, n52924, n52925, n52926, n52927, n52928, n52929, n52930, n52931, n52932, n52933, n52934, n52935, n52936, n52937, n52938, n52939, n52940, n52941, n52942, n52943, n52944, n52945, n52946, n52947, n52948, n52949, n52950, n52951, n52952, n52953, n52954, n52955, n52956, n52957, n52958, n52959, n52960, n52961, n52962, n52963, n52964, n52965, n52966, n52967, n52968, n52969, n52970, n52971, n52972, n52973, n52974, n52975, n52976, n52977, n52978, n52979, n52980, n52981, n52982, n52983, n52984, n52985, n52986, n52987, n52988, n52989, n52990, n52991, n52992, n52993, n52994, n52995, n52996, n52997, n52998, n52999, n53000, n53001, n53002, n53003, n53004, n53005, n53006, n53007, n53008, n53009, n53010, n53011, n53012, n53013, n53014, n53015, n53016, n53017, n53018, n53019, n53020, n53021, n53022, n53023, n53024, n53025, n53026, n53027, n53028, n53029, n53030, n53031, n53032, n53033, n53034, n53035, n53036, n53037, n53038, n53039, n53040, n53041, n53042, n53043, n53044, n53045, n53046, n53047, n53048, n53049, n53050, n53051, n53052, n53053, n53054, n53055, n53056, n53057, n53058, n53059, n53060, n53061, n53062, n53063, n53064, n53065, n53066, n53067, n53068, n53069, n53070, n53071, n53072, n53073, n53074, n53075, n53076, n53077, n53078, n53079, n53080, n53081, n53082, n53083, n53084, n53085, n53086, n53087, n53088, n53089, n53090, n53091, n53092, n53093, n53094, n53095, n53096, n53097, n53098, n53099, n53100, n53101, n53102, n53103, n53104, n53105, n53106, n53107, n53108, n53109, n53110, n53111, n53112, n53113, n53114, n53115, n53116, n53117, n53118, n53119, n53120, n53121, n53122, n53123, n53124, n53125, n53126, n53127, n53128, n53129, n53130, n53131, n53132, n53133, n53134, n53135, n53136, n53137, n53138, n53139, n53140, n53141, n53142, n53143, n53144, n53145, n53146, n53147, n53148, n53149, n53150, n53151, n53152, n53153, n53154, n53155, n53156, n53157, n53158, n53159, n53160, n53161, n53162, n53163, n53164, n53165, n53166, n53167, n53168, n53169, n53170, n53171, n53172, n53173, n53174, n53175, n53176, n53177, n53178, n53179, n53180, n53181, n53182, n53183, n53184, n53185, n53186, n53187, n53188, n53189, n53190, n53191, n53192, n53193, n53194, n53195, n53196, n53197, n53198, n53199, n53200, n53201, n53202, n53203, n53204, n53205, n53206, n53207, n53208, n53209, n53210, n53211, n53212, n53213, n53214, n53215, n53216, n53217, n53218, n53219, n53220, n53221, n53222, n53223, n53224, n53225, n53226, n53227, n53228, n53229, n53230, n53231, n53232, n53233, n53234, n53235, n53236, n53237, n53238, n53239, n53240, n53241, n53242, n53243, n53244, n53245, n53246, n53247, n53248, n53249, n53250, n53251, n53252, n53253, n53254, n53255, n53256, n53257, n53258, n53259, n53260, n53261, n53262, n53263, n53264, n53265, n53266, n53267, n53268, n53269, n53270, n53271, n53272, n53273, n53274, n53275, n53276, n53277, n53278, n53279, n53280, n53281, n53282, n53283, n53284, n53285, n53286, n53287, n53288, n53289, n53290, n53291, n53292, n53293, n53294, n53295, n53296, n53297, n53298, n53299, n53300, n53301, n53302, n53303, n53304, n53305, n53306, n53307, n53308, n53309, n53310, n53311, n53312, n53313, n53314, n53315, n53316, n53317, n53318, n53319, n53320, n53321, n53322, n53323, n53324, n53325, n53326, n53327, n53328, n53329, n53330, n53331, n53332, n53333, n53334, n53335, n53336, n53337, n53338, n53339, n53340, n53341, n53342, n53343, n53344, n53345, n53346, n53347, n53348, n53349, n53350, n53351, n53352, n53353, n53354, n53355, n53356, n53357, n53358, n53359, n53360, n53361, n53362, n53363, n53364, n53365, n53366, n53367, n53368, n53369, n53370, n53371, n53372, n53373, n53374, n53375, n53376, n53377, n53378, n53379, n53380, n53381, n53382, n53383, n53384, n53385, n53386, n53387, n53388, n53389, n53390, n53391, n53392, n53393, n53394, n53395, n53396, n53397, n53398, n53399, n53400, n53401, n53402, n53403, n53404, n53405, n53406, n53407, n53408, n53409, n53410, n53411, n53412, n53413, n53414, n53415, n53416, n53417, n53418, n53419, n53420, n53421, n53422, n53423, n53424, n53425, n53426, n53427, n53428, n53429, n53430, n53431, n53432, n53433, n53434, n53435, n53436, n53437, n53438, n53439, n53440, n53441, n53442, n53443, n53444, n53445, n53446, n53447, n53448, n53449, n53450, n53451, n53452, n53453, n53454, n53455, n53456, n53457, n53458, n53459, n53460, n53461, n53462, n53463, n53464, n53465, n53466, n53467, n53468, n53469, n53470, n53471, n53472, n53473, n53474, n53475, n53476, n53477, n53478, n53479, n53480, n53481, n53482, n53483, n53484, n53485, n53486, n53487, n53488, n53489, n53490, n53491, n53492, n53493, n53494, n53495, n53496, n53497, n53498, n53499, n53500, n53501, n53502, n53503, n53504, n53505, n53506, n53507, n53508, n53509, n53510, n53511, n53512, n53513, n53514, n53515, n53516, n53517, n53518, n53519, n53520, n53521, n53522, n53523, n53524, n53525, n53526, n53527, n53528, n53529, n53530, n53531, n53532, n53533, n53534, n53535, n53536, n53537, n53538, n53539, n53540, n53541, n53542, n53543, n53544, n53545, n53546, n53547, n53548, n53549, n53550, n53551, n53552, n53553, n53554, n53555, n53556, n53557, n53558, n53559, n53560, n53561, n53562, n53563, n53564, n53565, n53566, n53567, n53568, n53569, n53570, n53571, n53572, n53573, n53574, n53575, n53576, n53577, n53578, n53579, n53580, n53581, n53582, n53583, n53584, n53585, n53586, n53587, n53588, n53589, n53590, n53591, n53592, n53593, n53594, n53595, n53596, n53597, n53598, n53599, n53600, n53601, n53602, n53603, n53604, n53605, n53606, n53607, n53608, n53609, n53610, n53611, n53612, n53613, n53614, n53615, n53616, n53617, n53618, n53619, n53620, n53621, n53622, n53623, n53624, n53625, n53626, n53627, n53628, n53629, n53630, n53631, n53632, n53633, n53634, n53635, n53636, n53637, n53638, n53639, n53640, n53641, n53642, n53643, n53644, n53645, n53646, n53647, n53648, n53649, n53650, n53651, n53652, n53653, n53654, n53655, n53656, n53657, n53658, n53659, n53660, n53661, n53662, n53663, n53664, n53665, n53666, n53667, n53668, n53669, n53670, n53671, n53672, n53673, n53674, n53675, n53676, n53677, n53678, n53679, n53680, n53681, n53682, n53683, n53684, n53685, n53686, n53687, n53688, n53689, n53690, n53691, n53692, n53693, n53694, n53695, n53696, n53697, n53698, n53699, n53700, n53701, n53702, n53703, n53704, n53705, n53706, n53707, n53708, n53709, n53710, n53711, n53712, n53713, n53714, n53715, n53716, n53717, n53718, n53719, n53720, n53721, n53722, n53723, n53724, n53725, n53726, n53727, n53728, n53729, n53730, n53731, n53732, n53733, n53734, n53735, n53736, n53737, n53738, n53739, n53740, n53741, n53742, n53743, n53744, n53745, n53746, n53747, n53748, n53749, n53750, n53751, n53752, n53753, n53754, n53755, n53756, n53757, n53758, n53759, n53760, n53761, n53762, n53763, n53764, n53765, n53766, n53767, n53768, n53769, n53770, n53771, n53772, n53773, n53774, n53775, n53776, n53777, n53778, n53779, n53780, n53781, n53782, n53783, n53784, n53785, n53786, n53787, n53788, n53789, n53790, n53791, n53792, n53793, n53794, n53795, n53796, n53797, n53798, n53799, n53800, n53801, n53802, n53803, n53804, n53805, n53806, n53807, n53808, n53809, n53810, n53811, n53812, n53813, n53814, n53815, n53816, n53817, n53818, n53819, n53820, n53821, n53822, n53823, n53824, n53825, n53826, n53827, n53828, n53829, n53830, n53831, n53832, n53833, n53834, n53835, n53836, n53837, n53838, n53839, n53840, n53841, n53842, n53843, n53844, n53845, n53846, n53847, n53848, n53849, n53850, n53851, n53852, n53853, n53854, n53855, n53856, n53857, n53858, n53859, n53860, n53861, n53862, n53863, n53864, n53865, n53866, n53867, n53868, n53869, n53870, n53871, n53872, n53873, n53874, n53875, n53876, n53877, n53878, n53879, n53880, n53881, n53882, n53883, n53884, n53885, n53886, n53887, n53888, n53889, n53890, n53891, n53892, n53893, n53894, n53895, n53896, n53897, n53898, n53899, n53900, n53901, n53902, n53903, n53904, n53905, n53906, n53907, n53908, n53909, n53910, n53911, n53912, n53913, n53914, n53915, n53916, n53917, n53918, n53919, n53920, n53921, n53922, n53923, n53924, n53925, n53926, n53927, n53928, n53929, n53930, n53931, n53932, n53933, n53934, n53935, n53936, n53937, n53938, n53939, n53940, n53941, n53942, n53943, n53944, n53945, n53946, n53947, n53948, n53949, n53950, n53951, n53952, n53953, n53954, n53955, n53956, n53957, n53958, n53959, n53960, n53961, n53962, n53963, n53964, n53965, n53966, n53967, n53968, n53969, n53970, n53971, n53972, n53973, n53974, n53975, n53976, n53977, n53978, n53979, n53980, n53981, n53982, n53983, n53984, n53985, n53986, n53987, n53988, n53989, n53990, n53991, n53992, n53993, n53994, n53995, n53996, n53997, n53998, n53999, n54000, n54001, n54002, n54003, n54004, n54005, n54006, n54007, n54008, n54009, n54010, n54011, n54012, n54013, n54014, n54015, n54016, n54017, n54018, n54019, n54020, n54021, n54022, n54023, n54024, n54025, n54026, n54027, n54028, n54029, n54030, n54031, n54032, n54033, n54034, n54035, n54036, n54037, n54038, n54039, n54040, n54041, n54042, n54043, n54044, n54045, n54046, n54047, n54048, n54049, n54050, n54051, n54052, n54053, n54054, n54055, n54056, n54057, n54058, n54059, n54060, n54061, n54062, n54063, n54064, n54065, n54066, n54067, n54068, n54069, n54070, n54071, n54072, n54073, n54074, n54075, n54076, n54077, n54078, n54079, n54080, n54081, n54082, n54083, n54084, n54085, n54086, n54087, n54088, n54089, n54090, n54091, n54092, n54093, n54094, n54095, n54096, n54097, n54098, n54099, n54100, n54101, n54102, n54103, n54104, n54105, n54106, n54107, n54108, n54109, n54110, n54111, n54112, n54113, n54114, n54115, n54116, n54117, n54118, n54119, n54120, n54121, n54122, n54123, n54124, n54125, n54126, n54127, n54128, n54129, n54130, n54131, n54132, n54133, n54134, n54135, n54136, n54137, n54138, n54139, n54140, n54141, n54142, n54143, n54144, n54145, n54146, n54147, n54148, n54149, n54150, n54151, n54152, n54153, n54154, n54155, n54156, n54157, n54158, n54159, n54160, n54161, n54162, n54163, n54164, n54165, n54166, n54167, n54168, n54169, n54170, n54171, n54172, n54173, n54174, n54175, n54176, n54177, n54178, n54179, n54180, n54181, n54182, n54183, n54184, n54185, n54186, n54187, n54188, n54189, n54190, n54191, n54192, n54193, n54194, n54195, n54196, n54197, n54198, n54199, n54200, n54201, n54202, n54203, n54204, n54205, n54206, n54207, n54208, n54209, n54210, n54211, n54212, n54213, n54214, n54215, n54216, n54217, n54218, n54219, n54220, n54221, n54222, n54223, n54224, n54225, n54226, n54227, n54228, n54229, n54230, n54231, n54232, n54233, n54234, n54235, n54236, n54237, n54238, n54239, n54240, n54241, n54242, n54243, n54244, n54245, n54246, n54247, n54248, n54249, n54250, n54251, n54252, n54253, n54254, n54255, n54256, n54257, n54258, n54259, n54260, n54261, n54262, n54263, n54264, n54265, n54266, n54267, n54268, n54269, n54270, n54271, n54272, n54273, n54274, n54275, n54276, n54277, n54278, n54279, n54280, n54281, n54282, n54283, n54284, n54285, n54286, n54287, n54288, n54289, n54290, n54291, n54292, n54293, n54294, n54295, n54296, n54297, n54298, n54299, n54300, n54301, n54302, n54303, n54304, n54305, n54306, n54307, n54308, n54309, n54310, n54311, n54312, n54313, n54314, n54315, n54316, n54317, n54318, n54319, n54320, n54321, n54322, n54323, n54324, n54325, n54326, n54327, n54328, n54329, n54330, n54331, n54332, n54333, n54334, n54335, n54336, n54337, n54338, n54339, n54340, n54341, n54342, n54343, n54344, n54345, n54346, n54347, n54348, n54349, n54350, n54351, n54352, n54353, n54354, n54355, n54356, n54357, n54358, n54359, n54360, n54361, n54362, n54363, n54364, n54365, n54366, n54367, n54368, n54369, n54370, n54371, n54372, n54373, n54374, n54375, n54376, n54377, n54378, n54379, n54380, n54381, n54382, n54383, n54384, n54385, n54386, n54387, n54388, n54389, n54390, n54391, n54392, n54393, n54394, n54395, n54396, n54397, n54398, n54399, n54400, n54401, n54402, n54403, n54404, n54405, n54406, n54407, n54408, n54409, n54410, n54411, n54412, n54413, n54414, n54415, n54416, n54417, n54418, n54419, n54420, n54421, n54422, n54423, n54424, n54425, n54426, n54427, n54428, n54429, n54430, n54431, n54432, n54433, n54434, n54435, n54436, n54437, n54438, n54439, n54440, n54441, n54442, n54443, n54444, n54445, n54446, n54447, n54448, n54449, n54450, n54451, n54452, n54453, n54454, n54455, n54456, n54457, n54458, n54459, n54460, n54461, n54462, n54463, n54464, n54465, n54466, n54467, n54468, n54469, n54470, n54471, n54472, n54473, n54474, n54475, n54476, n54477, n54478, n54479, n54480, n54481, n54482, n54483, n54484, n54485, n54486, n54487, n54488, n54489, n54490, n54491, n54492, n54493, n54494, n54495, n54496, n54497, n54498, n54499, n54500, n54501, n54502, n54503, n54504, n54505, n54506, n54507, n54508, n54509, n54510, n54511, n54512, n54513, n54514, n54515, n54516, n54517, n54518, n54519, n54520, n54521, n54522, n54523, n54524, n54525, n54526, n54527, n54528, n54529, n54530, n54531, n54532, n54533, n54534, n54535, n54536, n54537, n54538, n54539, n54540, n54541, n54542, n54543, n54544, n54545, n54546, n54547, n54548, n54549, n54550, n54551, n54552, n54553, n54554, n54555, n54556, n54557, n54558, n54559, n54560, n54561, n54562, n54563, n54564, n54565, n54566, n54567, n54568, n54569, n54570, n54571, n54572, n54573, n54574, n54575, n54576, n54577, n54578, n54579, n54580, n54581, n54582, n54583, n54584, n54585, n54586, n54587, n54588, n54589, n54590, n54591, n54592, n54593, n54594, n54595, n54596, n54597, n54598, n54599, n54600, n54601, n54602, n54603, n54604, n54605, n54606, n54607, n54608, n54609, n54610, n54611, n54612, n54613, n54614, n54615, n54616, n54617, n54618, n54619, n54620, n54621, n54622, n54623, n54624, n54625, n54626, n54627, n54628, n54629, n54630, n54631, n54632, n54633, n54634, n54635, n54636, n54637, n54638, n54639, n54640, n54641, n54642, n54643, n54644, n54645, n54646, n54647, n54648, n54649, n54650, n54651, n54652, n54653, n54654, n54655, n54656, n54657, n54658, n54659, n54660, n54661, n54662, n54663, n54664, n54665, n54666, n54667, n54668, n54669, n54670, n54671, n54672, n54673, n54674, n54675, n54676, n54677, n54678, n54679, n54680, n54681, n54682, n54683, n54684, n54685, n54686, n54687, n54688, n54689, n54690, n54691, n54692, n54693, n54694, n54695, n54696, n54697, n54698, n54699, n54700, n54701, n54702, n54703, n54704, n54705, n54706, n54707, n54708, n54709, n54710, n54711, n54712, n54713, n54714, n54715, n54716, n54717, n54718, n54719, n54720, n54721, n54722, n54723, n54724, n54725, n54726, n54727, n54728, n54729, n54730, n54731, n54732, n54733, n54734, n54735, n54736, n54737, n54738, n54739, n54740, n54741, n54742, n54743, n54744, n54745, n54746, n54747, n54748, n54749, n54750, n54751, n54752, n54753, n54754, n54755, n54756, n54757, n54758, n54759, n54760, n54761, n54762, n54763, n54764, n54765, n54766, n54767, n54768, n54769, n54770, n54771, n54772, n54773, n54774, n54775, n54776, n54777, n54778, n54779, n54780, n54781, n54782, n54783, n54784, n54785, n54786, n54787, n54788, n54789, n54790, n54791, n54792, n54793, n54794, n54795, n54796, n54797, n54798, n54799, n54800, n54801, n54802, n54803, n54804, n54805, n54806, n54807, n54808, n54809, n54810, n54811, n54812, n54813, n54814, n54815, n54816, n54817, n54818, n54819, n54820, n54821, n54822, n54823, n54824, n54825, n54826, n54827, n54828, n54829, n54830, n54831, n54832, n54833, n54834, n54835, n54836, n54837, n54838, n54839, n54840, n54841, n54842, n54843, n54844, n54845, n54846, n54847, n54848, n54849, n54850, n54851, n54852, n54853, n54854, n54855, n54856, n54857, n54858, n54859, n54860, n54861, n54862, n54863, n54864, n54865, n54866, n54867, n54868, n54869, n54870, n54871, n54872, n54873, n54874, n54875, n54876, n54877, n54878, n54879, n54880, n54881, n54882, n54883, n54884, n54885, n54886, n54887, n54888, n54889, n54890, n54891, n54892, n54893, n54894, n54895, n54896, n54897, n54898, n54899, n54900, n54901, n54902, n54903, n54904, n54905, n54906, n54907, n54908, n54909, n54910, n54911, n54912, n54913, n54914, n54915, n54916, n54917, n54918, n54919, n54920, n54921, n54922, n54923, n54924, n54925, n54926, n54927, n54928, n54929, n54930, n54931, n54932, n54933, n54934, n54935, n54936, n54937, n54938, n54939, n54940, n54941, n54942, n54943, n54944, n54945, n54946, n54947, n54948, n54949, n54950, n54951, n54952, n54953, n54954, n54955, n54956, n54957, n54958, n54959, n54960, n54961, n54962, n54963, n54964, n54965, n54966, n54967, n54968, n54969, n54970, n54971, n54972, n54973, n54974, n54975, n54976, n54977, n54978, n54979, n54980, n54981, n54982, n54983, n54984, n54985, n54986, n54987, n54988, n54989, n54990, n54991, n54992, n54993, n54994, n54995, n54996, n54997, n54998, n54999, n55000, n55001, n55002, n55003, n55004, n55005, n55006, n55007, n55008, n55009, n55010, n55011, n55012, n55013, n55014, n55015, n55016, n55017, n55018, n55019, n55020, n55021, n55022, n55023, n55024, n55025, n55026, n55027, n55028, n55029, n55030, n55031, n55032, n55033, n55034, n55035, n55036, n55037, n55038, n55039, n55040, n55041, n55042, n55043, n55044, n55045, n55046, n55047, n55048, n55049, n55050, n55051, n55052, n55053, n55054, n55055, n55056, n55057, n55058, n55059, n55060, n55061, n55062, n55063, n55064, n55065, n55066, n55067, n55068, n55069, n55070, n55071, n55072, n55073, n55074, n55075, n55076, n55077, n55078, n55079, n55080, n55081, n55082, n55083, n55084, n55085, n55086, n55087, n55088, n55089, n55090, n55091, n55092, n55093, n55094, n55095, n55096, n55097, n55098, n55099, n55100, n55101, n55102, n55103, n55104, n55105, n55106, n55107, n55108, n55109, n55110, n55111, n55112, n55113, n55114, n55115, n55116, n55117, n55118, n55119, n55120, n55121, n55122, n55123, n55124, n55125, n55126, n55127, n55128, n55129, n55130, n55131, n55132, n55133, n55134, n55135, n55136, n55137, n55138, n55139, n55140, n55141, n55142, n55143, n55144, n55145, n55146, n55147, n55148, n55149, n55150, n55151, n55152, n55153, n55154, n55155, n55156, n55157, n55158, n55159, n55160, n55161, n55162, n55163, n55164, n55165, n55166, n55167, n55168, n55169, n55170, n55171, n55172, n55173, n55174, n55175, n55176, n55177, n55178, n55179, n55180, n55181, n55182, n55183, n55184, n55185, n55186, n55187, n55188, n55189, n55190, n55191, n55192, n55193, n55194, n55195, n55196, n55197, n55198, n55199, n55200, n55201, n55202, n55203, n55204, n55205, n55206, n55207, n55208, n55209, n55210, n55211, n55212, n55213, n55214, n55215, n55216, n55217, n55218, n55219, n55220, n55221, n55222, n55223, n55224, n55225, n55226, n55227, n55228, n55229, n55230, n55231, n55232, n55233, n55234, n55235, n55236, n55237, n55238, n55239, n55240, n55241, n55242, n55243, n55244, n55245, n55246, n55247, n55248, n55249, n55250, n55251, n55252, n55253, n55254, n55255, n55256, n55257, n55258, n55259, n55260, n55261, n55262, n55263, n55264, n55265, n55266, n55267, n55268, n55269, n55270, n55271, n55272, n55273, n55274, n55275, n55276, n55277, n55278, n55279, n55280, n55281, n55282, n55283, n55284, n55285, n55286, n55287, n55288, n55289, n55290, n55291, n55292, n55293, n55294, n55295, n55296, n55297, n55298, n55299, n55300, n55301, n55302, n55303, n55304, n55305, n55306, n55307, n55308, n55309, n55310, n55311, n55312, n55313, n55314, n55315, n55316, n55317, n55318, n55319, n55320, n55321, n55322, n55323, n55324, n55325, n55326, n55327, n55328, n55329, n55330, n55331, n55332, n55333, n55334, n55335, n55336, n55337, n55338, n55339, n55340, n55341, n55342, n55343, n55344, n55345, n55346, n55347, n55348, n55349, n55350, n55351, n55352, n55353, n55354, n55355, n55356, n55357, n55358, n55359, n55360, n55361, n55362, n55363, n55364, n55365, n55366, n55367, n55368, n55369, n55370, n55371, n55372, n55373, n55374, n55375, n55376, n55377, n55378, n55379, n55380, n55381, n55382, n55383, n55384, n55385, n55386, n55387, n55388, n55389, n55390, n55391, n55392, n55393, n55394, n55395, n55396, n55397, n55398, n55399, n55400, n55401, n55402, n55403, n55404, n55405, n55406, n55407, n55408, n55409, n55410, n55411, n55412, n55413, n55414, n55415, n55416, n55417, n55418, n55419, n55420, n55421, n55422, n55423, n55424, n55425, n55426, n55427, n55428, n55429, n55430, n55431, n55432, n55433, n55434, n55435, n55436, n55437, n55438, n55439, n55440, n55441, n55442, n55443, n55444, n55445, n55446, n55447, n55448, n55449, n55450, n55451, n55452, n55453, n55454, n55455, n55456, n55457, n55458, n55459, n55460, n55461, n55462, n55463, n55464, n55465, n55466, n55467, n55468, n55469, n55470, n55471, n55472, n55473, n55474, n55475, n55476, n55477, n55478, n55479, n55480, n55481, n55482, n55483, n55484, n55485, n55486, n55487, n55488, n55489, n55490, n55491, n55492, n55493, n55494, n55495, n55496, n55497, n55498, n55499, n55500, n55501, n55502, n55503, n55504, n55505, n55506, n55507, n55508, n55509, n55510, n55511, n55512, n55513, n55514, n55515, n55516, n55517, n55518, n55519, n55520, n55521, n55522, n55523, n55524, n55525, n55526, n55527, n55528, n55529, n55530, n55531, n55532, n55533, n55534, n55535, n55536, n55537, n55538, n55539, n55540, n55541, n55542, n55543, n55544, n55545, n55546, n55547, n55548, n55549, n55550, n55551, n55552, n55553, n55554, n55555, n55556, n55557, n55558, n55559, n55560, n55561, n55562, n55563, n55564, n55565, n55566, n55567, n55568, n55569, n55570, n55571, n55572, n55573, n55574, n55575, n55576, n55577, n55578, n55579, n55580, n55581, n55582, n55583, n55584, n55585, n55586, n55587, n55588, n55589, n55590, n55591, n55592, n55593, n55594, n55595, n55596, n55597, n55598, n55599, n55600, n55601, n55602, n55603, n55604, n55605, n55606, n55607, n55608, n55609, n55610, n55611, n55612, n55613, n55614, n55615, n55616, n55617, n55618, n55619, n55620, n55621, n55622, n55623, n55624, n55625, n55626, n55627, n55628, n55629, n55630, n55631, n55632, n55633, n55634, n55635, n55636, n55637, n55638, n55639, n55640, n55641, n55642, n55643, n55644, n55645, n55646, n55647, n55648, n55649, n55650, n55651, n55652, n55653, n55654, n55655, n55656, n55657, n55658, n55659, n55660, n55661, n55662, n55663, n55664, n55665, n55666, n55667, n55668, n55669, n55670, n55671, n55672, n55673, n55674, n55675, n55676, n55677, n55678, n55679, n55680, n55681, n55682, n55683, n55684, n55685, n55686, n55687, n55688, n55689, n55690, n55691, n55692, n55693, n55694, n55695, n55696, n55697, n55698, n55699, n55700, n55701, n55702, n55703, n55704, n55705, n55706, n55707, n55708, n55709, n55710, n55711, n55712, n55713, n55714, n55715, n55716, n55717, n55718, n55719, n55720, n55721, n55722, n55723, n55724, n55725, n55726, n55727, n55728, n55729, n55730, n55731, n55732, n55733, n55734, n55735, n55736, n55737, n55738, n55739, n55740, n55741, n55742, n55743, n55744, n55745, n55746, n55747, n55748, n55749, n55750, n55751, n55752, n55753, n55754, n55755, n55756, n55757, n55758, n55759, n55760, n55761, n55762, n55763, n55764, n55765, n55766, n55767, n55768, n55769, n55770, n55771, n55772, n55773, n55774, n55775, n55776, n55777, n55778, n55779, n55780, n55781, n55782, n55783, n55784, n55785, n55786, n55787, n55788, n55789, n55790, n55791, n55792, n55793, n55794, n55795, n55796, n55797, n55798, n55799, n55800, n55801, n55802, n55803, n55804, n55805, n55806, n55807, n55808, n55809, n55810, n55811, n55812, n55813, n55814, n55815, n55816, n55817, n55818, n55819, n55820, n55821, n55822, n55823, n55824, n55825, n55826, n55827, n55828, n55829, n55830, n55831, n55832, n55833, n55834, n55835, n55836, n55837, n55838, n55839, n55840, n55841, n55842, n55843, n55844, n55845, n55846, n55847, n55848, n55849, n55850, n55851, n55852, n55853, n55854, n55855, n55856, n55857, n55858, n55859, n55860, n55861, n55862, n55863, n55864, n55865, n55866, n55867, n55868, n55869, n55870, n55871, n55872, n55873, n55874, n55875, n55876, n55877, n55878, n55879, n55880, n55881, n55882, n55883, n55884, n55885, n55886, n55887, n55888, n55889, n55890, n55891, n55892, n55893, n55894, n55895, n55896, n55897, n55898, n55899, n55900, n55901, n55902, n55903, n55904, n55905, n55906, n55907, n55908, n55909, n55910, n55911, n55912, n55913, n55914, n55915, n55916, n55917, n55918, n55919, n55920, n55921, n55922, n55923, n55924, n55925, n55926, n55927, n55928, n55929, n55930, n55931, n55932, n55933, n55934, n55935, n55936, n55937, n55938, n55939, n55940, n55941, n55942, n55943, n55944, n55945, n55946, n55947, n55948, n55949, n55950, n55951, n55952, n55953, n55954, n55955, n55956, n55957, n55958, n55959, n55960, n55961, n55962, n55963, n55964, n55965, n55966, n55967, n55968, n55969, n55970, n55971, n55972, n55973, n55974, n55975, n55976, n55977, n55978, n55979, n55980, n55981, n55982, n55983, n55984, n55985, n55986, n55987, n55988, n55989, n55990, n55991, n55992, n55993, n55994, n55995, n55996, n55997, n55998, n55999, n56000, n56001, n56002, n56003, n56004, n56005, n56006, n56007, n56008, n56009, n56010, n56011, n56012, n56013, n56014, n56015, n56016, n56017, n56018, n56019, n56020, n56021, n56022, n56023, n56024, n56025, n56026, n56027, n56028, n56029, n56030, n56031, n56032, n56033, n56034, n56035, n56036, n56037, n56038, n56039, n56040, n56041, n56042, n56043, n56044, n56045, n56046, n56047, n56048, n56049, n56050, n56051, n56052, n56053, n56054, n56055, n56056, n56057, n56058, n56059, n56060, n56061, n56062, n56063, n56064, n56065, n56066, n56067, n56068, n56069, n56070, n56071, n56072, n56073, n56074, n56075, n56076, n56077, n56078, n56079, n56080, n56081, n56082, n56083, n56084, n56085, n56086, n56087, n56088, n56089, n56090, n56091, n56092, n56093, n56094, n56095, n56096, n56097, n56098, n56099, n56100, n56101, n56102, n56103, n56104, n56105, n56106, n56107, n56108, n56109, n56110, n56111, n56112, n56113, n56114, n56115, n56116, n56117, n56118, n56119, n56120, n56121, n56122, n56123, n56124, n56125, n56126, n56127, n56128, n56129, n56130, n56131, n56132, n56133, n56134, n56135, n56136, n56137, n56138, n56139, n56140, n56141, n56142, n56143, n56144, n56145, n56146, n56147, n56148, n56149, n56150, n56151, n56152, n56153, n56154, n56155, n56156, n56157, n56158, n56159, n56160, n56161, n56162, n56163, n56164, n56165, n56166, n56167, n56168, n56169, n56170, n56171, n56172, n56173, n56174, n56175, n56176, n56177, n56178, n56179, n56180, n56181, n56182, n56183, n56184, n56185, n56186, n56187, n56188, n56189, n56190, n56191, n56192, n56193, n56194, n56195, n56196, n56197, n56198, n56199, n56200, n56201, n56202, n56203, n56204, n56205, n56206, n56207, n56208, n56209, n56210, n56211, n56212, n56213, n56214, n56215, n56216, n56217, n56218, n56219, n56220, n56221, n56222, n56223, n56224, n56225, n56226, n56227, n56228, n56229, n56230, n56231, n56232, n56233, n56234, n56235, n56236, n56237, n56238, n56239, n56240, n56241, n56242, n56243, n56244, n56245, n56246, n56247, n56248, n56249, n56250, n56251, n56252, n56253, n56254, n56255, n56256, n56257, n56258, n56259, n56260, n56261, n56262, n56263, n56264, n56265, n56266, n56267, n56268, n56269, n56270, n56271, n56272, n56273, n56274, n56275, n56276, n56277, n56278, n56279, n56280, n56281, n56282, n56283, n56284, n56285, n56286, n56287, n56288, n56289, n56290, n56291, n56292, n56293, n56294, n56295, n56296, n56297, n56298, n56299, n56300, n56301, n56302, n56303, n56304, n56305, n56306, n56307, n56308, n56309, n56310, n56311, n56312, n56313, n56314, n56315, n56316, n56317, n56318, n56319, n56320, n56321, n56322, n56323, n56324, n56325, n56326, n56327, n56328, n56329, n56330, n56331, n56332, n56333, n56334, n56335, n56336, n56337, n56338, n56339, n56340, n56341, n56342, n56343, n56344, n56345, n56346, n56347, n56348, n56349, n56350, n56351, n56352, n56353, n56354, n56355, n56356, n56357, n56358, n56359, n56360, n56361, n56362, n56363, n56364, n56365, n56366, n56367, n56368, n56369, n56370, n56371, n56372, n56373, n56374, n56375, n56376, n56377, n56378, n56379, n56380, n56381, n56382, n56383, n56384, n56385, n56386, n56387, n56388, n56389, n56390, n56391, n56392, n56393, n56394, n56395, n56396, n56397, n56398, n56399, n56400, n56401, n56402, n56403, n56404, n56405, n56406, n56407, n56408, n56409, n56410, n56411, n56412, n56413, n56414, n56415, n56416, n56417, n56418, n56419, n56420, n56421, n56422, n56423, n56424, n56425, n56426, n56427, n56428, n56429, n56430, n56431, n56432, n56433, n56434, n56435, n56436, n56437, n56438, n56439, n56440, n56441, n56442, n56443, n56444, n56445, n56446, n56447, n56448, n56449, n56450, n56451, n56452, n56453, n56454, n56455, n56456, n56457, n56458, n56459, n56460, n56461, n56462, n56463, n56464, n56465, n56466, n56467, n56468, n56469, n56470, n56471, n56472, n56473, n56474, n56475, n56476, n56477, n56478, n56479, n56480, n56481, n56482, n56483, n56484, n56485, n56486, n56487, n56488, n56489, n56490, n56491, n56492, n56493, n56494, n56495, n56496, n56497, n56498, n56499, n56500, n56501, n56502, n56503, n56504, n56505, n56506, n56507, n56508, n56509, n56510, n56511, n56512, n56513, n56514, n56515, n56516, n56517, n56518, n56519, n56520, n56521, n56522, n56523, n56524, n56525, n56526, n56527, n56528, n56529, n56530, n56531, n56532, n56533, n56534, n56535, n56536, n56537, n56538, n56539, n56540, n56541, n56542, n56543, n56544, n56545, n56546, n56547, n56548, n56549, n56550, n56551, n56552, n56553, n56554, n56555, n56556, n56557, n56558, n56559, n56560, n56561, n56562, n56563, n56564, n56565, n56566, n56567, n56568, n56569, n56570, n56571, n56572, n56573, n56574, n56575, n56576, n56577, n56578, n56579, n56580, n56581, n56582, n56583, n56584, n56585, n56586, n56587, n56588, n56589, n56590, n56591, n56592, n56593, n56594, n56595, n56596, n56597, n56598, n56599, n56600, n56601, n56602, n56603, n56604, n56605, n56606, n56607, n56608, n56609, n56610, n56611, n56612, n56613, n56614, n56615, n56616, n56617, n56618, n56619, n56620, n56621, n56622, n56623, n56624, n56625, n56626, n56627, n56628, n56629, n56630, n56631, n56632, n56633, n56634, n56635, n56636, n56637, n56638, n56639, n56640, n56641, n56642, n56643, n56644, n56645, n56646, n56647, n56648, n56649, n56650, n56651, n56652, n56653, n56654, n56655, n56656, n56657, n56658, n56659, n56660, n56661, n56662, n56663, n56664, n56665, n56666, n56667, n56668, n56669, n56670, n56671, n56672, n56673, n56674, n56675, n56676, n56677, n56678, n56679, n56680, n56681, n56682, n56683, n56684, n56685, n56686, n56687, n56688, n56689, n56690, n56691, n56692, n56693, n56694, n56695, n56696, n56697, n56698, n56699, n56700, n56701, n56702, n56703, n56704, n56705, n56706, n56707, n56708, n56709, n56710, n56711, n56712, n56713, n56714, n56715, n56716, n56717, n56718, n56719, n56720, n56721, n56722, n56723, n56724, n56725, n56726, n56727, n56728, n56729, n56730, n56731, n56732, n56733, n56734, n56735, n56736, n56737, n56738, n56739, n56740, n56741, n56742, n56743, n56744, n56745, n56746, n56747, n56748, n56749, n56750, n56751, n56752, n56753, n56754, n56755, n56756, n56757, n56758, n56759, n56760, n56761, n56762, n56763, n56764, n56765, n56766, n56767, n56768, n56769, n56770, n56771, n56772, n56773, n56774, n56775, n56776, n56777, n56778, n56779, n56780, n56781, n56782, n56783, n56784, n56785, n56786, n56787, n56788, n56789, n56790, n56791, n56792, n56793, n56794, n56795, n56796, n56797, n56798, n56799, n56800, n56801, n56802, n56803, n56804, n56805, n56806, n56807, n56808, n56809, n56810, n56811, n56812, n56813, n56814, n56815, n56816, n56817, n56818, n56819, n56820, n56821, n56822, n56823, n56824, n56825, n56826, n56827, n56828, n56829, n56830, n56831, n56832, n56833, n56834, n56835, n56836, n56837, n56838, n56839, n56840, n56841, n56842, n56843, n56844, n56845, n56846, n56847, n56848, n56849, n56850, n56851, n56852, n56853, n56854, n56855, n56856, n56857, n56858, n56859, n56860, n56861, n56862, n56863, n56864, n56865, n56866, n56867, n56868, n56869, n56870, n56871, n56872, n56873, n56874, n56875, n56876, n56877, n56878, n56879, n56880, n56881, n56882, n56883, n56884, n56885, n56886, n56887, n56888, n56889, n56890, n56891, n56892, n56893, n56894, n56895, n56896, n56897, n56898, n56899, n56900, n56901, n56902, n56903, n56904, n56905, n56906, n56907, n56908, n56909, n56910, n56911, n56912, n56913, n56914, n56915, n56916, n56917, n56918, n56919, n56920, n56921, n56922, n56923, n56924, n56925, n56926, n56927, n56928, n56929, n56930, n56931, n56932, n56933, n56934, n56935, n56936, n56937, n56938, n56939, n56940, n56941, n56942, n56943, n56944, n56945, n56946, n56947, n56948, n56949, n56950, n56951, n56952, n56953, n56954, n56955, n56956, n56957, n56958, n56959, n56960, n56961, n56962, n56963, n56964, n56965, n56966, n56967, n56968, n56969, n56970, n56971, n56972, n56973, n56974, n56975, n56976, n56977, n56978, n56979, n56980, n56981, n56982, n56983, n56984, n56985, n56986, n56987, n56988, n56989, n56990, n56991, n56992, n56993, n56994, n56995, n56996, n56997, n56998, n56999, n57000, n57001, n57002, n57003, n57004, n57005, n57006, n57007, n57008, n57009, n57010, n57011, n57012, n57013, n57014, n57015, n57016, n57017, n57018, n57019, n57020, n57021, n57022, n57023, n57024, n57025, n57026, n57027, n57028, n57029, n57030, n57031, n57032, n57033, n57034, n57035, n57036, n57037, n57038, n57039, n57040, n57041, n57042, n57043, n57044, n57045, n57046, n57047, n57048, n57049, n57050, n57051, n57052, n57053, n57054, n57055, n57056, n57057, n57058, n57059, n57060, n57061, n57062, n57063, n57064, n57065, n57066, n57067, n57068, n57069, n57070, n57071, n57072, n57073, n57074, n57075, n57076, n57077, n57078, n57079, n57080, n57081, n57082, n57083, n57084, n57085, n57086, n57087, n57088, n57089, n57090, n57091, n57092, n57093, n57094, n57095, n57096, n57097, n57098, n57099, n57100, n57101, n57102, n57103, n57104, n57105, n57106, n57107, n57108, n57109, n57110, n57111, n57112, n57113, n57114, n57115, n57116, n57117, n57118, n57119, n57120, n57121, n57122, n57123, n57124, n57125, n57126, n57127, n57128, n57129, n57130, n57131, n57132, n57133, n57134, n57135, n57136, n57137, n57138, n57139, n57140, n57141, n57142, n57143, n57144, n57145, n57146, n57147, n57148, n57149, n57150, n57151, n57152, n57153, n57154, n57155, n57156, n57157, n57158, n57159, n57160, n57161, n57162, n57163, n57164, n57165, n57166, n57167, n57168, n57169, n57170, n57171, n57172, n57173, n57174, n57175, n57176, n57177, n57178, n57179, n57180, n57181, n57182, n57183, n57184, n57185, n57186, n57187, n57188, n57189, n57190, n57191, n57192, n57193, n57194, n57195, n57196, n57197, n57198, n57199, n57200, n57201, n57202, n57203, n57204, n57205, n57206, n57207, n57208, n57209, n57210, n57211, n57212, n57213, n57214, n57215, n57216, n57217, n57218, n57219, n57220, n57221, n57222, n57223, n57224, n57225, n57226, n57227, n57228, n57229, n57230, n57231, n57232, n57233, n57234, n57235, n57236, n57237, n57238, n57239, n57240, n57241, n57242, n57243, n57244, n57245, n57246, n57247, n57248, n57249, n57250, n57251, n57252, n57253, n57254, n57255, n57256, n57257, n57258, n57259, n57260, n57261, n57262, n57263, n57264, n57265, n57266, n57267, n57268, n57269, n57270, n57271, n57272, n57273, n57274, n57275, n57276, n57277, n57278, n57279, n57280, n57281, n57282, n57283, n57284, n57285, n57286, n57287, n57288, n57289, n57290, n57291, n57292, n57293, n57294, n57295, n57296, n57297, n57298, n57299, n57300, n57301, n57302, n57303, n57304, n57305, n57306, n57307, n57308, n57309, n57310, n57311, n57312, n57313, n57314, n57315, n57316, n57317, n57318, n57319, n57320, n57321, n57322, n57323, n57324, n57325, n57326, n57327, n57328, n57329, n57330, n57331, n57332, n57333, n57334, n57335, n57336, n57337, n57338, n57339, n57340, n57341, n57342, n57343, n57344, n57345, n57346, n57347, n57348, n57349, n57350, n57351, n57352, n57353, n57354, n57355, n57356, n57357, n57358, n57359, n57360, n57361, n57362, n57363, n57364, n57365, n57366, n57367, n57368, n57369, n57370, n57371, n57372, n57373, n57374, n57375, n57376, n57377, n57378, n57379, n57380, n57381, n57382, n57383, n57384, n57385, n57386, n57387, n57388, n57389, n57390, n57391, n57392, n57393, n57394, n57395, n57396, n57397, n57398, n57399, n57400, n57401, n57402, n57403, n57404, n57405, n57406, n57407, n57408, n57409, n57410, n57411, n57412, n57413, n57414, n57415, n57416, n57417, n57418, n57419, n57420, n57421, n57422, n57423, n57424, n57425, n57426, n57427, n57428, n57429, n57430, n57431, n57432, n57433, n57434, n57435, n57436, n57437, n57438, n57439, n57440, n57441, n57442, n57443, n57444, n57445, n57446, n57447, n57448, n57449, n57450, n57451, n57452, n57453, n57454, n57455, n57456, n57457, n57458, n57459, n57460, n57461, n57462, n57463, n57464, n57465, n57466, n57467, n57468, n57469, n57470, n57471, n57472, n57473, n57474, n57475, n57476, n57477, n57478, n57479, n57480, n57481, n57482, n57483, n57484, n57485, n57486, n57487, n57488, n57489, n57490, n57491, n57492, n57493, n57494, n57495, n57496, n57497, n57498, n57499, n57500, n57501, n57502, n57503, n57504, n57505, n57506, n57507, n57508, n57509, n57510, n57511, n57512, n57513, n57514, n57515, n57516, n57517, n57518, n57519, n57520, n57521, n57522, n57523, n57524, n57525, n57526, n57527, n57528, n57529, n57530, n57531, n57532, n57533, n57534, n57535, n57536, n57537, n57538, n57539, n57540, n57541, n57542, n57543, n57544, n57545, n57546, n57547, n57548, n57549, n57550, n57551, n57552, n57553, n57554, n57555, n57556, n57557, n57558, n57559, n57560, n57561, n57562, n57563, n57564, n57565, n57566, n57567, n57568, n57569, n57570, n57571, n57572, n57573, n57574, n57575, n57576, n57577, n57578, n57579, n57580, n57581, n57582, n57583, n57584, n57585, n57586, n57587, n57588, n57589, n57590, n57591, n57592, n57593, n57594, n57595, n57596, n57597, n57598, n57599, n57600, n57601, n57602, n57603, n57604, n57605, n57606, n57607, n57608, n57609, n57610, n57611, n57612, n57613, n57614, n57615, n57616, n57617, n57618, n57619, n57620, n57621, n57622, n57623, n57624, n57625, n57626, n57627, n57628, n57629, n57630, n57631, n57632, n57633, n57634, n57635, n57636, n57637, n57638, n57639, n57640, n57641, n57642, n57643, n57644, n57645, n57646, n57647, n57648, n57649, n57650, n57651, n57652, n57653, n57654, n57655, n57656, n57657, n57658, n57659, n57660, n57661, n57662, n57663, n57664, n57665, n57666, n57667, n57668, n57669, n57670, n57671, n57672, n57673, n57674, n57675, n57676, n57677, n57678, n57679, n57680, n57681, n57682, n57683, n57684, n57685, n57686, n57687, n57688, n57689, n57690, n57691, n57692, n57693, n57694, n57695, n57696, n57697, n57698, n57699, n57700, n57701, n57702, n57703, n57704, n57705, n57706, n57707, n57708, n57709, n57710, n57711, n57712, n57713, n57714, n57715, n57716, n57717, n57718, n57719, n57720, n57721, n57722, n57723, n57724, n57725, n57726, n57727, n57728, n57729, n57730, n57731, n57732, n57733, n57734, n57735, n57736, n57737, n57738, n57739, n57740, n57741, n57742, n57743, n57744, n57745, n57746, n57747, n57748, n57749, n57750, n57751, n57752, n57753, n57754, n57755, n57756, n57757, n57758, n57759, n57760, n57761, n57762, n57763, n57764, n57765, n57766, n57767, n57768, n57769, n57770, n57771, n57772, n57773, n57774, n57775, n57776, n57777, n57778, n57779, n57780, n57781, n57782, n57783, n57784, n57785, n57786, n57787, n57788, n57789, n57790, n57791, n57792, n57793, n57794, n57795, n57796, n57797, n57798, n57799, n57800, n57801, n57802, n57803, n57804, n57805, n57806, n57807, n57808, n57809, n57810, n57811, n57812, n57813, n57814, n57815, n57816, n57817, n57818, n57819, n57820, n57821, n57822, n57823, n57824, n57825, n57826, n57827, n57828, n57829, n57830, n57831, n57832, n57833, n57834, n57835, n57836, n57837, n57838, n57839, n57840, n57841, n57842, n57843, n57844, n57845, n57846, n57847, n57848, n57849, n57850, n57851, n57852, n57853, n57854, n57855, n57856, n57857, n57858, n57859, n57860, n57861, n57862, n57863, n57864, n57865, n57866, n57867, n57868, n57869, n57870, n57871, n57872, n57873, n57874, n57875, n57876, n57877, n57878, n57879, n57880, n57881, n57882, n57883, n57884, n57885, n57886, n57887, n57888, n57889, n57890, n57891, n57892, n57893, n57894, n57895, n57896, n57897, n57898, n57899, n57900, n57901, n57902, n57903, n57904, n57905, n57906, n57907, n57908, n57909, n57910, n57911, n57912, n57913, n57914, n57915, n57916, n57917, n57918, n57919, n57920, n57921, n57922, n57923, n57924, n57925, n57926, n57927, n57928, n57929, n57930, n57931, n57932, n57933, n57934, n57935, n57936, n57937, n57938, n57939, n57940, n57941, n57942, n57943, n57944, n57945, n57946, n57947, n57948, n57949, n57950, n57951, n57952, n57953, n57954, n57955, n57956, n57957, n57958, n57959, n57960, n57961, n57962, n57963, n57964, n57965, n57966, n57967, n57968, n57969, n57970, n57971, n57972, n57973, n57974, n57975, n57976, n57977, n57978, n57979, n57980, n57981, n57982, n57983, n57984, n57985, n57986, n57987, n57988, n57989, n57990, n57991, n57992, n57993, n57994, n57995, n57996, n57997, n57998, n57999, n58000, n58001, n58002, n58003, n58004, n58005, n58006, n58007, n58008, n58009, n58010, n58011, n58012, n58013, n58014, n58015, n58016, n58017, n58018, n58019, n58020, n58021, n58022, n58023, n58024, n58025, n58026, n58027, n58028, n58029, n58030, n58031, n58032, n58033, n58034, n58035, n58036, n58037, n58038, n58039, n58040, n58041, n58042, n58043, n58044, n58045, n58046, n58047, n58048, n58049, n58050, n58051, n58052, n58053, n58054, n58055, n58056, n58057, n58058, n58059, n58060, n58061, n58062, n58063, n58064, n58065, n58066, n58067, n58068, n58069, n58070, n58071, n58072, n58073, n58074, n58075, n58076, n58077, n58078, n58079, n58080, n58081, n58082, n58083, n58084, n58085, n58086, n58087, n58088, n58089, n58090, n58091, n58092, n58093, n58094, n58095, n58096, n58097, n58098, n58099, n58100, n58101, n58102, n58103, n58104, n58105, n58106, n58107, n58108, n58109, n58110, n58111, n58112, n58113, n58114, n58115, n58116, n58117, n58118, n58119, n58120, n58121, n58122, n58123, n58124, n58125, n58126, n58127, n58128, n58129, n58130, n58131, n58132, n58133, n58134, n58135, n58136, n58137, n58138, n58139, n58140, n58141, n58142, n58143, n58144, n58145, n58146, n58147, n58148, n58149, n58150, n58151, n58152, n58153, n58154, n58155, n58156, n58157, n58158, n58159, n58160, n58161, n58162, n58163, n58164, n58165, n58166, n58167, n58168, n58169, n58170, n58171, n58172, n58173, n58174, n58175, n58176, n58177, n58178, n58179, n58180, n58181, n58182, n58183, n58184, n58185, n58186, n58187, n58188, n58189, n58190, n58191, n58192, n58193, n58194, n58195, n58196, n58197, n58198, n58199, n58200, n58201, n58202, n58203, n58204, n58205, n58206, n58207, n58208, n58209, n58210, n58211, n58212, n58213, n58214, n58215, n58216, n58217, n58218, n58219, n58220, n58221, n58222, n58223, n58224, n58225, n58226, n58227, n58228, n58229, n58230, n58231, n58232, n58233, n58234, n58235, n58236, n58237, n58238, n58239, n58240, n58241, n58242, n58243, n58244, n58245, n58246, n58247, n58248, n58249, n58250, n58251, n58252, n58253, n58254, n58255, n58256, n58257, n58258, n58259, n58260, n58261, n58262, n58263, n58264, n58265, n58266, n58267, n58268, n58269, n58270, n58271, n58272, n58273, n58274, n58275, n58276, n58277, n58278, n58279, n58280, n58281, n58282, n58283, n58284, n58285, n58286, n58287, n58288, n58289, n58290, n58291, n58292, n58293, n58294, n58295, n58296, n58297, n58298, n58299, n58300, n58301, n58302, n58303, n58304, n58305, n58306, n58307, n58308, n58309, n58310, n58311, n58312, n58313, n58314, n58315, n58316, n58317, n58318, n58319, n58320, n58321, n58322, n58323, n58324, n58325, n58326, n58327, n58328, n58329, n58330, n58331, n58332, n58333, n58334, n58335, n58336, n58337, n58338, n58339, n58340, n58341, n58342, n58343, n58344, n58345, n58346, n58347, n58348, n58349, n58350, n58351, n58352, n58353, n58354, n58355, n58356, n58357, n58358, n58359, n58360, n58361, n58362, n58363, n58364, n58365, n58366, n58367, n58368, n58369, n58370, n58371, n58372, n58373, n58374, n58375, n58376, n58377, n58378, n58379, n58380, n58381, n58382, n58383, n58384, n58385, n58386, n58387, n58388, n58389, n58390, n58391, n58392, n58393, n58394, n58395, n58396, n58397, n58398, n58399, n58400, n58401, n58402, n58403, n58404, n58405, n58406, n58407, n58408, n58409, n58410, n58411, n58412, n58413, n58414, n58415, n58416, n58417, n58418, n58419, n58420, n58421, n58422, n58423, n58424, n58425, n58426, n58427, n58428, n58429, n58430, n58431, n58432, n58433, n58434, n58435, n58436, n58437, n58438, n58439, n58440, n58441, n58442, n58443, n58444, n58445, n58446, n58447, n58448, n58449, n58450, n58451, n58452, n58453, n58454, n58455, n58456, n58457, n58458, n58459, n58460, n58461, n58462, n58463, n58464, n58465, n58466, n58467, n58468, n58469, n58470, n58471, n58472, n58473, n58474, n58475, n58476, n58477, n58478, n58479, n58480, n58481, n58482, n58483, n58484, n58485, n58486, n58487, n58488, n58489, n58490, n58491, n58492, n58493, n58494, n58495, n58496, n58497, n58498, n58499, n58500, n58501, n58502, n58503, n58504, n58505, n58506, n58507, n58508, n58509, n58510, n58511, n58512, n58513, n58514, n58515, n58516, n58517, n58518, n58519, n58520, n58521, n58522, n58523, n58524, n58525, n58526, n58527, n58528, n58529, n58530, n58531, n58532, n58533, n58534, n58535, n58536, n58537, n58538, n58539, n58540, n58541, n58542, n58543, n58544, n58545, n58546, n58547, n58548, n58549, n58550, n58551, n58552, n58553, n58554, n58555, n58556, n58557, n58558, n58559, n58560, n58561, n58562, n58563, n58564, n58565, n58566, n58567, n58568, n58569, n58570, n58571, n58572, n58573, n58574, n58575, n58576, n58577, n58578, n58579, n58580, n58581, n58582, n58583, n58584, n58585, n58586, n58587, n58588, n58589, n58590, n58591, n58592, n58593, n58594, n58595, n58596, n58597, n58598, n58599, n58600, n58601, n58602, n58603, n58604, n58605, n58606, n58607, n58608, n58609, n58610, n58611, n58612, n58613, n58614, n58615, n58616, n58617, n58618, n58619, n58620, n58621, n58622, n58623, n58624, n58625, n58626, n58627, n58628, n58629, n58630, n58631, n58632, n58633, n58634, n58635, n58636, n58637, n58638, n58639, n58640, n58641, n58642, n58643, n58644, n58645, n58646, n58647, n58648, n58649, n58650, n58651, n58652, n58653, n58654, n58655, n58656, n58657, n58658, n58659, n58660, n58661, n58662, n58663, n58664, n58665, n58666, n58667, n58668, n58669, n58670, n58671, n58672, n58673, n58674, n58675, n58676, n58677, n58678, n58679, n58680, n58681, n58682, n58683, n58684, n58685, n58686, n58687, n58688, n58689, n58690, n58691, n58692, n58693, n58694, n58695, n58696, n58697, n58698, n58699, n58700, n58701, n58702, n58703, n58704, n58705, n58706, n58707, n58708, n58709, n58710, n58711, n58712, n58713, n58714, n58715, n58716, n58717, n58718, n58719, n58720, n58721, n58722, n58723, n58724, n58725, n58726, n58727, n58728, n58729, n58730, n58731, n58732, n58733, n58734, n58735, n58736, n58737, n58738, n58739, n58740, n58741, n58742, n58743, n58744, n58745, n58746, n58747, n58748, n58749, n58750, n58751, n58752, n58753, n58754, n58755, n58756, n58757, n58758, n58759, n58760, n58761, n58762, n58763, n58764, n58765, n58766, n58767, n58768, n58769, n58770, n58771, n58772, n58773, n58774, n58775, n58776, n58777, n58778, n58779, n58780, n58781, n58782, n58783, n58784, n58785, n58786, n58787, n58788, n58789, n58790, n58791, n58792, n58793, n58794, n58795, n58796, n58797, n58798, n58799, n58800, n58801, n58802, n58803, n58804, n58805, n58806, n58807, n58808, n58809, n58810, n58811, n58812, n58813, n58814, n58815, n58816, n58817, n58818, n58819, n58820, n58821, n58822, n58823, n58824, n58825, n58826, n58827, n58828, n58829, n58830, n58831, n58832, n58833, n58834, n58835, n58836, n58837, n58838, n58839, n58840, n58841, n58842, n58843, n58844, n58845, n58846, n58847, n58848, n58849, n58850, n58851, n58852, n58853, n58854, n58855, n58856, n58857, n58858, n58859, n58860, n58861, n58862, n58863, n58864, n58865, n58866, n58867, n58868, n58869, n58870, n58871, n58872, n58873, n58874, n58875, n58876, n58877, n58878, n58879, n58880, n58881, n58882, n58883, n58884, n58885, n58886, n58887, n58888, n58889, n58890, n58891, n58892, n58893, n58894, n58895, n58896, n58897, n58898, n58899, n58900, n58901, n58902, n58903, n58904, n58905, n58906, n58907, n58908, n58909, n58910, n58911, n58912, n58913, n58914, n58915, n58916, n58917, n58918, n58919, n58920, n58921, n58922, n58923, n58924, n58925, n58926, n58927, n58928, n58929, n58930, n58931, n58932, n58933, n58934, n58935, n58936, n58937, n58938, n58939, n58940, n58941, n58942, n58943, n58944, n58945, n58946, n58947, n58948, n58949, n58950, n58951, n58952, n58953, n58954, n58955, n58956, n58957, n58958, n58959, n58960, n58961, n58962, n58963, n58964, n58965, n58966, n58967, n58968, n58969, n58970, n58971, n58972, n58973, n58974, n58975, n58976, n58977, n58978, n58979, n58980, n58981, n58982, n58983, n58984, n58985, n58986, n58987, n58988, n58989, n58990, n58991, n58992, n58993, n58994, n58995, n58996, n58997, n58998, n58999, n59000, n59001, n59002, n59003, n59004, n59005, n59006, n59007, n59008, n59009, n59010, n59011, n59012, n59013, n59014, n59015, n59016, n59017, n59018, n59019, n59020, n59021, n59022, n59023, n59024, n59025, n59026, n59027, n59028, n59029, n59030, n59031, n59032, n59033, n59034, n59035, n59036, n59037, n59038, n59039, n59040, n59041, n59042, n59043, n59044, n59045, n59046, n59047, n59048, n59049, n59050, n59051, n59052, n59053, n59054, n59055, n59056, n59057, n59058, n59059, n59060, n59061, n59062, n59063, n59064, n59065, n59066, n59067, n59068, n59069, n59070, n59071, n59072, n59073, n59074, n59075, n59076, n59077, n59078, n59079, n59080, n59081, n59082, n59083, n59084, n59085, n59086, n59087, n59088, n59089, n59090, n59091, n59092, n59093, n59094, n59095, n59096, n59097, n59098, n59099, n59100, n59101, n59102, n59103, n59104, n59105, n59106, n59107, n59108, n59109, n59110, n59111, n59112, n59113, n59114, n59115, n59116, n59117, n59118, n59119, n59120, n59121, n59122, n59123, n59124, n59125, n59126, n59127, n59128, n59129, n59130, n59131, n59132, n59133, n59134, n59135, n59136, n59137, n59138, n59139, n59140, n59141, n59142, n59143, n59144, n59145, n59146, n59147, n59148, n59149, n59150, n59151, n59152, n59153, n59154, n59155, n59156, n59157, n59158, n59159, n59160, n59161, n59162, n59163, n59164, n59165, n59166, n59167, n59168, n59169, n59170, n59171, n59172, n59173, n59174, n59175, n59176, n59177, n59178, n59179, n59180, n59181, n59182, n59183, n59184, n59185, n59186, n59187, n59188, n59189, n59190, n59191, n59192, n59193, n59194, n59195, n59196, n59197, n59198, n59199, n59200, n59201, n59202, n59203, n59204, n59205, n59206, n59207, n59208, n59209, n59210, n59211, n59212, n59213, n59214, n59215, n59216, n59217, n59218, n59219, n59220, n59221, n59222, n59223, n59224, n59225, n59226, n59227, n59228, n59229, n59230, n59231, n59232, n59233, n59234, n59235, n59236, n59237, n59238, n59239, n59240, n59241, n59242, n59243, n59244, n59245, n59246, n59247, n59248, n59249, n59250, n59251, n59252, n59253, n59254, n59255, n59256, n59257, n59258, n59259, n59260, n59261, n59262, n59263, n59264, n59265, n59266, n59267, n59268, n59269, n59270, n59271, n59272, n59273, n59274, n59275, n59276, n59277, n59278, n59279, n59280, n59281, n59282, n59283, n59284, n59285, n59286, n59287, n59288, n59289, n59290, n59291, n59292, n59293, n59294, n59295, n59296, n59297, n59298, n59299, n59300, n59301, n59302, n59303, n59304, n59305, n59306, n59307, n59308, n59309, n59310, n59311, n59312, n59313, n59314, n59315, n59316, n59317, n59318, n59319, n59320, n59321, n59322, n59323, n59324, n59325, n59326, n59327, n59328, n59329, n59330, n59331, n59332, n59333, n59334, n59335, n59336, n59337, n59338, n59339, n59340, n59341, n59342, n59343, n59344, n59345, n59346, n59347, n59348, n59349, n59350, n59351, n59352, n59353, n59354, n59355, n59356, n59357, n59358, n59359, n59360, n59361, n59362, n59363, n59364, n59365, n59366, n59367, n59368, n59369, n59370, n59371, n59372, n59373, n59374, n59375, n59376, n59377, n59378, n59379, n59380, n59381, n59382, n59383, n59384, n59385, n59386, n59387, n59388, n59389, n59390, n59391, n59392, n59393, n59394, n59395, n59396, n59397, n59398, n59399, n59400, n59401, n59402, n59403, n59404, n59405, n59406, n59407, n59408, n59409, n59410, n59411, n59412, n59413, n59414, n59415, n59416, n59417, n59418, n59419, n59420, n59421, n59422, n59423, n59424, n59425, n59426, n59427, n59428, n59429, n59430, n59431, n59432, n59433, n59434, n59435, n59436, n59437, n59438, n59439, n59440, n59441, n59442, n59443, n59444, n59445, n59446, n59447, n59448, n59449, n59450, n59451, n59452, n59453, n59454, n59455, n59456, n59457, n59458, n59459, n59460, n59461, n59462, n59463, n59464, n59465, n59466, n59467, n59468, n59469, n59470, n59471, n59472, n59473, n59474, n59475, n59476, n59477, n59478, n59479, n59480, n59481, n59482, n59483, n59484, n59485, n59486, n59487, n59488, n59489, n59490, n59491, n59492, n59493, n59494, n59495, n59496, n59497, n59498, n59499, n59500, n59501, n59502, n59503, n59504, n59505, n59506, n59507, n59508, n59509, n59510, n59511, n59512, n59513, n59514, n59515, n59516, n59517, n59518, n59519, n59520, n59521, n59522, n59523, n59524, n59525, n59526, n59527, n59528, n59529, n59530, n59531, n59532, n59533, n59534, n59535, n59536, n59537, n59538, n59539, n59540, n59541, n59542, n59543, n59544, n59545, n59546, n59547, n59548, n59549, n59550, n59551, n59552, n59553, n59554, n59555, n59556, n59557, n59558, n59559, n59560, n59561, n59562, n59563, n59564, n59565, n59566, n59567, n59568, n59569, n59570, n59571, n59572, n59573, n59574, n59575, n59576, n59577, n59578, n59579, n59580, n59581, n59582, n59583, n59584, n59585, n59586, n59587, n59588, n59589, n59590, n59591, n59592, n59593, n59594, n59595, n59596, n59597, n59598, n59599, n59600, n59601, n59602, n59603, n59604, n59605, n59606, n59607, n59608, n59609, n59610, n59611, n59612, n59613, n59614, n59615, n59616, n59617, n59618, n59619, n59620, n59621, n59622, n59623, n59624, n59625, n59626, n59627, n59628, n59629, n59630, n59631, n59632, n59633, n59634, n59635, n59636, n59637, n59638, n59639, n59640, n59641, n59642, n59643, n59644, n59645, n59646, n59647, n59648, n59649, n59650, n59651, n59652, n59653, n59654, n59655, n59656, n59657, n59658, n59659, n59660, n59661, n59662, n59663, n59664, n59665, n59666, n59667, n59668, n59669, n59670, n59671, n59672, n59673, n59674, n59675, n59676, n59677, n59678, n59679, n59680, n59681, n59682, n59683, n59684, n59685, n59686, n59687, n59688, n59689, n59690, n59691, n59692, n59693, n59694, n59695, n59696, n59697, n59698, n59699, n59700, n59701, n59702, n59703, n59704, n59705, n59706, n59707, n59708, n59709, n59710, n59711, n59712, n59713, n59714, n59715, n59716, n59717, n59718, n59719, n59720, n59721, n59722, n59723, n59724, n59725, n59726, n59727, n59728, n59729, n59730, n59731, n59732, n59733, n59734, n59735, n59736, n59737, n59738, n59739, n59740, n59741, n59742, n59743, n59744, n59745, n59746, n59747, n59748, n59749, n59750, n59751, n59752, n59753, n59754, n59755, n59756, n59757, n59758, n59759, n59760, n59761, n59762, n59763, n59764, n59765, n59766, n59767, n59768, n59769, n59770, n59771, n59772, n59773, n59774, n59775, n59776, n59777, n59778, n59779, n59780, n59781, n59782, n59783, n59784, n59785, n59786, n59787, n59788, n59789, n59790, n59791, n59792, n59793, n59794, n59795, n59796, n59797, n59798, n59799, n59800, n59801, n59802, n59803, n59804, n59805, n59806, n59807, n59808, n59809, n59810, n59811, n59812, n59813, n59814, n59815, n59816, n59817, n59818, n59819, n59820, n59821, n59822, n59823, n59824, n59825, n59826, n59827, n59828, n59829, n59830, n59831, n59832, n59833, n59834, n59835, n59836, n59837, n59838, n59839, n59840, n59841, n59842, n59843, n59844, n59845, n59846, n59847, n59848, n59849, n59850, n59851, n59852, n59853, n59854, n59855, n59856, n59857, n59858, n59859, n59860, n59861, n59862, n59863, n59864, n59865, n59866, n59867, n59868, n59869, n59870, n59871, n59872, n59873, n59874, n59875, n59876, n59877, n59878, n59879, n59880, n59881, n59882, n59883, n59884, n59885, n59886, n59887, n59888, n59889, n59890, n59891, n59892, n59893, n59894, n59895, n59896, n59897, n59898, n59899, n59900, n59901, n59902, n59903, n59904, n59905, n59906, n59907, n59908, n59909, n59910, n59911, n59912, n59913, n59914, n59915, n59916, n59917, n59918, n59919, n59920, n59921, n59922, n59923, n59924, n59925, n59926, n59927, n59928, n59929, n59930, n59931, n59932, n59933, n59934, n59935, n59936, n59937, n59938, n59939, n59940, n59941, n59942, n59943, n59944, n59945, n59946, n59947, n59948, n59949, n59950, n59951, n59952, n59953, n59954, n59955, n59956, n59957, n59958, n59959, n59960, n59961, n59962, n59963, n59964, n59965, n59966, n59967, n59968, n59969, n59970, n59971, n59972, n59973, n59974, n59975, n59976, n59977, n59978, n59979, n59980, n59981, n59982, n59983, n59984, n59985, n59986, n59987, n59988, n59989, n59990, n59991, n59992, n59993, n59994, n59995, n59996, n59997, n59998, n59999, n60000, n60001, n60002, n60003, n60004, n60005, n60006, n60007, n60008, n60009, n60010, n60011, n60012, n60013, n60014, n60015, n60016, n60017, n60018, n60019, n60020, n60021, n60022, n60023, n60024, n60025, n60026, n60027, n60028, n60029, n60030, n60031, n60032, n60033, n60034, n60035, n60036, n60037, n60038, n60039, n60040, n60041, n60042, n60043, n60044, n60045, n60046, n60047, n60048, n60049, n60050, n60051, n60052, n60053, n60054, n60055, n60056, n60057, n60058, n60059, n60060, n60061, n60062, n60063, n60064, n60065, n60066, n60067, n60068, n60069, n60070, n60071, n60072, n60073, n60074, n60075, n60076, n60077, n60078, n60079, n60080, n60081, n60082, n60083, n60084, n60085, n60086, n60087, n60088, n60089, n60090, n60091, n60092, n60093, n60094, n60095, n60096, n60097, n60098, n60099, n60100, n60101, n60102, n60103, n60104, n60105, n60106, n60107, n60108, n60109, n60110, n60111, n60112, n60113, n60114, n60115, n60116, n60117, n60118, n60119, n60120, n60121, n60122, n60123, n60124, n60125, n60126, n60127, n60128, n60129, n60130, n60131, n60132, n60133, n60134, n60135, n60136, n60137, n60138, n60139, n60140, n60141, n60142, n60143, n60144, n60145, n60146, n60147, n60148, n60149, n60150, n60151, n60152, n60153, n60154, n60155, n60156, n60157, n60158, n60159, n60160, n60161, n60162, n60163, n60164, n60165, n60166, n60167, n60168, n60169, n60170, n60171, n60172, n60173, n60174, n60175, n60176, n60177, n60178, n60179, n60180, n60181, n60182, n60183, n60184, n60185, n60186, n60187, n60188, n60189, n60190, n60191, n60192, n60193, n60194, n60195, n60196, n60197, n60198, n60199, n60200, n60201, n60202, n60203, n60204, n60205, n60206, n60207, n60208, n60209, n60210, n60211, n60212, n60213, n60214, n60215, n60216, n60217, n60218, n60219, n60220, n60221, n60222, n60223, n60224, n60225, n60226, n60227, n60228, n60229, n60230, n60231, n60232, n60233, n60234, n60235, n60236, n60237, n60238, n60239, n60240, n60241, n60242, n60243, n60244, n60245, n60246, n60247, n60248, n60249, n60250, n60251, n60252, n60253, n60254, n60255, n60256, n60257, n60258, n60259, n60260, n60261, n60262, n60263, n60264, n60265, n60266, n60267, n60268, n60269, n60270, n60271, n60272, n60273, n60274, n60275, n60276, n60277, n60278, n60279, n60280, n60281, n60282, n60283, n60284, n60285, n60286, n60287, n60288, n60289, n60290, n60291, n60292, n60293, n60294, n60295, n60296, n60297, n60298, n60299, n60300, n60301, n60302, n60303, n60304, n60305, n60306, n60307, n60308, n60309, n60310, n60311, n60312, n60313, n60314, n60315, n60316, n60317, n60318, n60319, n60320, n60321, n60322, n60323, n60324, n60325, n60326, n60327, n60328, n60329, n60330, n60331, n60332, n60333, n60334, n60335, n60336, n60337, n60338, n60339, n60340, n60341, n60342, n60343, n60344, n60345, n60346, n60347, n60348, n60349, n60350, n60351, n60352, n60353, n60354, n60355, n60356, n60357, n60358, n60359, n60360, n60361, n60362, n60363, n60364, n60365, n60366, n60367, n60368, n60369, n60370, n60371, n60372, n60373, n60374, n60375, n60376, n60377, n60378, n60379, n60380, n60381, n60382, n60383, n60384, n60385, n60386, n60387, n60388, n60389, n60390, n60391, n60392, n60393, n60394, n60395, n60396, n60397, n60398, n60399, n60400, n60401, n60402, n60403, n60404, n60405, n60406, n60407, n60408, n60409, n60410, n60411, n60412, n60413, n60414, n60415, n60416, n60417, n60418, n60419, n60420, n60421, n60422, n60423, n60424, n60425, n60426, n60427, n60428, n60429, n60430, n60431, n60432, n60433, n60434, n60435, n60436, n60437, n60438, n60439, n60440, n60441, n60442, n60443, n60444, n60445, n60446, n60447, n60448, n60449, n60450, n60451, n60452, n60453, n60454, n60455, n60456, n60457, n60458, n60459, n60460, n60461, n60462, n60463, n60464, n60465, n60466, n60467, n60468, n60469, n60470, n60471, n60472, n60473, n60474, n60475, n60476, n60477, n60478, n60479, n60480, n60481, n60482, n60483, n60484, n60485, n60486, n60487, n60488, n60489, n60490, n60491, n60492, n60493, n60494, n60495, n60496, n60497, n60498, n60499, n60500, n60501, n60502, n60503, n60504, n60505, n60506, n60507, n60508, n60509, n60510, n60511, n60512, n60513, n60514, n60515, n60516, n60517, n60518, n60519, n60520, n60521, n60522, n60523, n60524, n60525, n60526, n60527, n60528, n60529, n60530, n60531, n60532, n60533, n60534, n60535, n60536, n60537, n60538, n60539, n60540, n60541, n60542, n60543, n60544, n60545, n60546, n60547, n60548, n60549, n60550, n60551, n60552, n60553, n60554, n60555, n60556, n60557, n60558, n60559, n60560, n60561, n60562, n60563, n60564, n60565, n60566, n60567, n60568, n60569, n60570, n60571, n60572, n60573, n60574, n60575, n60576, n60577, n60578, n60579, n60580, n60581, n60582, n60583, n60584, n60585, n60586, n60587, n60588, n60589, n60590, n60591, n60592, n60593, n60594, n60595, n60596, n60597, n60598, n60599, n60600, n60601, n60602, n60603, n60604, n60605, n60606, n60607, n60608, n60609, n60610, n60611, n60612, n60613, n60614, n60615, n60616, n60617, n60618, n60619, n60620, n60621, n60622, n60623, n60624, n60625, n60626, n60627, n60628, n60629, n60630, n60631, n60632, n60633, n60634, n60635, n60636, n60637, n60638, n60639, n60640, n60641, n60642, n60643, n60644, n60645, n60646, n60647, n60648, n60649, n60650, n60651, n60652, n60653, n60654, n60655, n60656, n60657, n60658, n60659, n60660, n60661, n60662, n60663, n60664, n60665, n60666, n60667, n60668, n60669, n60670, n60671, n60672, n60673, n60674, n60675, n60676, n60677, n60678, n60679, n60680, n60681, n60682, n60683, n60684, n60685, n60686, n60687, n60688, n60689, n60690, n60691, n60692, n60693, n60694, n60695, n60696, n60697, n60698, n60699, n60700, n60701, n60702, n60703, n60704, n60705, n60706, n60707, n60708, n60709, n60710, n60711, n60712, n60713, n60714, n60715, n60716, n60717, n60718, n60719, n60720, n60721, n60722, n60723, n60724, n60725, n60726, n60727, n60728, n60729, n60730, n60731, n60732, n60733, n60734, n60735, n60736, n60737, n60738, n60739, n60740, n60741, n60742, n60743, n60744, n60745, n60746, n60747, n60748, n60749, n60750, n60751, n60752, n60753, n60754, n60755, n60756, n60757, n60758, n60759, n60760, n60761, n60762, n60763, n60764, n60765, n60766, n60767, n60768, n60769, n60770, n60771, n60772, n60773, n60774, n60775, n60776, n60777, n60778, n60779, n60780, n60781, n60782, n60783, n60784, n60785, n60786, n60787, n60788, n60789, n60790, n60791, n60792, n60793, n60794, n60795, n60796, n60797, n60798, n60799, n60800, n60801, n60802, n60803, n60804, n60805, n60806, n60807, n60808, n60809, n60810, n60811, n60812, n60813, n60814, n60815, n60816, n60817, n60818, n60819, n60820, n60821, n60822, n60823, n60824, n60825, n60826, n60827, n60828, n60829, n60830, n60831, n60832, n60833, n60834, n60835, n60836, n60837, n60838, n60839, n60840, n60841, n60842, n60843, n60844, n60845, n60846, n60847, n60848, n60849, n60850, n60851, n60852, n60853, n60854, n60855, n60856, n60857, n60858, n60859, n60860, n60861, n60862, n60863, n60864, n60865, n60866, n60867, n60868, n60869, n60870, n60871, n60872, n60873, n60874, n60875, n60876, n60877, n60878, n60879, n60880, n60881, n60882, n60883, n60884, n60885, n60886, n60887, n60888, n60889, n60890, n60891, n60892, n60893, n60894, n60895, n60896, n60897, n60898, n60899, n60900, n60901, n60902, n60903, n60904, n60905, n60906, n60907, n60908, n60909, n60910, n60911, n60912, n60913, n60914, n60915, n60916, n60917, n60918, n60919, n60920, n60921, n60922, n60923, n60924, n60925, n60926, n60927, n60928, n60929, n60930, n60931, n60932, n60933, n60934, n60935, n60936, n60937, n60938, n60939, n60940, n60941, n60942, n60943, n60944, n60945, n60946, n60947, n60948, n60949, n60950, n60951, n60952, n60953, n60954, n60955, n60956, n60957, n60958, n60959, n60960, n60961, n60962, n60963, n60964, n60965, n60966, n60967, n60968, n60969, n60970, n60971, n60972, n60973, n60974, n60975, n60976, n60977, n60978, n60979, n60980, n60981, n60982, n60983, n60984, n60985, n60986, n60987, n60988, n60989, n60990, n60991, n60992, n60993, n60994, n60995, n60996, n60997, n60998, n60999, n61000, n61001, n61002, n61003, n61004, n61005, n61006, n61007, n61008, n61009, n61010, n61011, n61012, n61013, n61014, n61015, n61016, n61017, n61018, n61019, n61020, n61021, n61022, n61023, n61024, n61025, n61026, n61027, n61028, n61029, n61030, n61031, n61032, n61033, n61034, n61035, n61036, n61037, n61038, n61039, n61040, n61041, n61042, n61043, n61044, n61045, n61046, n61047, n61048, n61049, n61050, n61051, n61052, n61053, n61054, n61055, n61056, n61057, n61058, n61059, n61060, n61061, n61062, n61063, n61064, n61065, n61066, n61067, n61068, n61069, n61070, n61071, n61072, n61073, n61074, n61075, n61076, n61077, n61078, n61079, n61080, n61081, n61082, n61083, n61084, n61085, n61086, n61087, n61088, n61089, n61090, n61091, n61092, n61093, n61094, n61095, n61096, n61097, n61098, n61099, n61100, n61101, n61102, n61103, n61104, n61105, n61106, n61107, n61108, n61109, n61110, n61111, n61112, n61113, n61114, n61115, n61116, n61117, n61118, n61119, n61120, n61121, n61122, n61123, n61124, n61125, n61126, n61127, n61128, n61129, n61130, n61131, n61132, n61133, n61134, n61135, n61136, n61137, n61138, n61139, n61140, n61141, n61142, n61143, n61144, n61145, n61146, n61147, n61148, n61149, n61150, n61151, n61152, n61153, n61154, n61155, n61156, n61157, n61158, n61159, n61160, n61161, n61162, n61163, n61164, n61165, n61166, n61167, n61168, n61169, n61170, n61171, n61172, n61173, n61174, n61175, n61176, n61177, n61178, n61179, n61180, n61181, n61182, n61183, n61184, n61185, n61186, n61187, n61188, n61189, n61190, n61191, n61192, n61193, n61194, n61195, n61196, n61197, n61198, n61199, n61200, n61201, n61202, n61203, n61204, n61205, n61206, n61207, n61208, n61209, n61210, n61211, n61212, n61213, n61214, n61215, n61216, n61217, n61218, n61219, n61220, n61221, n61222, n61223, n61224, n61225, n61226, n61227, n61228, n61229, n61230, n61231, n61232, n61233, n61234, n61235, n61236, n61237, n61238, n61239, n61240, n61241, n61242, n61243, n61244, n61245, n61246, n61247, n61248, n61249, n61250, n61251, n61252, n61253, n61254, n61255, n61256, n61257, n61258, n61259, n61260, n61261, n61262, n61263, n61264, n61265, n61266, n61267, n61268, n61269, n61270, n61271, n61272, n61273, n61274, n61275, n61276, n61277, n61278, n61279, n61280, n61281, n61282, n61283, n61284, n61285, n61286, n61287, n61288, n61289, n61290, n61291, n61292, n61293, n61294, n61295, n61296, n61297, n61298, n61299, n61300, n61301, n61302, n61303, n61304, n61305, n61306, n61307, n61308, n61309, n61310, n61311, n61312, n61313, n61314, n61315, n61316, n61317, n61318, n61319, n61320, n61321, n61322, n61323, n61324, n61325, n61326, n61327, n61328, n61329, n61330, n61331, n61332, n61333, n61334, n61335, n61336, n61337, n61338, n61339, n61340, n61341, n61342, n61343, n61344, n61345, n61346, n61347, n61348, n61349, n61350, n61351, n61352, n61353, n61354, n61355, n61356, n61357, n61358, n61359, n61360, n61361, n61362, n61363, n61364, n61365, n61366, n61367, n61368, n61369, n61370, n61371, n61372, n61373, n61374, n61375, n61376, n61377, n61378, n61379, n61380, n61381, n61382, n61383, n61384, n61385, n61386, n61387, n61388, n61389, n61390, n61391, n61392, n61393, n61394, n61395, n61396, n61397, n61398, n61399, n61400, n61401, n61402, n61403, n61404, n61405, n61406, n61407, n61408, n61409, n61410, n61411, n61412, n61413, n61414, n61415, n61416, n61417, n61418, n61419, n61420, n61421, n61422, n61423, n61424, n61425, n61426, n61427, n61428, n61429, n61430, n61431, n61432, n61433, n61434, n61435, n61436, n61437, n61438, n61439, n61440, n61441, n61442, n61443, n61444, n61445, n61446, n61447, n61448, n61449, n61450, n61451, n61452, n61453, n61454, n61455, n61456, n61457, n61458, n61459, n61460, n61461, n61462, n61463, n61464, n61465, n61466, n61467, n61468, n61469, n61470, n61471, n61472, n61473, n61474, n61475, n61476, n61477, n61478, n61479, n61480, n61481, n61482, n61483, n61484, n61485, n61486, n61487, n61488, n61489, n61490, n61491, n61492, n61493, n61494, n61495, n61496, n61497, n61498, n61499, n61500, n61501, n61502, n61503, n61504, n61505, n61506, n61507, n61508, n61509, n61510, n61511, n61512, n61513, n61514, n61515, n61516, n61517, n61518, n61519, n61520, n61521, n61522, n61523, n61524, n61525, n61526, n61527, n61528, n61529, n61530, n61531, n61532, n61533, n61534, n61535, n61536, n61537, n61538, n61539, n61540, n61541, n61542, n61543, n61544, n61545, n61546, n61547, n61548, n61549, n61550, n61551, n61552, n61553, n61554, n61555, n61556, n61557, n61558, n61559, n61560, n61561, n61562, n61563, n61564, n61565, n61566, n61567, n61568, n61569, n61570, n61571, n61572, n61573, n61574, n61575, n61576, n61577, n61578, n61579, n61580, n61581, n61582, n61583, n61584, n61585, n61586, n61587, n61588, n61589, n61590, n61591, n61592, n61593, n61594, n61595, n61596, n61597, n61598, n61599, n61600, n61601, n61602, n61603, n61604, n61605, n61606, n61607, n61608, n61609, n61610, n61611, n61612, n61613, n61614, n61615, n61616, n61617, n61618, n61619, n61620, n61621, n61622, n61623, n61624, n61625, n61626, n61627, n61628, n61629, n61630, n61631, n61632, n61633, n61634, n61635, n61636, n61637, n61638, n61639, n61640, n61641, n61642, n61643, n61644, n61645, n61646, n61647, n61648, n61649, n61650, n61651, n61652, n61653, n61654, n61655, n61656, n61657, n61658, n61659, n61660, n61661, n61662, n61663, n61664, n61665, n61666, n61667, n61668, n61669, n61670, n61671, n61672, n61673, n61674, n61675, n61676, n61677, n61678, n61679, n61680, n61681, n61682, n61683, n61684, n61685, n61686, n61687, n61688, n61689, n61690, n61691, n61692, n61693, n61694, n61695, n61696, n61697, n61698, n61699, n61700, n61701, n61702, n61703, n61704, n61705, n61706, n61707, n61708, n61709, n61710, n61711, n61712, n61713, n61714, n61715, n61716, n61717, n61718, n61719, n61720, n61721, n61722, n61723, n61724, n61725, n61726, n61727, n61728, n61729, n61730, n61731, n61732, n61733, n61734, n61735, n61736, n61737, n61738, n61739, n61740, n61741, n61742, n61743, n61744, n61745, n61746, n61747, n61748, n61749, n61750, n61751, n61752, n61753, n61754, n61755, n61756, n61757, n61758, n61759, n61760, n61761, n61762, n61763, n61764, n61765, n61766, n61767, n61768, n61769, n61770, n61771, n61772, n61773, n61774, n61775, n61776, n61777, n61778, n61779, n61780, n61781, n61782, n61783, n61784, n61785, n61786, n61787, n61788, n61789, n61790, n61791, n61792, n61793, n61794, n61795, n61796, n61797, n61798, n61799, n61800, n61801, n61802, n61803, n61804, n61805, n61806, n61807, n61808, n61809, n61810, n61811, n61812, n61813, n61814, n61815, n61816, n61817, n61818, n61819, n61820, n61821, n61822, n61823, n61824, n61825, n61826, n61827, n61828, n61829, n61830, n61831, n61832, n61833, n61834, n61835, n61836, n61837, n61838, n61839, n61840, n61841, n61842, n61843, n61844, n61845, n61846, n61847, n61848, n61849, n61850, n61851, n61852, n61853, n61854, n61855, n61856, n61857, n61858, n61859, n61860, n61861, n61862, n61863, n61864, n61865, n61866, n61867, n61868, n61869, n61870, n61871, n61872, n61873, n61874, n61875, n61876, n61877, n61878, n61879, n61880, n61881, n61882, n61883, n61884, n61885, n61886, n61887, n61888, n61889, n61890, n61891, n61892, n61893, n61894, n61895, n61896, n61897, n61898, n61899, n61900, n61901, n61902, n61903, n61904, n61905, n61906, n61907, n61908, n61909, n61910, n61911, n61912, n61913, n61914, n61915, n61916, n61917, n61918, n61919, n61920, n61921, n61922, n61923, n61924, n61925, n61926, n61927, n61928, n61929, n61930, n61931, n61932, n61933, n61934, n61935, n61936, n61937, n61938, n61939, n61940, n61941, n61942, n61943, n61944, n61945, n61946, n61947, n61948, n61949, n61950, n61951, n61952, n61953, n61954, n61955, n61956, n61957, n61958, n61959, n61960, n61961, n61962, n61963, n61964, n61965, n61966, n61967, n61968, n61969, n61970, n61971, n61972, n61973, n61974, n61975, n61976, n61977, n61978, n61979, n61980, n61981, n61982, n61983, n61984, n61985, n61986, n61987, n61988, n61989, n61990, n61991, n61992, n61993, n61994, n61995, n61996, n61997, n61998, n61999, n62000, n62001, n62002, n62003, n62004, n62005, n62006, n62007, n62008, n62009, n62010, n62011, n62012, n62013, n62014, n62015, n62016, n62017, n62018, n62019, n62020, n62021, n62022, n62023, n62024, n62025, n62026, n62027, n62028, n62029, n62030, n62031, n62032, n62033, n62034, n62035, n62036, n62037, n62038, n62039, n62040, n62041, n62042, n62043, n62044, n62045, n62046, n62047, n62048, n62049, n62050, n62051, n62052, n62053, n62054, n62055, n62056, n62057, n62058, n62059, n62060, n62061, n62062, n62063, n62064, n62065, n62066, n62067, n62068, n62069, n62070, n62071, n62072, n62073, n62074, n62075, n62076, n62077, n62078, n62079, n62080, n62081, n62082, n62083, n62084, n62085, n62086, n62087, n62088, n62089, n62090, n62091, n62092, n62093, n62094, n62095, n62096, n62097, n62098, n62099, n62100, n62101, n62102, n62103, n62104, n62105, n62106, n62107, n62108, n62109, n62110, n62111, n62112, n62113, n62114, n62115, n62116, n62117, n62118, n62119, n62120, n62121, n62122, n62123, n62124, n62125, n62126, n62127, n62128, n62129, n62130, n62131, n62132, n62133, n62134, n62135, n62136, n62137, n62138, n62139, n62140, n62141, n62142, n62143, n62144, n62145, n62146, n62147, n62148, n62149, n62150, n62151, n62152, n62153, n62154, n62155, n62156, n62157, n62158, n62159, n62160, n62161, n62162, n62163, n62164, n62165, n62166, n62167, n62168, n62169, n62170, n62171, n62172, n62173, n62174, n62175, n62176, n62177, n62178, n62179, n62180, n62181, n62182, n62183, n62184, n62185, n62186, n62187, n62188, n62189, n62190, n62191, n62192, n62193, n62194, n62195, n62196, n62197, n62198, n62199, n62200, n62201, n62202, n62203, n62204, n62205, n62206, n62207, n62208, n62209, n62210, n62211, n62212, n62213, n62214, n62215, n62216, n62217, n62218, n62219, n62220, n62221, n62222, n62223, n62224, n62225, n62226, n62227, n62228, n62229, n62230, n62231, n62232, n62233, n62234, n62235, n62236, n62237, n62238, n62239, n62240, n62241, n62242, n62243, n62244, n62245, n62246, n62247, n62248, n62249, n62250, n62251, n62252, n62253, n62254, n62255, n62256, n62257, n62258, n62259, n62260, n62261, n62262, n62263, n62264, n62265, n62266, n62267, n62268, n62269, n62270, n62271, n62272, n62273, n62274, n62275, n62276, n62277, n62278, n62279, n62280, n62281, n62282, n62283, n62284, n62285, n62286, n62287, n62288, n62289, n62290, n62291, n62292, n62293, n62294, n62295, n62296, n62297, n62298, n62299, n62300, n62301, n62302, n62303, n62304, n62305, n62306, n62307, n62308, n62309, n62310, n62311, n62312, n62313, n62314, n62315, n62316, n62317, n62318, n62319, n62320, n62321, n62322, n62323, n62324, n62325, n62326, n62327, n62328, n62329, n62330, n62331, n62332, n62333, n62334, n62335, n62336, n62337, n62338, n62339, n62340, n62341, n62342, n62343, n62344, n62345, n62346, n62347, n62348, n62349, n62350, n62351, n62352, n62353, n62354, n62355, n62356, n62357, n62358, n62359, n62360, n62361, n62362, n62363, n62364, n62365, n62366, n62367, n62368, n62369, n62370, n62371, n62372, n62373, n62374, n62375, n62376, n62377, n62378, n62379, n62380, n62381, n62382, n62383, n62384, n62385, n62386, n62387, n62388, n62389, n62390, n62391, n62392, n62393, n62394, n62395, n62396, n62397, n62398, n62399, n62400, n62401, n62402, n62403, n62404, n62405, n62406, n62407, n62408, n62409, n62410, n62411, n62412, n62413, n62414, n62415, n62416, n62417, n62418, n62419, n62420, n62421, n62422, n62423, n62424, n62425, n62426, n62427, n62428, n62429, n62430, n62431, n62432, n62433, n62434, n62435, n62436, n62437, n62438, n62439, n62440, n62441, n62442, n62443, n62444, n62445, n62446, n62447, n62448, n62449, n62450, n62451, n62452, n62453, n62454, n62455, n62456, n62457, n62458, n62459, n62460, n62461, n62462, n62463, n62464, n62465, n62466, n62467, n62468, n62469, n62470, n62471, n62472, n62473, n62474, n62475, n62476, n62477, n62478, n62479, n62480, n62481, n62482, n62483, n62484, n62485, n62486, n62487, n62488, n62489, n62490, n62491, n62492, n62493, n62494, n62495, n62496, n62497, n62498, n62499, n62500, n62501, n62502, n62503, n62504, n62505, n62506, n62507, n62508, n62509, n62510, n62511, n62512, n62513, n62514, n62515, n62516, n62517, n62518, n62519, n62520, n62521, n62522, n62523, n62524, n62525, n62526, n62527, n62528, n62529, n62530, n62531, n62532, n62533, n62534, n62535, n62536, n62537, n62538, n62539, n62540, n62541, n62542, n62543, n62544, n62545, n62546, n62547, n62548, n62549, n62550, n62551, n62552, n62553, n62554, n62555, n62556, n62557, n62558, n62559, n62560, n62561, n62562, n62563, n62564, n62565, n62566, n62567, n62568, n62569, n62570, n62571, n62572, n62573, n62574, n62575, n62576, n62577, n62578, n62579, n62580, n62581, n62582, n62583, n62584, n62585, n62586, n62587, n62588, n62589, n62590, n62591, n62592, n62593, n62594, n62595, n62596, n62597, n62598, n62599, n62600, n62601, n62602, n62603, n62604, n62605, n62606, n62607, n62608, n62609, n62610, n62611, n62612, n62613, n62614, n62615, n62616, n62617, n62618, n62619, n62620, n62621, n62622, n62623, n62624, n62625, n62626, n62627, n62628, n62629, n62630, n62631, n62632, n62633, n62634, n62635, n62636, n62637, n62638, n62639, n62640, n62641, n62642, n62643, n62644, n62645, n62646, n62647, n62648, n62649, n62650, n62651, n62652, n62653, n62654, n62655, n62656, n62657, n62658, n62659, n62660, n62661, n62662, n62663, n62664, n62665, n62666, n62667, n62668, n62669, n62670, n62671, n62672, n62673, n62674, n62675, n62676, n62677, n62678, n62679, n62680, n62681, n62682, n62683, n62684, n62685, n62686, n62687, n62688, n62689, n62690, n62691, n62692, n62693, n62694, n62695, n62696, n62697, n62698, n62699, n62700, n62701, n62702, n62703, n62704, n62705, n62706, n62707, n62708, n62709, n62710, n62711, n62712, n62713, n62714, n62715, n62716, n62717, n62718, n62719, n62720, n62721, n62722, n62723, n62724, n62725, n62726, n62727, n62728, n62729, n62730, n62731, n62732, n62733, n62734, n62735, n62736, n62737, n62738, n62739, n62740, n62741, n62742, n62743, n62744, n62745, n62746, n62747, n62748, n62749, n62750, n62751, n62752, n62753, n62754, n62755, n62756, n62757, n62758, n62759, n62760, n62761, n62762, n62763, n62764, n62765, n62766, n62767, n62768, n62769, n62770, n62771, n62772, n62773, n62774, n62775, n62776, n62777, n62778, n62779, n62780, n62781, n62782, n62783, n62784, n62785, n62786, n62787, n62788, n62789, n62790, n62791, n62792, n62793, n62794, n62795, n62796, n62797, n62798, n62799, n62800, n62801, n62802, n62803, n62804, n62805, n62806, n62807, n62808, n62809, n62810, n62811, n62812, n62813, n62814, n62815, n62816, n62817, n62818, n62819, n62820, n62821, n62822, n62823, n62824, n62825, n62826, n62827, n62828, n62829, n62830, n62831, n62832, n62833, n62834, n62835, n62836, n62837, n62838, n62839, n62840, n62841, n62842, n62843, n62844, n62845, n62846, n62847, n62848, n62849, n62850, n62851, n62852, n62853, n62854, n62855, n62856, n62857, n62858, n62859, n62860, n62861, n62862, n62863, n62864, n62865, n62866, n62867, n62868, n62869, n62870, n62871, n62872, n62873, n62874, n62875, n62876, n62877, n62878, n62879, n62880, n62881, n62882, n62883, n62884, n62885, n62886, n62887, n62888, n62889, n62890, n62891, n62892, n62893, n62894, n62895, n62896, n62897, n62898, n62899, n62900, n62901, n62902, n62903, n62904, n62905, n62906, n62907, n62908, n62909, n62910, n62911, n62912, n62913, n62914, n62915, n62916, n62917, n62918, n62919, n62920, n62921, n62922, n62923, n62924, n62925, n62926, n62927, n62928, n62929, n62930, n62931, n62932, n62933, n62934, n62935, n62936, n62937, n62938, n62939, n62940, n62941, n62942, n62943, n62944, n62945, n62946, n62947, n62948, n62949, n62950, n62951, n62952, n62953, n62954, n62955, n62956, n62957, n62958, n62959, n62960, n62961, n62962, n62963, n62964, n62965, n62966, n62967, n62968, n62969, n62970, n62971, n62972, n62973, n62974, n62975, n62976, n62977, n62978, n62979, n62980, n62981, n62982, n62983, n62984, n62985, n62986, n62987, n62988, n62989, n62990, n62991, n62992, n62993, n62994, n62995, n62996, n62997, n62998, n62999, n63000, n63001, n63002, n63003, n63004, n63005, n63006, n63007, n63008, n63009, n63010, n63011, n63012, n63013, n63014, n63015, n63016, n63017, n63018, n63019, n63020, n63021, n63022, n63023, n63024, n63025, n63026, n63027, n63028, n63029, n63030, n63031, n63032, n63033, n63034, n63035, n63036, n63037, n63038, n63039, n63040, n63041, n63042, n63043, n63044, n63045, n63046, n63047, n63048, n63049, n63050, n63051, n63052, n63053, n63054, n63055, n63056, n63057, n63058, n63059, n63060, n63061, n63062, n63063, n63064, n63065, n63066, n63067, n63068, n63069, n63070, n63071, n63072, n63073, n63074, n63075, n63076, n63077, n63078, n63079, n63080, n63081, n63082, n63083, n63084, n63085, n63086, n63087, n63088, n63089, n63090, n63091, n63092, n63093, n63094, n63095, n63096, n63097, n63098, n63099, n63100, n63101, n63102, n63103, n63104, n63105, n63106, n63107, n63108, n63109, n63110, n63111, n63112, n63113, n63114, n63115, n63116, n63117, n63118, n63119, n63120, n63121, n63122, n63123, n63124, n63125, n63126, n63127, n63128, n63129, n63130, n63131, n63132, n63133, n63134, n63135, n63136, n63137, n63138, n63139, n63140, n63141, n63142, n63143, n63144, n63145, n63146, n63147, n63148, n63149, n63150, n63151, n63152, n63153, n63154, n63155, n63156, n63157, n63158, n63159, n63160, n63161, n63162, n63163, n63164, n63165, n63166, n63167, n63168, n63169, n63170, n63171, n63172, n63173, n63174, n63175, n63176, n63177, n63178, n63179, n63180, n63181, n63182, n63183, n63184, n63185, n63186, n63187, n63188, n63189, n63190, n63191, n63192, n63193, n63194, n63195, n63196, n63197, n63198, n63199, n63200, n63201, n63202, n63203, n63204, n63205, n63206, n63207, n63208, n63209, n63210, n63211, n63212, n63213, n63214, n63215, n63216, n63217, n63218, n63219, n63220, n63221, n63222, n63223, n63224, n63225, n63226, n63227, n63228, n63229, n63230, n63231, n63232, n63233, n63234, n63235, n63236, n63237, n63238, n63239, n63240, n63241, n63242, n63243, n63244, n63245, n63246, n63247, n63248, n63249, n63250, n63251, n63252, n63253, n63254, n63255, n63256, n63257, n63258, n63259, n63260, n63261, n63262, n63263, n63264, n63265, n63266, n63267, n63268, n63269, n63270, n63271, n63272, n63273, n63274, n63275, n63276, n63277, n63278, n63279, n63280, n63281, n63282, n63283, n63284, n63285, n63286, n63287, n63288, n63289, n63290, n63291, n63292, n63293, n63294, n63295, n63296, n63297, n63298, n63299, n63300, n63301, n63302, n63303, n63304, n63305, n63306, n63307, n63308, n63309, n63310, n63311, n63312, n63313, n63314, n63315, n63316, n63317, n63318, n63319, n63320, n63321, n63322, n63323, n63324, n63325, n63326, n63327, n63328, n63329, n63330, n63331, n63332, n63333, n63334, n63335, n63336, n63337, n63338, n63339, n63340, n63341, n63342, n63343, n63344, n63345, n63346, n63347, n63348, n63349, n63350, n63351, n63352, n63353, n63354, n63355, n63356, n63357, n63358, n63359, n63360, n63361, n63362, n63363, n63364, n63365, n63366, n63367, n63368, n63369, n63370, n63371, n63372, n63373, n63374, n63375, n63376, n63377, n63378, n63379, n63380, n63381, n63382, n63383, n63384, n63385, n63386, n63387, n63388, n63389, n63390, n63391, n63392, n63393, n63394, n63395, n63396, n63397, n63398, n63399, n63400, n63401, n63402, n63403, n63404, n63405, n63406, n63407, n63408, n63409, n63410, n63411, n63412, n63413, n63414, n63415, n63416, n63417, n63418, n63419, n63420, n63421, n63422, n63423, n63424, n63425, n63426, n63427, n63428, n63429, n63430, n63431, n63432, n63433, n63434, n63435, n63436, n63437, n63438, n63439, n63440, n63441, n63442, n63443, n63444, n63445, n63446, n63447, n63448, n63449, n63450, n63451, n63452, n63453, n63454, n63455, n63456, n63457, n63458, n63459, n63460, n63461, n63462, n63463, n63464, n63465, n63466, n63467, n63468, n63469, n63470, n63471, n63472, n63473, n63474, n63475, n63476, n63477, n63478, n63479, n63480, n63481, n63482, n63483, n63484, n63485, n63486, n63487, n63488, n63489, n63490, n63491, n63492, n63493, n63494, n63495, n63496, n63497, n63498, n63499, n63500, n63501, n63502, n63503, n63504, n63505, n63506, n63507, n63508, n63509, n63510, n63511, n63512, n63513, n63514, n63515, n63516, n63517, n63518, n63519, n63520, n63521, n63522, n63523, n63524, n63525, n63526, n63527, n63528, n63529, n63530, n63531, n63532, n63533, n63534, n63535, n63536, n63537, n63538, n63539, n63540, n63541, n63542, n63543, n63544, n63545, n63546, n63547, n63548, n63549, n63550, n63551, n63552, n63553, n63554, n63555, n63556, n63557, n63558, n63559, n63560, n63561, n63562, n63563, n63564, n63565, n63566, n63567, n63568, n63569, n63570, n63571, n63572, n63573, n63574, n63575, n63576, n63577, n63578, n63579, n63580, n63581, n63582, n63583, n63584, n63585, n63586, n63587, n63588, n63589, n63590, n63591, n63592, n63593, n63594, n63595, n63596, n63597, n63598, n63599, n63600, n63601, n63602, n63603, n63604, n63605, n63606, n63607, n63608, n63609, n63610, n63611, n63612, n63613, n63614, n63615, n63616, n63617, n63618, n63619, n63620, n63621, n63622, n63623, n63624, n63625, n63626, n63627, n63628, n63629, n63630, n63631, n63632, n63633, n63634, n63635, n63636, n63637, n63638, n63639, n63640, n63641, n63642, n63643, n63644, n63645, n63646, n63647, n63648, n63649, n63650, n63651, n63652, n63653, n63654, n63655, n63656, n63657, n63658, n63659, n63660, n63661, n63662, n63663, n63664, n63665, n63666, n63667, n63668, n63669, n63670, n63671, n63672, n63673, n63674, n63675, n63676, n63677, n63678, n63679, n63680, n63681, n63682, n63683, n63684, n63685, n63686, n63687, n63688, n63689, n63690, n63691, n63692, n63693, n63694, n63695, n63696, n63697, n63698, n63699, n63700, n63701, n63702, n63703, n63704, n63705, n63706, n63707, n63708, n63709, n63710, n63711, n63712, n63713, n63714, n63715, n63716, n63717, n63718, n63719, n63720, n63721, n63722, n63723, n63724, n63725, n63726, n63727, n63728, n63729, n63730, n63731, n63732, n63733, n63734, n63735, n63736, n63737, n63738, n63739, n63740, n63741, n63742, n63743, n63744, n63745, n63746, n63747, n63748, n63749, n63750, n63751, n63752, n63753, n63754, n63755, n63756, n63757, n63758, n63759, n63760, n63761, n63762, n63763, n63764, n63765, n63766, n63767, n63768, n63769, n63770, n63771, n63772, n63773, n63774, n63775, n63776, n63777, n63778, n63779, n63780, n63781, n63782, n63783, n63784, n63785, n63786, n63787, n63788, n63789, n63790, n63791, n63792, n63793, n63794, n63795, n63796, n63797, n63798, n63799, n63800, n63801, n63802, n63803, n63804, n63805, n63806, n63807, n63808, n63809, n63810, n63811, n63812, n63813, n63814, n63815, n63816, n63817, n63818, n63819, n63820, n63821, n63822, n63823, n63824, n63825, n63826, n63827, n63828, n63829, n63830, n63831, n63832, n63833, n63834, n63835, n63836, n63837, n63838, n63839, n63840, n63841, n63842, n63843, n63844, n63845, n63846, n63847, n63848, n63849, n63850, n63851, n63852, n63853, n63854, n63855, n63856, n63857, n63858, n63859, n63860, n63861, n63862, n63863, n63864, n63865, n63866, n63867, n63868, n63869, n63870, n63871, n63872, n63873, n63874, n63875, n63876, n63877, n63878, n63879, n63880, n63881, n63882, n63883, n63884, n63885, n63886, n63887, n63888, n63889, n63890, n63891, n63892, n63893, n63894, n63895, n63896, n63897, n63898, n63899, n63900, n63901, n63902, n63903, n63904, n63905, n63906, n63907, n63908, n63909, n63910, n63911, n63912, n63913, n63914, n63915, n63916, n63917, n63918, n63919, n63920, n63921, n63922, n63923, n63924, n63925, n63926, n63927, n63928, n63929, n63930, n63931, n63932, n63933, n63934, n63935, n63936, n63937, n63938, n63939, n63940, n63941, n63942, n63943, n63944, n63945, n63946, n63947, n63948, n63949, n63950, n63951, n63952, n63953, n63954, n63955, n63956, n63957, n63958, n63959, n63960, n63961, n63962, n63963, n63964, n63965, n63966, n63967, n63968, n63969, n63970, n63971, n63972, n63973, n63974, n63975, n63976, n63977, n63978, n63979, n63980, n63981, n63982, n63983, n63984, n63985, n63986, n63987, n63988, n63989, n63990, n63991, n63992, n63993, n63994, n63995, n63996, n63997, n63998, n63999, n64000, n64001, n64002, n64003, n64004, n64005, n64006, n64007, n64008, n64009, n64010, n64011, n64012, n64013, n64014, n64015, n64016, n64017, n64018, n64019, n64020, n64021, n64022, n64023, n64024, n64025, n64026, n64027, n64028, n64029, n64030, n64031, n64032, n64033, n64034, n64035, n64036, n64037, n64038, n64039, n64040, n64041, n64042, n64043, n64044, n64045, n64046, n64047, n64048, n64049, n64050, n64051, n64052, n64053, n64054, n64055, n64056, n64057, n64058, n64059, n64060, n64061, n64062, n64063, n64064, n64065, n64066, n64067, n64068, n64069, n64070, n64071, n64072, n64073, n64074, n64075, n64076, n64077, n64078, n64079, n64080, n64081, n64082, n64083, n64084, n64085, n64086, n64087, n64088, n64089, n64090, n64091, n64092, n64093, n64094, n64095, n64096, n64097, n64098, n64099, n64100, n64101, n64102, n64103, n64104, n64105, n64106, n64107, n64108, n64109, n64110, n64111, n64112, n64113, n64114, n64115, n64116, n64117, n64118, n64119, n64120, n64121, n64122, n64123, n64124, n64125, n64126, n64127, n64128, n64129, n64130, n64131, n64132, n64133, n64134, n64135, n64136, n64137, n64138, n64139, n64140, n64141, n64142, n64143, n64144, n64145, n64146, n64147, n64148, n64149, n64150, n64151, n64152, n64153, n64154, n64155, n64156, n64157, n64158, n64159, n64160, n64161, n64162, n64163, n64164, n64165, n64166, n64167, n64168, n64169, n64170, n64171, n64172, n64173, n64174, n64175, n64176, n64177, n64178, n64179, n64180, n64181, n64182, n64183, n64184, n64185, n64186, n64187, n64188, n64189, n64190, n64191, n64192, n64193, n64194, n64195, n64196, n64197, n64198, n64199, n64200, n64201, n64202, n64203, n64204, n64205, n64206, n64207, n64208, n64209, n64210, n64211, n64212, n64213, n64214, n64215, n64216, n64217, n64218, n64219, n64220, n64221, n64222, n64223, n64224, n64225, n64226, n64227, n64228, n64229, n64230, n64231, n64232, n64233, n64234, n64235, n64236, n64237, n64238, n64239, n64240, n64241, n64242, n64243, n64244, n64245, n64246, n64247, n64248, n64249, n64250, n64251, n64252, n64253, n64254, n64255, n64256, n64257, n64258, n64259, n64260, n64261, n64262, n64263, n64264, n64265, n64266, n64267, n64268, n64269, n64270, n64271, n64272, n64273, n64274, n64275, n64276, n64277, n64278, n64279, n64280, n64281, n64282, n64283, n64284, n64285, n64286, n64287, n64288, n64289, n64290, n64291, n64292, n64293, n64294, n64295, n64296, n64297, n64298, n64299, n64300, n64301, n64302, n64303, n64304, n64305, n64306, n64307, n64308, n64309, n64310, n64311, n64312, n64313, n64314, n64315, n64316, n64317, n64318, n64319, n64320, n64321, n64322, n64323, n64324, n64325, n64326, n64327, n64328, n64329, n64330, n64331, n64332, n64333, n64334, n64335, n64336, n64337, n64338, n64339, n64340, n64341, n64342, n64343, n64344, n64345, n64346, n64347, n64348, n64349, n64350, n64351, n64352, n64353, n64354, n64355, n64356, n64357, n64358, n64359, n64360, n64361, n64362, n64363, n64364, n64365, n64366, n64367, n64368, n64369, n64370, n64371, n64372, n64373, n64374, n64375, n64376, n64377, n64378, n64379, n64380, n64381, n64382, n64383, n64384, n64385, n64386, n64387, n64388, n64389, n64390, n64391, n64392, n64393, n64394, n64395, n64396, n64397, n64398, n64399, n64400, n64401, n64402, n64403, n64404, n64405, n64406, n64407, n64408, n64409, n64410, n64411, n64412, n64413, n64414, n64415, n64416, n64417, n64418, n64419, n64420, n64421, n64422, n64423, n64424, n64425, n64426, n64427, n64428, n64429, n64430, n64431, n64432, n64433, n64434, n64435, n64436, n64437, n64438, n64439, n64440, n64441, n64442, n64443, n64444, n64445, n64446, n64447, n64448, n64449, n64450, n64451, n64452, n64453, n64454, n64455, n64456, n64457, n64458, n64459, n64460, n64461, n64462, n64463, n64464, n64465, n64466, n64467, n64468, n64469, n64470, n64471, n64472, n64473, n64474, n64475, n64476, n64477, n64478, n64479, n64480, n64481, n64482, n64483, n64484, n64485, n64486, n64487, n64488, n64489, n64490, n64491, n64492, n64493, n64494, n64495, n64496, n64497, n64498, n64499, n64500, n64501, n64502, n64503, n64504, n64505, n64506, n64507, n64508, n64509, n64510, n64511, n64512, n64513, n64514, n64515, n64516, n64517, n64518, n64519, n64520, n64521, n64522, n64523, n64524, n64525, n64526, n64527, n64528, n64529, n64530, n64531, n64532, n64533, n64534, n64535, n64536, n64537, n64538, n64539, n64540, n64541, n64542, n64543, n64544, n64545, n64546, n64547, n64548, n64549, n64550, n64551, n64552, n64553, n64554, n64555, n64556, n64557, n64558, n64559, n64560, n64561, n64562, n64563, n64564, n64565, n64566, n64567, n64568, n64569, n64570, n64571, n64572, n64573, n64574, n64575, n64576, n64577, n64578, n64579, n64580, n64581, n64582, n64583, n64584, n64585, n64586, n64587, n64588, n64589, n64590, n64591, n64592, n64593, n64594, n64595, n64596, n64597, n64598, n64599, n64600, n64601, n64602, n64603, n64604, n64605, n64606, n64607, n64608, n64609, n64610, n64611, n64612, n64613, n64614, n64615, n64616, n64617, n64618, n64619, n64620, n64621, n64622, n64623, n64624, n64625, n64626, n64627, n64628, n64629, n64630, n64631, n64632, n64633, n64634, n64635, n64636, n64637, n64638, n64639, n64640, n64641, n64642, n64643, n64644, n64645, n64646, n64647, n64648, n64649, n64650, n64651, n64652, n64653, n64654, n64655, n64656, n64657, n64658, n64659, n64660, n64661, n64662, n64663, n64664, n64665, n64666, n64667, n64668, n64669, n64670, n64671, n64672, n64673, n64674, n64675, n64676, n64677, n64678, n64679, n64680, n64681, n64682, n64683, n64684, n64685, n64686, n64687, n64688, n64689, n64690, n64691, n64692, n64693, n64694, n64695, n64696, n64697, n64698, n64699, n64700, n64701, n64702, n64703, n64704, n64705, n64706, n64707, n64708, n64709, n64710, n64711, n64712, n64713, n64714, n64715, n64716, n64717, n64718, n64719, n64720, n64721, n64722, n64723, n64724, n64725, n64726, n64727, n64728, n64729, n64730, n64731, n64732, n64733, n64734, n64735, n64736, n64737, n64738, n64739, n64740, n64741, n64742, n64743, n64744, n64745, n64746, n64747, n64748, n64749, n64750, n64751, n64752, n64753, n64754, n64755, n64756, n64757, n64758, n64759, n64760, n64761, n64762, n64763, n64764, n64765, n64766, n64767, n64768, n64769, n64770, n64771, n64772, n64773, n64774, n64775, n64776, n64777, n64778, n64779, n64780, n64781, n64782, n64783, n64784, n64785, n64786, n64787, n64788, n64789, n64790, n64791, n64792, n64793, n64794, n64795, n64796, n64797, n64798, n64799, n64800, n64801, n64802, n64803, n64804, n64805, n64806, n64807, n64808, n64809, n64810, n64811, n64812, n64813, n64814, n64815, n64816, n64817, n64818, n64819, n64820, n64821, n64822, n64823, n64824, n64825, n64826, n64827, n64828, n64829, n64830, n64831, n64832, n64833, n64834, n64835, n64836, n64837, n64838, n64839, n64840, n64841, n64842, n64843, n64844, n64845, n64846, n64847, n64848, n64849, n64850, n64851, n64852, n64853, n64854, n64855, n64856, n64857, n64858, n64859, n64860, n64861, n64862, n64863, n64864, n64865, n64866, n64867, n64868, n64869, n64870, n64871, n64872, n64873, n64874, n64875, n64876, n64877, n64878, n64879, n64880, n64881, n64882, n64883, n64884, n64885, n64886, n64887, n64888, n64889, n64890, n64891, n64892, n64893, n64894, n64895, n64896, n64897, n64898, n64899, n64900, n64901, n64902, n64903, n64904, n64905, n64906, n64907, n64908, n64909, n64910, n64911, n64912, n64913, n64914, n64915, n64916, n64917, n64918, n64919, n64920, n64921, n64922, n64923, n64924, n64925, n64926, n64927, n64928, n64929, n64930, n64931, n64932, n64933, n64934, n64935, n64936, n64937, n64938, n64939, n64940, n64941, n64942, n64943, n64944, n64945, n64946, n64947, n64948, n64949, n64950, n64951, n64952, n64953, n64954, n64955, n64956, n64957, n64958, n64959, n64960, n64961, n64962, n64963, n64964, n64965, n64966, n64967, n64968, n64969, n64970, n64971, n64972, n64973, n64974, n64975, n64976, n64977, n64978, n64979, n64980, n64981, n64982, n64983, n64984, n64985, n64986, n64987, n64988, n64989, n64990, n64991, n64992, n64993, n64994, n64995, n64996, n64997, n64998, n64999, n65000, n65001, n65002, n65003, n65004, n65005, n65006, n65007, n65008, n65009, n65010, n65011, n65012, n65013, n65014, n65015, n65016, n65017, n65018, n65019, n65020, n65021, n65022, n65023, n65024, n65025, n65026, n65027, n65028, n65029, n65030, n65031, n65032, n65033, n65034, n65035, n65036, n65037, n65038, n65039, n65040, n65041, n65042, n65043, n65044, n65045, n65046, n65047, n65048, n65049, n65050, n65051, n65052, n65053, n65054, n65055, n65056, n65057, n65058, n65059, n65060, n65061, n65062, n65063, n65064, n65065, n65066, n65067, n65068, n65069, n65070, n65071, n65072, n65073, n65074, n65075, n65076, n65077, n65078, n65079, n65080, n65081, n65082, n65083, n65084, n65085, n65086, n65087, n65088, n65089, n65090, n65091, n65092, n65093, n65094, n65095, n65096, n65097, n65098, n65099, n65100, n65101, n65102, n65103, n65104, n65105, n65106, n65107, n65108, n65109, n65110, n65111, n65112, n65113, n65114, n65115, n65116, n65117, n65118, n65119, n65120, n65121, n65122, n65123, n65124, n65125, n65126, n65127, n65128, n65129, n65130, n65131, n65132, n65133, n65134, n65135, n65136, n65137, n65138, n65139, n65140, n65141, n65142, n65143, n65144, n65145, n65146, n65147, n65148, n65149, n65150, n65151, n65152, n65153, n65154, n65155, n65156, n65157, n65158, n65159, n65160, n65161, n65162, n65163, n65164, n65165, n65166, n65167, n65168, n65169, n65170, n65171, n65172, n65173, n65174, n65175, n65176, n65177, n65178, n65179, n65180, n65181, n65182, n65183, n65184, n65185, n65186, n65187, n65188, n65189, n65190, n65191, n65192, n65193, n65194, n65195, n65196, n65197, n65198, n65199, n65200, n65201, n65202, n65203, n65204, n65205, n65206, n65207, n65208, n65209, n65210, n65211, n65212, n65213, n65214, n65215, n65216, n65217, n65218, n65219, n65220, n65221, n65222, n65223, n65224, n65225, n65226, n65227, n65228, n65229, n65230, n65231, n65232, n65233, n65234, n65235, n65236, n65237, n65238, n65239, n65240, n65241, n65242, n65243, n65244, n65245, n65246, n65247, n65248, n65249, n65250, n65251, n65252, n65253, n65254, n65255, n65256, n65257, n65258, n65259, n65260, n65261, n65262, n65263, n65264, n65265, n65266, n65267, n65268, n65269, n65270, n65271, n65272, n65273, n65274, n65275, n65276, n65277, n65278, n65279, n65280, n65281, n65282, n65283, n65284, n65285, n65286, n65287, n65288, n65289, n65290, n65291, n65292, n65293, n65294, n65295, n65296, n65297, n65298, n65299, n65300, n65301, n65302, n65303, n65304, n65305, n65306, n65307, n65308, n65309, n65310, n65311, n65312, n65313, n65314, n65315, n65316, n65317, n65318, n65319, n65320, n65321, n65322, n65323, n65324, n65325, n65326, n65327, n65328, n65329, n65330, n65331, n65332, n65333, n65334, n65335, n65336, n65337, n65338, n65339, n65340, n65341, n65342, n65343, n65344, n65345, n65346, n65347, n65348, n65349, n65350, n65351, n65352, n65353, n65354, n65355, n65356, n65357, n65358, n65359, n65360, n65361, n65362, n65363, n65364, n65365, n65366, n65367, n65368, n65369, n65370, n65371, n65372, n65373, n65374, n65375, n65376, n65377, n65378, n65379, n65380, n65381, n65382, n65383, n65384, n65385, n65386, n65387, n65388, n65389, n65390, n65391, n65392, n65393, n65394, n65395, n65396, n65397, n65398, n65399, n65400, n65401, n65402, n65403, n65404, n65405, n65406, n65407, n65408, n65409, n65410, n65411, n65412, n65413, n65414, n65415, n65416, n65417, n65418, n65419, n65420, n65421, n65422, n65423, n65424, n65425, n65426, n65427, n65428, n65429, n65430, n65431, n65432, n65433, n65434, n65435, n65436, n65437, n65438, n65439, n65440, n65441, n65442, n65443, n65444, n65445, n65446, n65447, n65448, n65449, n65450, n65451, n65452, n65453, n65454, n65455, n65456, n65457, n65458, n65459, n65460, n65461, n65462, n65463, n65464, n65465, n65466, n65467, n65468, n65469, n65470, n65471, n65472, n65473, n65474, n65475, n65476, n65477, n65478, n65479, n65480, n65481, n65482, n65483, n65484, n65485, n65486, n65487, n65488, n65489, n65490, n65491, n65492, n65493, n65494, n65495, n65496, n65497, n65498, n65499, n65500, n65501, n65502, n65503, n65504, n65505, n65506, n65507, n65508, n65509, n65510, n65511, n65512, n65513, n65514, n65515, n65516, n65517, n65518, n65519, n65520, n65521, n65522, n65523, n65524, n65525, n65526, n65527, n65528, n65529, n65530, n65531, n65532, n65533, n65534, n65535, n65536, n65537, n65538, n65539, n65540, n65541, n65542, n65543, n65544, n65545, n65546, n65547, n65548, n65549, n65550, n65551, n65552, n65553, n65554, n65555, n65556, n65557, n65558, n65559, n65560, n65561, n65562, n65563, n65564, n65565, n65566, n65567, n65568, n65569, n65570, n65571, n65572, n65573, n65574, n65575, n65576, n65577, n65578, n65579, n65580, n65581, n65582, n65583, n65584, n65585, n65586, n65587, n65588, n65589, n65590, n65591, n65592, n65593, n65594, n65595, n65596, n65597, n65598, n65599, n65600, n65601, n65602, n65603, n65604, n65605, n65606, n65607, n65608, n65609, n65610, n65611, n65612, n65613, n65614, n65615, n65616, n65617, n65618, n65619, n65620, n65621, n65622, n65623, n65624, n65625, n65626, n65627, n65628, n65629, n65630, n65631, n65632, n65633, n65634, n65635, n65636, n65637, n65638, n65639, n65640, n65641, n65642, n65643, n65644, n65645, n65646, n65647, n65648, n65649, n65650, n65651, n65652, n65653, n65654, n65655, n65656, n65657, n65658, n65659, n65660, n65661, n65662, n65663, n65664, n65665, n65666, n65667, n65668, n65669, n65670, n65671, n65672, n65673, n65674, n65675, n65676, n65677, n65678, n65679, n65680, n65681, n65682, n65683, n65684, n65685, n65686, n65687, n65688, n65689, n65690, n65691, n65692, n65693, n65694, n65695, n65696, n65697, n65698, n65699, n65700, n65701, n65702, n65703, n65704, n65705, n65706, n65707, n65708, n65709, n65710, n65711, n65712, n65713, n65714, n65715, n65716, n65717, n65718, n65719, n65720, n65721, n65722, n65723, n65724, n65725, n65726, n65727, n65728, n65729, n65730, n65731, n65732, n65733, n65734, n65735, n65736, n65737, n65738, n65739, n65740, n65741, n65742, n65743, n65744, n65745, n65746, n65747, n65748, n65749, n65750, n65751, n65752, n65753, n65754, n65755, n65756, n65757, n65758, n65759, n65760, n65761, n65762, n65763, n65764, n65765, n65766, n65767, n65768, n65769, n65770, n65771, n65772, n65773, n65774, n65775, n65776, n65777, n65778, n65779, n65780, n65781, n65782, n65783, n65784, n65785, n65786, n65787, n65788, n65789, n65790, n65791, n65792, n65793, n65794, n65795, n65796, n65797, n65798, n65799, n65800, n65801, n65802, n65803, n65804, n65805, n65806, n65807, n65808, n65809, n65810, n65811, n65812, n65813, n65814, n65815, n65816, n65817, n65818, n65819, n65820, n65821, n65822, n65823, n65824, n65825, n65826, n65827, n65828, n65829, n65830, n65831, n65832, n65833, n65834, n65835, n65836, n65837, n65838, n65839, n65840, n65841, n65842, n65843, n65844, n65845, n65846, n65847, n65848, n65849, n65850, n65851, n65852, n65853, n65854, n65855, n65856, n65857, n65858, n65859, n65860, n65861, n65862, n65863, n65864, n65865, n65866, n65867, n65868, n65869, n65870, n65871, n65872, n65873, n65874, n65875, n65876, n65877, n65878, n65879, n65880, n65881, n65882, n65883, n65884, n65885, n65886, n65887, n65888, n65889, n65890, n65891, n65892, n65893, n65894, n65895, n65896, n65897, n65898, n65899, n65900, n65901, n65902, n65903, n65904, n65905, n65906, n65907, n65908, n65909, n65910, n65911, n65912, n65913, n65914, n65915, n65916, n65917, n65918, n65919, n65920, n65921, n65922, n65923, n65924, n65925, n65926, n65927, n65928, n65929, n65930, n65931, n65932, n65933, n65934, n65935, n65936, n65937, n65938, n65939, n65940, n65941, n65942, n65943, n65944, n65945, n65946, n65947, n65948, n65949, n65950, n65951, n65952, n65953, n65954, n65955, n65956, n65957, n65958, n65959, n65960, n65961, n65962, n65963, n65964, n65965, n65966, n65967, n65968, n65969, n65970, n65971, n65972, n65973, n65974, n65975, n65976, n65977, n65978, n65979, n65980, n65981, n65982, n65983, n65984, n65985, n65986, n65987, n65988, n65989, n65990, n65991, n65992, n65993, n65994, n65995, n65996, n65997, n65998, n65999, n66000, n66001, n66002, n66003, n66004, n66005, n66006, n66007, n66008, n66009, n66010, n66011, n66012, n66013, n66014, n66015, n66016, n66017, n66018, n66019, n66020, n66021, n66022, n66023, n66024, n66025, n66026, n66027, n66028, n66029, n66030, n66031, n66032, n66033, n66034, n66035, n66036, n66037, n66038, n66039, n66040, n66041, n66042, n66043, n66044, n66045, n66046, n66047, n66048, n66049, n66050, n66051, n66052, n66053, n66054, n66055, n66056, n66057, n66058, n66059, n66060, n66061, n66062, n66063, n66064, n66065, n66066, n66067, n66068, n66069, n66070, n66071, n66072, n66073, n66074, n66075, n66076, n66077, n66078, n66079, n66080, n66081, n66082, n66083, n66084, n66085, n66086, n66087, n66088, n66089, n66090, n66091, n66092, n66093, n66094, n66095, n66096, n66097, n66098, n66099, n66100, n66101, n66102, n66103, n66104, n66105, n66106, n66107, n66108, n66109, n66110, n66111, n66112, n66113, n66114, n66115, n66116, n66117, n66118, n66119, n66120, n66121, n66122, n66123, n66124, n66125, n66126, n66127, n66128, n66129, n66130, n66131, n66132, n66133, n66134, n66135, n66136, n66137, n66138, n66139, n66140, n66141, n66142, n66143, n66144, n66145, n66146, n66147, n66148, n66149, n66150, n66151, n66152, n66153, n66154, n66155, n66156, n66157, n66158, n66159, n66160, n66161, n66162, n66163, n66164, n66165, n66166, n66167, n66168, n66169, n66170, n66171, n66172, n66173, n66174, n66175, n66176, n66177, n66178, n66179, n66180, n66181, n66182, n66183, n66184, n66185, n66186, n66187, n66188, n66189, n66190, n66191, n66192, n66193, n66194, n66195, n66196, n66197, n66198, n66199, n66200, n66201, n66202, n66203, n66204, n66205, n66206, n66207, n66208, n66209, n66210, n66211, n66212, n66213, n66214, n66215, n66216, n66217, n66218, n66219, n66220, n66221, n66222, n66223, n66224, n66225, n66226, n66227, n66228, n66229, n66230, n66231, n66232, n66233, n66234, n66235, n66236, n66237, n66238, n66239, n66240, n66241, n66242, n66243, n66244, n66245, n66246, n66247, n66248, n66249, n66250, n66251, n66252, n66253, n66254, n66255, n66256, n66257, n66258, n66259, n66260, n66261, n66262, n66263, n66264, n66265, n66266, n66267, n66268, n66269, n66270, n66271, n66272, n66273, n66274, n66275, n66276, n66277, n66278, n66279, n66280, n66281, n66282, n66283, n66284, n66285, n66286, n66287, n66288, n66289, n66290, n66291, n66292, n66293, n66294, n66295, n66296, n66297, n66298, n66299, n66300, n66301, n66302, n66303, n66304, n66305, n66306, n66307, n66308, n66309, n66310, n66311, n66312, n66313, n66314, n66315, n66316, n66317, n66318, n66319, n66320, n66321, n66322, n66323, n66324, n66325, n66326, n66327, n66328, n66329, n66330, n66331, n66332, n66333, n66334, n66335, n66336, n66337, n66338, n66339, n66340, n66341, n66342, n66343, n66344, n66345, n66346, n66347, n66348, n66349, n66350, n66351, n66352, n66353, n66354, n66355, n66356, n66357, n66358, n66359, n66360, n66361, n66362, n66363, n66364, n66365, n66366, n66367, n66368, n66369, n66370, n66371, n66372, n66373, n66374, n66375, n66376, n66377, n66378, n66379, n66380, n66381, n66382, n66383, n66384, n66385, n66386, n66387, n66388, n66389, n66390, n66391, n66392, n66393, n66394, n66395, n66396, n66397, n66398, n66399, n66400, n66401, n66402, n66403, n66404, n66405, n66406, n66407, n66408, n66409, n66410, n66411, n66412, n66413, n66414, n66415, n66416, n66417, n66418, n66419, n66420, n66421, n66422, n66423, n66424, n66425, n66426, n66427, n66428, n66429, n66430, n66431, n66432, n66433, n66434, n66435, n66436, n66437, n66438, n66439, n66440, n66441, n66442, n66443, n66444, n66445, n66446, n66447, n66448, n66449, n66450, n66451, n66452, n66453, n66454, n66455, n66456, n66457, n66458, n66459, n66460, n66461, n66462, n66463, n66464, n66465, n66466, n66467, n66468, n66469, n66470, n66471, n66472, n66473, n66474, n66475, n66476, n66477, n66478, n66479, n66480, n66481, n66482, n66483, n66484, n66485, n66486, n66487, n66488, n66489, n66490, n66491, n66492, n66493, n66494, n66495, n66496, n66497, n66498, n66499, n66500, n66501, n66502, n66503, n66504, n66505, n66506, n66507, n66508, n66509, n66510, n66511, n66512, n66513, n66514, n66515, n66516, n66517, n66518, n66519, n66520, n66521, n66522, n66523, n66524, n66525, n66526, n66527, n66528, n66529, n66530, n66531, n66532, n66533, n66534, n66535, n66536, n66537, n66538, n66539, n66540, n66541, n66542, n66543, n66544, n66545, n66546, n66547, n66548, n66549, n66550, n66551, n66552, n66553, n66554, n66555, n66556, n66557, n66558, n66559, n66560, n66561, n66562, n66563, n66564, n66565, n66566, n66567, n66568, n66569, n66570, n66571, n66572, n66573, n66574, n66575, n66576, n66577, n66578, n66579, n66580, n66581, n66582, n66583, n66584, n66585, n66586, n66587, n66588, n66589, n66590, n66591, n66592, n66593, n66594, n66595, n66596, n66597, n66598, n66599, n66600, n66601, n66602, n66603, n66604, n66605, n66606, n66607, n66608, n66609, n66610, n66611, n66612, n66613, n66614, n66615, n66616, n66617, n66618, n66619, n66620, n66621, n66622, n66623, n66624, n66625, n66626, n66627, n66628, n66629, n66630, n66631, n66632, n66633, n66634, n66635, n66636, n66637, n66638, n66639, n66640, n66641, n66642, n66643, n66644, n66645, n66646, n66647, n66648, n66649, n66650, n66651, n66652, n66653, n66654, n66655, n66656, n66657, n66658, n66659, n66660, n66661, n66662, n66663, n66664, n66665, n66666, n66667, n66668, n66669, n66670, n66671, n66672, n66673, n66674, n66675, n66676, n66677, n66678, n66679, n66680, n66681, n66682, n66683, n66684, n66685, n66686, n66687, n66688, n66689, n66690, n66691, n66692, n66693, n66694, n66695, n66696, n66697, n66698, n66699, n66700, n66701, n66702, n66703, n66704, n66705, n66706, n66707, n66708, n66709, n66710, n66711, n66712, n66713, n66714, n66715, n66716, n66717, n66718, n66719, n66720, n66721, n66722, n66723, n66724, n66725, n66726, n66727, n66728, n66729, n66730, n66731, n66732, n66733, n66734, n66735, n66736, n66737, n66738, n66739, n66740, n66741, n66742, n66743, n66744, n66745, n66746, n66747, n66748, n66749, n66750, n66751, n66752, n66753, n66754, n66755, n66756, n66757, n66758, n66759, n66760, n66761, n66762, n66763, n66764, n66765, n66766, n66767, n66768, n66769, n66770, n66771, n66772, n66773, n66774, n66775, n66776, n66777, n66778, n66779, n66780, n66781, n66782, n66783, n66784, n66785, n66786, n66787, n66788, n66789, n66790, n66791, n66792, n66793, n66794, n66795, n66796, n66797, n66798, n66799, n66800, n66801, n66802, n66803, n66804, n66805, n66806, n66807, n66808, n66809, n66810, n66811, n66812, n66813, n66814, n66815, n66816, n66817, n66818, n66819, n66820, n66821, n66822, n66823, n66824, n66825, n66826, n66827, n66828, n66829, n66830, n66831, n66832, n66833, n66834, n66835, n66836, n66837, n66838, n66839, n66840, n66841, n66842, n66843, n66844, n66845, n66846, n66847, n66848, n66849, n66850, n66851, n66852, n66853, n66854, n66855, n66856, n66857, n66858, n66859, n66860, n66861, n66862, n66863, n66864, n66865, n66866, n66867, n66868, n66869, n66870, n66871, n66872, n66873, n66874, n66875, n66876, n66877, n66878, n66879, n66880, n66881, n66882, n66883, n66884, n66885, n66886, n66887, n66888, n66889, n66890, n66891, n66892, n66893, n66894, n66895, n66896, n66897, n66898, n66899, n66900, n66901, n66902, n66903, n66904, n66905, n66906, n66907, n66908, n66909, n66910, n66911, n66912, n66913, n66914, n66915, n66916, n66917, n66918, n66919, n66920, n66921, n66922, n66923, n66924, n66925, n66926, n66927, n66928, n66929, n66930, n66931, n66932, n66933, n66934, n66935, n66936, n66937, n66938, n66939, n66940, n66941, n66942, n66943, n66944, n66945, n66946, n66947, n66948, n66949, n66950, n66951, n66952, n66953, n66954, n66955, n66956, n66957, n66958, n66959, n66960, n66961, n66962, n66963, n66964, n66965, n66966, n66967, n66968, n66969, n66970, n66971, n66972, n66973, n66974, n66975, n66976, n66977, n66978, n66979, n66980, n66981, n66982, n66983, n66984, n66985, n66986, n66987, n66988, n66989, n66990, n66991, n66992, n66993, n66994, n66995, n66996, n66997, n66998, n66999, n67000, n67001, n67002, n67003, n67004, n67005, n67006, n67007, n67008, n67009, n67010, n67011, n67012, n67013, n67014, n67015, n67016, n67017, n67018, n67019, n67020, n67021, n67022, n67023, n67024, n67025, n67026, n67027, n67028, n67029, n67030, n67031, n67032, n67033, n67034, n67035, n67036, n67037, n67038, n67039, n67040, n67041, n67042, n67043, n67044, n67045, n67046, n67047, n67048, n67049, n67050, n67051, n67052, n67053, n67054, n67055, n67056, n67057, n67058, n67059, n67060, n67061, n67062, n67063, n67064, n67065, n67066, n67067, n67068, n67069, n67070, n67071, n67072, n67073, n67074, n67075, n67076, n67077, n67078, n67079, n67080, n67081, n67082, n67083, n67084, n67085, n67086, n67087, n67088, n67089, n67090, n67091, n67092, n67093, n67094, n67095, n67096, n67097, n67098, n67099, n67100, n67101, n67102, n67103, n67104, n67105, n67106, n67107, n67108, n67109, n67110, n67111, n67112, n67113, n67114, n67115, n67116, n67117, n67118, n67119, n67120, n67121, n67122, n67123, n67124, n67125, n67126, n67127, n67128, n67129, n67130, n67131, n67132, n67133, n67134, n67135, n67136, n67137, n67138, n67139, n67140, n67141, n67142, n67143, n67144, n67145, n67146, n67147, n67148, n67149, n67150, n67151, n67152, n67153, n67154, n67155, n67156, n67157, n67158, n67159, n67160, n67161, n67162, n67163, n67164, n67165, n67166, n67167, n67168, n67169, n67170, n67171, n67172, n67173, n67174, n67175, n67176, n67177, n67178, n67179, n67180, n67181, n67182, n67183, n67184, n67185, n67186, n67187, n67188, n67189, n67190, n67191, n67192, n67193, n67194, n67195, n67196, n67197, n67198, n67199, n67200, n67201, n67202, n67203, n67204, n67205, n67206, n67207, n67208, n67209, n67210, n67211, n67212, n67213, n67214, n67215, n67216, n67217, n67218, n67219, n67220, n67221, n67222, n67223, n67224, n67225, n67226, n67227, n67228, n67229, n67230, n67231, n67232, n67233, n67234, n67235, n67236, n67237, n67238, n67239, n67240, n67241, n67242, n67243, n67244, n67245, n67246, n67247, n67248, n67249, n67250, n67251, n67252, n67253, n67254, n67255, n67256, n67257, n67258, n67259, n67260, n67261, n67262, n67263, n67264, n67265, n67266, n67267, n67268, n67269, n67270, n67271, n67272, n67273, n67274, n67275, n67276, n67277, n67278, n67279, n67280, n67281, n67282, n67283, n67284, n67285, n67286, n67287, n67288, n67289, n67290, n67291, n67292, n67293, n67294, n67295, n67296, n67297, n67298, n67299, n67300, n67301, n67302, n67303, n67304, n67305, n67306, n67307, n67308, n67309, n67310, n67311, n67312, n67313, n67314, n67315, n67316, n67317, n67318, n67319, n67320, n67321, n67322, n67323, n67324, n67325, n67326, n67327, n67328, n67329, n67330, n67331, n67332, n67333, n67334, n67335, n67336, n67337, n67338, n67339, n67340, n67341, n67342, n67343, n67344, n67345, n67346, n67347, n67348, n67349, n67350, n67351, n67352, n67353, n67354, n67355, n67356, n67357, n67358, n67359, n67360, n67361, n67362, n67363, n67364, n67365, n67366, n67367, n67368, n67369, n67370, n67371, n67372, n67373, n67374, n67375, n67376, n67377, n67378, n67379, n67380, n67381, n67382, n67383, n67384, n67385, n67386, n67387, n67388, n67389, n67390, n67391, n67392, n67393, n67394, n67395, n67396, n67397, n67398, n67399, n67400, n67401, n67402, n67403, n67404, n67405, n67406, n67407, n67408, n67409, n67410, n67411, n67412, n67413, n67414, n67415, n67416, n67417, n67418, n67419, n67420, n67421, n67422, n67423, n67424, n67425, n67426, n67427, n67428, n67429, n67430, n67431, n67432, n67433, n67434, n67435, n67436, n67437, n67438, n67439, n67440, n67441, n67442, n67443, n67444, n67445, n67446, n67447, n67448, n67449, n67450, n67451, n67452, n67453, n67454, n67455, n67456, n67457, n67458, n67459, n67460, n67461, n67462, n67463, n67464, n67465, n67466, n67467, n67468, n67469, n67470, n67471, n67472, n67473, n67474, n67475, n67476, n67477, n67478, n67479, n67480, n67481, n67482, n67483, n67484, n67485, n67486, n67487, n67488, n67489, n67490, n67491, n67492, n67493, n67494, n67495, n67496, n67497, n67498, n67499, n67500, n67501, n67502, n67503, n67504, n67505, n67506, n67507, n67508, n67509, n67510, n67511, n67512, n67513, n67514, n67515, n67516, n67517, n67518, n67519, n67520, n67521, n67522, n67523, n67524, n67525, n67526, n67527, n67528, n67529, n67530, n67531, n67532, n67533, n67534, n67535, n67536, n67537, n67538, n67539, n67540, n67541, n67542, n67543, n67544, n67545, n67546, n67547, n67548, n67549, n67550, n67551, n67552, n67553, n67554, n67555, n67556, n67557, n67558, n67559, n67560, n67561, n67562, n67563, n67564, n67565, n67566, n67567, n67568, n67569, n67570, n67571, n67572, n67573, n67574, n67575, n67576, n67577, n67578, n67579, n67580, n67581, n67582, n67583, n67584, n67585, n67586, n67587, n67588, n67589, n67590, n67591, n67592, n67593, n67594, n67595, n67596, n67597, n67598, n67599, n67600, n67601, n67602, n67603, n67604, n67605, n67606, n67607, n67608, n67609, n67610, n67611, n67612, n67613, n67614, n67615, n67616, n67617, n67618, n67619, n67620, n67621, n67622, n67623, n67624, n67625, n67626, n67627, n67628, n67629, n67630, n67631, n67632, n67633, n67634, n67635, n67636, n67637, n67638, n67639, n67640, n67641, n67642, n67643, n67644, n67645, n67646, n67647, n67648, n67649, n67650, n67651, n67652, n67653, n67654, n67655, n67656, n67657, n67658, n67659, n67660, n67661, n67662, n67663, n67664, n67665, n67666, n67667, n67668, n67669, n67670, n67671, n67672, n67673, n67674, n67675, n67676, n67677, n67678, n67679, n67680, n67681, n67682, n67683, n67684, n67685, n67686, n67687, n67688, n67689, n67690, n67691, n67692, n67693, n67694, n67695, n67696, n67697, n67698, n67699, n67700, n67701, n67702, n67703, n67704, n67705, n67706, n67707, n67708, n67709, n67710, n67711, n67712, n67713, n67714, n67715, n67716, n67717, n67718, n67719, n67720, n67721, n67722, n67723, n67724, n67725, n67726, n67727, n67728, n67729, n67730, n67731, n67732, n67733, n67734, n67735, n67736, n67737, n67738, n67739, n67740, n67741, n67742, n67743, n67744, n67745, n67746, n67747, n67748, n67749, n67750, n67751, n67752, n67753, n67754, n67755, n67756, n67757, n67758, n67759, n67760, n67761, n67762, n67763, n67764, n67765, n67766, n67767, n67768, n67769, n67770, n67771, n67772, n67773, n67774, n67775, n67776, n67777, n67778, n67779, n67780, n67781, n67782, n67783, n67784, n67785, n67786, n67787, n67788, n67789, n67790, n67791, n67792, n67793, n67794, n67795, n67796, n67797, n67798, n67799, n67800, n67801, n67802, n67803, n67804, n67805, n67806, n67807, n67808, n67809, n67810, n67811, n67812, n67813, n67814, n67815, n67816, n67817, n67818, n67819, n67820, n67821, n67822, n67823, n67824, n67825, n67826, n67827, n67828, n67829, n67830, n67831, n67832, n67833, n67834, n67835, n67836, n67837, n67838, n67839, n67840, n67841, n67842, n67843, n67844, n67845, n67846, n67847, n67848, n67849, n67850, n67851, n67852, n67853, n67854, n67855, n67856, n67857, n67858, n67859, n67860, n67861, n67862, n67863, n67864, n67865, n67866, n67867, n67868, n67869, n67870, n67871, n67872, n67873, n67874, n67875, n67876, n67877, n67878, n67879, n67880, n67881, n67882, n67883, n67884, n67885, n67886, n67887, n67888, n67889, n67890, n67891, n67892, n67893, n67894, n67895, n67896, n67897, n67898, n67899, n67900, n67901, n67902, n67903, n67904, n67905, n67906, n67907, n67908, n67909, n67910, n67911, n67912, n67913, n67914, n67915, n67916, n67917, n67918, n67919, n67920, n67921, n67922, n67923, n67924, n67925, n67926, n67927, n67928, n67929, n67930, n67931, n67932, n67933, n67934, n67935, n67936, n67937, n67938, n67939, n67940, n67941, n67942, n67943, n67944, n67945, n67946, n67947, n67948, n67949, n67950, n67951, n67952, n67953, n67954, n67955, n67956, n67957, n67958, n67959, n67960, n67961, n67962, n67963, n67964, n67965, n67966, n67967, n67968, n67969, n67970, n67971, n67972, n67973, n67974, n67975, n67976, n67977, n67978, n67979, n67980, n67981, n67982, n67983, n67984, n67985, n67986, n67987, n67988, n67989, n67990, n67991, n67992, n67993, n67994, n67995, n67996, n67997, n67998, n67999, n68000, n68001, n68002, n68003, n68004, n68005, n68006, n68007, n68008, n68009, n68010, n68011, n68012, n68013, n68014, n68015, n68016, n68017, n68018, n68019, n68020, n68021, n68022, n68023, n68024, n68025, n68026, n68027, n68028, n68029, n68030, n68031, n68032, n68033, n68034, n68035, n68036, n68037, n68038, n68039, n68040, n68041, n68042, n68043, n68044, n68045, n68046, n68047, n68048, n68049, n68050, n68051, n68052, n68053, n68054, n68055, n68056, n68057, n68058, n68059, n68060, n68061, n68062, n68063, n68064, n68065, n68066, n68067, n68068, n68069, n68070, n68071, n68072, n68073, n68074, n68075, n68076, n68077, n68078, n68079, n68080, n68081, n68082, n68083, n68084, n68085, n68086, n68087, n68088, n68089, n68090, n68091, n68092, n68093, n68094, n68095, n68096, n68097, n68098, n68099, n68100, n68101, n68102, n68103, n68104, n68105, n68106, n68107, n68108, n68109, n68110, n68111, n68112, n68113, n68114, n68115, n68116, n68117, n68118, n68119, n68120, n68121, n68122, n68123, n68124, n68125, n68126, n68127, n68128, n68129, n68130, n68131, n68132, n68133, n68134, n68135, n68136, n68137, n68138, n68139, n68140, n68141, n68142, n68143, n68144, n68145, n68146, n68147, n68148, n68149, n68150, n68151, n68152, n68153, n68154, n68155, n68156, n68157, n68158, n68159, n68160, n68161, n68162, n68163, n68164, n68165, n68166, n68167, n68168, n68169, n68170, n68171, n68172, n68173, n68174, n68175, n68176, n68177, n68178, n68179, n68180, n68181, n68182, n68183, n68184, n68185, n68186, n68187, n68188, n68189, n68190, n68191, n68192, n68193, n68194, n68195, n68196, n68197, n68198, n68199, n68200, n68201, n68202, n68203, n68204, n68205, n68206, n68207, n68208, n68209, n68210, n68211, n68212, n68213, n68214, n68215, n68216, n68217, n68218, n68219, n68220, n68221, n68222, n68223, n68224, n68225, n68226, n68227, n68228, n68229, n68230, n68231, n68232, n68233, n68234, n68235, n68236, n68237, n68238, n68239, n68240, n68241, n68242, n68243, n68244, n68245, n68246, n68247, n68248, n68249, n68250, n68251, n68252, n68253, n68254, n68255, n68256, n68257, n68258, n68259, n68260, n68261, n68262, n68263, n68264, n68265, n68266, n68267, n68268, n68269, n68270, n68271, n68272, n68273, n68274, n68275, n68276, n68277, n68278, n68279, n68280, n68281, n68282, n68283, n68284, n68285, n68286, n68287, n68288, n68289, n68290, n68291, n68292, n68293, n68294, n68295, n68296, n68297, n68298, n68299, n68300, n68301, n68302, n68303, n68304, n68305, n68306, n68307, n68308, n68309, n68310, n68311, n68312, n68313, n68314, n68315, n68316, n68317, n68318, n68319, n68320, n68321, n68322, n68323, n68324, n68325, n68326, n68327, n68328, n68329, n68330, n68331, n68332, n68333, n68334, n68335, n68336, n68337, n68338, n68339, n68340, n68341, n68342, n68343, n68344, n68345, n68346, n68347, n68348, n68349, n68350, n68351, n68352, n68353, n68354, n68355, n68356, n68357, n68358, n68359, n68360, n68361, n68362, n68363, n68364, n68365, n68366, n68367, n68368, n68369, n68370, n68371, n68372, n68373, n68374, n68375, n68376, n68377, n68378, n68379, n68380, n68381, n68382, n68383, n68384, n68385, n68386, n68387, n68388, n68389, n68390, n68391, n68392, n68393, n68394, n68395, n68396, n68397, n68398, n68399, n68400, n68401, n68402, n68403, n68404, n68405, n68406, n68407, n68408, n68409, n68410, n68411, n68412, n68413, n68414, n68415, n68416, n68417, n68418, n68419, n68420, n68421, n68422, n68423, n68424, n68425, n68426, n68427, n68428, n68429, n68430, n68431, n68432, n68433, n68434, n68435, n68436, n68437, n68438, n68439, n68440, n68441, n68442, n68443, n68444, n68445, n68446, n68447, n68448, n68449, n68450, n68451, n68452, n68453, n68454, n68455, n68456, n68457, n68458, n68459, n68460, n68461, n68462, n68463, n68464, n68465, n68466, n68467, n68468, n68469, n68470, n68471, n68472, n68473, n68474, n68475, n68476, n68477, n68478, n68479, n68480, n68481, n68482, n68483, n68484, n68485, n68486, n68487, n68488, n68489, n68490, n68491, n68492, n68493, n68494, n68495, n68496, n68497, n68498, n68499, n68500, n68501, n68502, n68503, n68504, n68505, n68506, n68507, n68508, n68509, n68510, n68511, n68512, n68513, n68514, n68515, n68516, n68517, n68518, n68519, n68520, n68521, n68522, n68523, n68524, n68525, n68526, n68527, n68528, n68529, n68530, n68531, n68532, n68533, n68534, n68535, n68536, n68537, n68538, n68539, n68540, n68541, n68542, n68543, n68544, n68545, n68546, n68547, n68548, n68549, n68550, n68551, n68552, n68553, n68554, n68555, n68556, n68557, n68558, n68559, n68560, n68561, n68562, n68563, n68564, n68565, n68566, n68567, n68568, n68569, n68570, n68571, n68572, n68573, n68574, n68575, n68576, n68577, n68578, n68579, n68580, n68581, n68582, n68583, n68584, n68585, n68586, n68587, n68588, n68589, n68590, n68591, n68592, n68593, n68594, n68595, n68596, n68597, n68598, n68599, n68600, n68601, n68602, n68603, n68604, n68605, n68606, n68607, n68608, n68609, n68610, n68611, n68612, n68613, n68614, n68615, n68616, n68617, n68618, n68619, n68620, n68621, n68622, n68623, n68624, n68625, n68626, n68627, n68628, n68629, n68630, n68631, n68632, n68633, n68634, n68635, n68636, n68637, n68638, n68639, n68640, n68641, n68642, n68643, n68644, n68645, n68646, n68647, n68648, n68649, n68650, n68651, n68652, n68653, n68654, n68655, n68656, n68657, n68658, n68659, n68660, n68661, n68662, n68663, n68664, n68665, n68666, n68667, n68668, n68669, n68670, n68671, n68672, n68673, n68674, n68675, n68676, n68677, n68678, n68679, n68680, n68681, n68682, n68683, n68684, n68685, n68686, n68687, n68688, n68689, n68690, n68691, n68692, n68693, n68694, n68695, n68696, n68697, n68698, n68699, n68700, n68701, n68702, n68703, n68704, n68705, n68706, n68707, n68708, n68709, n68710, n68711, n68712, n68713, n68714, n68715, n68716, n68717, n68718, n68719, n68720, n68721, n68722, n68723, n68724, n68725, n68726, n68727, n68728, n68729, n68730, n68731, n68732, n68733, n68734, n68735, n68736, n68737, n68738, n68739, n68740, n68741, n68742, n68743, n68744, n68745, n68746, n68747, n68748, n68749, n68750, n68751, n68752, n68753, n68754, n68755, n68756, n68757, n68758, n68759, n68760, n68761, n68762, n68763, n68764, n68765, n68766, n68767, n68768, n68769, n68770, n68771, n68772, n68773, n68774, n68775, n68776, n68777, n68778, n68779, n68780, n68781, n68782, n68783, n68784, n68785, n68786, n68787, n68788, n68789, n68790, n68791, n68792, n68793, n68794, n68795, n68796, n68797, n68798, n68799, n68800, n68801, n68802, n68803, n68804, n68805, n68806, n68807, n68808, n68809, n68810, n68811, n68812, n68813, n68814, n68815, n68816, n68817, n68818, n68819, n68820, n68821, n68822, n68823, n68824, n68825, n68826, n68827, n68828, n68829, n68830, n68831, n68832, n68833, n68834, n68835, n68836, n68837, n68838, n68839, n68840, n68841, n68842, n68843, n68844, n68845, n68846, n68847, n68848, n68849, n68850, n68851, n68852, n68853, n68854, n68855, n68856, n68857, n68858, n68859, n68860, n68861, n68862, n68863, n68864, n68865, n68866, n68867, n68868, n68869, n68870, n68871, n68872, n68873, n68874, n68875, n68876, n68877, n68878, n68879, n68880, n68881, n68882, n68883, n68884, n68885, n68886, n68887, n68888, n68889, n68890, n68891, n68892, n68893, n68894, n68895, n68896, n68897, n68898, n68899, n68900, n68901, n68902, n68903, n68904, n68905, n68906, n68907, n68908, n68909, n68910, n68911, n68912, n68913, n68914, n68915, n68916, n68917, n68918, n68919, n68920, n68921, n68922, n68923, n68924, n68925, n68926, n68927, n68928, n68929, n68930, n68931, n68932, n68933, n68934, n68935, n68936, n68937, n68938, n68939, n68940, n68941, n68942, n68943, n68944, n68945, n68946, n68947, n68948, n68949, n68950, n68951, n68952, n68953, n68954, n68955, n68956, n68957, n68958, n68959, n68960, n68961, n68962, n68963, n68964, n68965, n68966, n68967, n68968, n68969, n68970, n68971, n68972, n68973, n68974, n68975, n68976, n68977, n68978, n68979, n68980, n68981, n68982, n68983, n68984, n68985, n68986, n68987, n68988, n68989, n68990, n68991, n68992, n68993, n68994, n68995, n68996, n68997, n68998, n68999, n69000, n69001, n69002, n69003, n69004, n69005, n69006, n69007, n69008, n69009, n69010, n69011, n69012, n69013, n69014, n69015, n69016, n69017, n69018, n69019, n69020, n69021, n69022, n69023, n69024, n69025, n69026, n69027, n69028, n69029, n69030, n69031, n69032, n69033, n69034, n69035, n69036, n69037, n69038, n69039, n69040, n69041, n69042, n69043, n69044, n69045, n69046, n69047, n69048, n69049, n69050, n69051, n69052, n69053, n69054, n69055, n69056, n69057, n69058, n69059, n69060, n69061, n69062, n69063, n69064, n69065, n69066, n69067, n69068, n69069, n69070, n69071, n69072, n69073, n69074, n69075, n69076, n69077, n69078, n69079, n69080, n69081, n69082, n69083, n69084, n69085, n69086, n69087, n69088, n69089, n69090, n69091, n69092, n69093, n69094, n69095, n69096, n69097, n69098, n69099, n69100, n69101, n69102, n69103, n69104, n69105, n69106, n69107, n69108, n69109, n69110, n69111, n69112, n69113, n69114, n69115, n69116, n69117, n69118, n69119, n69120, n69121, n69122, n69123, n69124, n69125, n69126, n69127, n69128, n69129, n69130, n69131, n69132, n69133, n69134, n69135, n69136, n69137, n69138, n69139, n69140, n69141, n69142, n69143, n69144, n69145, n69146, n69147, n69148, n69149, n69150, n69151, n69152, n69153, n69154, n69155, n69156, n69157, n69158, n69159, n69160, n69161, n69162, n69163, n69164, n69165, n69166, n69167, n69168, n69169, n69170, n69171, n69172, n69173, n69174, n69175, n69176, n69177, n69178, n69179, n69180, n69181, n69182, n69183, n69184, n69185, n69186, n69187, n69188, n69189, n69190, n69191, n69192, n69193, n69194, n69195, n69196, n69197, n69198, n69199, n69200, n69201, n69202, n69203, n69204, n69205, n69206, n69207, n69208, n69209, n69210, n69211, n69212, n69213, n69214, n69215, n69216, n69217, n69218, n69219, n69220, n69221, n69222, n69223, n69224, n69225, n69226, n69227, n69228, n69229, n69230, n69231, n69232, n69233, n69234, n69235, n69236, n69237, n69238, n69239, n69240, n69241, n69242, n69243, n69244, n69245, n69246, n69247, n69248, n69249, n69250, n69251, n69252, n69253, n69254, n69255, n69256, n69257, n69258, n69259, n69260, n69261, n69262, n69263, n69264, n69265, n69266, n69267, n69268, n69269, n69270, n69271, n69272, n69273, n69274, n69275, n69276, n69277, n69278, n69279, n69280, n69281, n69282, n69283, n69284, n69285, n69286, n69287, n69288, n69289, n69290, n69291, n69292, n69293, n69294, n69295, n69296, n69297, n69298, n69299, n69300, n69301, n69302, n69303, n69304, n69305, n69306, n69307, n69308, n69309, n69310, n69311, n69312, n69313, n69314, n69315, n69316, n69317, n69318, n69319, n69320, n69321, n69322, n69323, n69324, n69325, n69326, n69327, n69328, n69329, n69330, n69331, n69332, n69333, n69334, n69335, n69336, n69337, n69338, n69339, n69340, n69341, n69342, n69343, n69344, n69345, n69346, n69347, n69348, n69349, n69350, n69351, n69352, n69353, n69354, n69355, n69356, n69357, n69358, n69359, n69360, n69361, n69362, n69363, n69364, n69365, n69366, n69367, n69368, n69369, n69370, n69371, n69372, n69373, n69374, n69375, n69376, n69377, n69378, n69379, n69380, n69381, n69382, n69383, n69384, n69385, n69386, n69387, n69388, n69389, n69390, n69391, n69392, n69393, n69394, n69395, n69396, n69397, n69398, n69399, n69400, n69401, n69402, n69403, n69404, n69405, n69406, n69407, n69408, n69409, n69410, n69411, n69412, n69413, n69414, n69415, n69416, n69417, n69418, n69419, n69420, n69421, n69422, n69423, n69424, n69425, n69426, n69427, n69428, n69429, n69430, n69431, n69432, n69433, n69434, n69435, n69436, n69437, n69438, n69439, n69440, n69441, n69442, n69443, n69444, n69445, n69446, n69447, n69448, n69449, n69450, n69451, n69452, n69453, n69454, n69455, n69456, n69457, n69458, n69459, n69460, n69461, n69462, n69463, n69464, n69465, n69466, n69467, n69468, n69469, n69470, n69471, n69472, n69473, n69474, n69475, n69476, n69477, n69478, n69479, n69480, n69481, n69482, n69483, n69484, n69485, n69486, n69487, n69488, n69489, n69490, n69491, n69492, n69493, n69494, n69495, n69496, n69497, n69498, n69499, n69500, n69501, n69502, n69503, n69504, n69505, n69506, n69507, n69508, n69509, n69510, n69511, n69512, n69513, n69514, n69515, n69516, n69517, n69518, n69519, n69520, n69521, n69522, n69523, n69524, n69525, n69526, n69527, n69528, n69529, n69530, n69531, n69532, n69533, n69534, n69535, n69536, n69537, n69538, n69539, n69540, n69541, n69542, n69543, n69544, n69545, n69546, n69547, n69548, n69549, n69550, n69551, n69552, n69553, n69554, n69555, n69556, n69557, n69558, n69559, n69560, n69561, n69562, n69563, n69564, n69565, n69566, n69567, n69568, n69569, n69570, n69571, n69572, n69573, n69574, n69575, n69576, n69577, n69578, n69579, n69580, n69581, n69582, n69583, n69584, n69585, n69586, n69587, n69588, n69589, n69590, n69591, n69592, n69593, n69594, n69595, n69596, n69597, n69598, n69599, n69600, n69601, n69602, n69603, n69604, n69605, n69606, n69607, n69608, n69609, n69610, n69611, n69612, n69613, n69614, n69615, n69616, n69617, n69618, n69619, n69620, n69621, n69622, n69623, n69624, n69625, n69626, n69627, n69628, n69629, n69630, n69631, n69632, n69633, n69634, n69635, n69636, n69637, n69638, n69639, n69640, n69641, n69642, n69643, n69644, n69645, n69646, n69647, n69648, n69649, n69650, n69651, n69652, n69653, n69654, n69655, n69656, n69657, n69658, n69659, n69660, n69661, n69662, n69663, n69664, n69665, n69666, n69667, n69668, n69669, n69670, n69671, n69672, n69673, n69674, n69675, n69676, n69677, n69678, n69679, n69680, n69681, n69682, n69683, n69684, n69685, n69686, n69687, n69688, n69689, n69690, n69691, n69692, n69693, n69694, n69695, n69696, n69697, n69698, n69699, n69700, n69701, n69702, n69703, n69704, n69705, n69706, n69707, n69708, n69709, n69710, n69711, n69712, n69713, n69714, n69715, n69716, n69717, n69718, n69719, n69720, n69721, n69722, n69723, n69724, n69725, n69726, n69727, n69728, n69729, n69730, n69731, n69732, n69733, n69734, n69735, n69736, n69737, n69738, n69739, n69740, n69741, n69742, n69743, n69744, n69745, n69746, n69747, n69748, n69749, n69750, n69751, n69752, n69753, n69754, n69755, n69756, n69757, n69758, n69759, n69760, n69761, n69762, n69763, n69764, n69765, n69766, n69767, n69768, n69769, n69770, n69771, n69772, n69773, n69774, n69775, n69776, n69777, n69778, n69779, n69780, n69781, n69782, n69783, n69784, n69785, n69786, n69787, n69788, n69789, n69790, n69791, n69792, n69793, n69794, n69795, n69796, n69797, n69798, n69799, n69800, n69801, n69802, n69803, n69804, n69805, n69806, n69807, n69808, n69809, n69810, n69811, n69812, n69813, n69814, n69815, n69816, n69817, n69818, n69819, n69820, n69821, n69822, n69823, n69824, n69825, n69826, n69827, n69828, n69829, n69830, n69831, n69832, n69833, n69834, n69835, n69836, n69837, n69838, n69839, n69840, n69841, n69842, n69843, n69844, n69845, n69846, n69847, n69848, n69849, n69850, n69851, n69852, n69853, n69854, n69855, n69856, n69857, n69858, n69859, n69860, n69861, n69862, n69863, n69864, n69865, n69866, n69867, n69868, n69869, n69870, n69871, n69872, n69873, n69874, n69875, n69876, n69877, n69878, n69879, n69880, n69881, n69882, n69883, n69884, n69885, n69886, n69887, n69888, n69889, n69890, n69891, n69892, n69893, n69894, n69895, n69896, n69897, n69898, n69899, n69900, n69901, n69902, n69903, n69904, n69905, n69906, n69907, n69908, n69909, n69910, n69911, n69912, n69913, n69914, n69915, n69916, n69917, n69918, n69919, n69920, n69921, n69922, n69923, n69924, n69925, n69926, n69927, n69928, n69929, n69930, n69931, n69932, n69933, n69934, n69935, n69936, n69937, n69938, n69939, n69940, n69941, n69942, n69943, n69944, n69945, n69946, n69947, n69948, n69949, n69950, n69951, n69952, n69953, n69954, n69955, n69956, n69957, n69958, n69959, n69960, n69961, n69962, n69963, n69964, n69965, n69966, n69967, n69968, n69969, n69970, n69971, n69972, n69973, n69974, n69975, n69976, n69977, n69978, n69979, n69980, n69981, n69982, n69983, n69984, n69985, n69986, n69987, n69988, n69989, n69990, n69991, n69992, n69993, n69994, n69995, n69996, n69997, n69998, n69999, n70000, n70001, n70002, n70003, n70004, n70005, n70006, n70007, n70008, n70009, n70010, n70011, n70012, n70013, n70014, n70015, n70016, n70017, n70018, n70019, n70020, n70021, n70022, n70023, n70024, n70025, n70026, n70027, n70028, n70029, n70030, n70031, n70032, n70033, n70034, n70035, n70036, n70037, n70038, n70039, n70040, n70041, n70042, n70043, n70044, n70045, n70046, n70047, n70048, n70049, n70050, n70051, n70052, n70053, n70054, n70055, n70056, n70057, n70058, n70059, n70060, n70061, n70062, n70063, n70064, n70065, n70066, n70067, n70068, n70069, n70070, n70071, n70072, n70073, n70074, n70075, n70076, n70077, n70078, n70079, n70080, n70081, n70082, n70083, n70084, n70085, n70086, n70087, n70088, n70089, n70090, n70091, n70092, n70093, n70094, n70095, n70096, n70097, n70098, n70099, n70100, n70101, n70102, n70103, n70104, n70105, n70106, n70107, n70108, n70109, n70110, n70111, n70112, n70113, n70114, n70115, n70116, n70117, n70118, n70119, n70120, n70121, n70122, n70123, n70124, n70125, n70126, n70127, n70128, n70129, n70130, n70131, n70132, n70133, n70134, n70135, n70136, n70137, n70138, n70139, n70140, n70141, n70142, n70143, n70144, n70145, n70146, n70147, n70148, n70149, n70150, n70151, n70152, n70153, n70154, n70155, n70156, n70157, n70158, n70159, n70160, n70161, n70162, n70163, n70164, n70165, n70166, n70167, n70168, n70169, n70170, n70171, n70172, n70173, n70174, n70175, n70176, n70177, n70178, n70179, n70180, n70181, n70182, n70183, n70184, n70185, n70186, n70187, n70188, n70189, n70190, n70191, n70192, n70193, n70194, n70195, n70196, n70197, n70198, n70199, n70200, n70201, n70202, n70203, n70204, n70205, n70206, n70207, n70208, n70209, n70210, n70211, n70212, n70213, n70214, n70215, n70216, n70217, n70218, n70219, n70220, n70221, n70222, n70223, n70224, n70225, n70226, n70227, n70228, n70229, n70230, n70231, n70232, n70233, n70234, n70235, n70236, n70237, n70238, n70239, n70240, n70241, n70242, n70243, n70244, n70245, n70246, n70247, n70248, n70249, n70250, n70251, n70252, n70253, n70254, n70255, n70256, n70257, n70258, n70259, n70260, n70261, n70262, n70263, n70264, n70265, n70266, n70267, n70268, n70269, n70270, n70271, n70272, n70273, n70274, n70275, n70276, n70277, n70278, n70279, n70280, n70281, n70282, n70283, n70284, n70285, n70286, n70287, n70288, n70289, n70290, n70291, n70292, n70293, n70294, n70295, n70296, n70297, n70298, n70299, n70300, n70301, n70302, n70303, n70304, n70305, n70306, n70307, n70308, n70309, n70310, n70311, n70312, n70313, n70314, n70315, n70316, n70317, n70318, n70319, n70320, n70321, n70322, n70323, n70324, n70325, n70326, n70327, n70328, n70329, n70330, n70331, n70332, n70333, n70334, n70335, n70336, n70337, n70338, n70339, n70340, n70341, n70342, n70343, n70344, n70345, n70346, n70347, n70348, n70349, n70350, n70351, n70352, n70353, n70354, n70355, n70356, n70357, n70358, n70359, n70360, n70361, n70362, n70363, n70364, n70365, n70366, n70367, n70368, n70369, n70370, n70371, n70372, n70373, n70374, n70375, n70376, n70377, n70378, n70379, n70380, n70381, n70382, n70383, n70384, n70385, n70386, n70387, n70388, n70389, n70390, n70391, n70392, n70393, n70394, n70395, n70396, n70397, n70398, n70399, n70400, n70401, n70402, n70403, n70404, n70405, n70406, n70407, n70408, n70409, n70410, n70411, n70412, n70413, n70414, n70415, n70416, n70417, n70418, n70419, n70420, n70421, n70422, n70423, n70424, n70425, n70426, n70427, n70428, n70429, n70430, n70431, n70432, n70433, n70434, n70435, n70436, n70437, n70438, n70439, n70440, n70441, n70442, n70443, n70444, n70445, n70446, n70447, n70448, n70449, n70450, n70451, n70452, n70453, n70454, n70455, n70456, n70457, n70458, n70459, n70460, n70461, n70462, n70463, n70464, n70465, n70466, n70467, n70468, n70469, n70470, n70471, n70472, n70473, n70474, n70475, n70476, n70477, n70478, n70479, n70480, n70481, n70482, n70483, n70484, n70485, n70486, n70487, n70488, n70489, n70490, n70491, n70492, n70493, n70494, n70495, n70496, n70497, n70498, n70499, n70500, n70501, n70502, n70503, n70504, n70505, n70506, n70507, n70508, n70509, n70510, n70511, n70512, n70513, n70514, n70515, n70516, n70517, n70518, n70519, n70520, n70521, n70522, n70523, n70524, n70525, n70526, n70527, n70528, n70529, n70530, n70531, n70532, n70533, n70534, n70535, n70536, n70537, n70538, n70539, n70540, n70541, n70542, n70543, n70544, n70545, n70546, n70547, n70548, n70549, n70550, n70551, n70552, n70553, n70554, n70555, n70556, n70557, n70558, n70559, n70560, n70561, n70562, n70563, n70564, n70565, n70566, n70567, n70568, n70569, n70570, n70571, n70572, n70573, n70574, n70575, n70576, n70577, n70578, n70579, n70580, n70581, n70582, n70583, n70584, n70585, n70586, n70587, n70588, n70589, n70590, n70591, n70592, n70593, n70594, n70595, n70596, n70597, n70598, n70599, n70600, n70601, n70602, n70603, n70604, n70605, n70606, n70607, n70608, n70609, n70610, n70611, n70612, n70613, n70614, n70615, n70616, n70617, n70618, n70619, n70620, n70621, n70622, n70623, n70624, n70625, n70626, n70627, n70628, n70629, n70630, n70631, n70632, n70633, n70634, n70635, n70636, n70637, n70638, n70639, n70640, n70641, n70642, n70643, n70644, n70645, n70646, n70647, n70648, n70649, n70650, n70651, n70652, n70653, n70654, n70655, n70656, n70657, n70658, n70659, n70660, n70661, n70662, n70663, n70664, n70665, n70666, n70667, n70668, n70669, n70670, n70671, n70672, n70673, n70674, n70675, n70676, n70677, n70678, n70679, n70680, n70681, n70682, n70683, n70684, n70685, n70686, n70687, n70688, n70689, n70690, n70691, n70692, n70693, n70694, n70695, n70696, n70697, n70698, n70699, n70700, n70701, n70702, n70703, n70704, n70705, n70706, n70707, n70708, n70709, n70710, n70711, n70712, n70713, n70714, n70715, n70716, n70717, n70718, n70719, n70720, n70721, n70722, n70723, n70724, n70725, n70726, n70727, n70728, n70729, n70730, n70731, n70732, n70733, n70734, n70735, n70736, n70737, n70738, n70739, n70740, n70741, n70742, n70743, n70744, n70745, n70746, n70747, n70748, n70749, n70750, n70751, n70752, n70753, n70754, n70755, n70756, n70757, n70758, n70759, n70760, n70761, n70762, n70763, n70764, n70765, n70766, n70767, n70768, n70769, n70770, n70771, n70772, n70773, n70774, n70775, n70776, n70777, n70778, n70779, n70780, n70781, n70782, n70783, n70784, n70785, n70786, n70787, n70788, n70789, n70790, n70791, n70792, n70793, n70794, n70795, n70796, n70797, n70798, n70799, n70800, n70801, n70802, n70803, n70804, n70805, n70806, n70807, n70808, n70809, n70810, n70811, n70812, n70813, n70814, n70815, n70816, n70817, n70818, n70819, n70820, n70821, n70822, n70823, n70824, n70825, n70826, n70827, n70828, n70829, n70830, n70831, n70832, n70833, n70834, n70835, n70836, n70837, n70838, n70839, n70840, n70841, n70842, n70843, n70844, n70845, n70846, n70847, n70848, n70849, n70850, n70851, n70852, n70853, n70854, n70855, n70856, n70857, n70858, n70859, n70860, n70861, n70862, n70863, n70864, n70865, n70866, n70867, n70868, n70869, n70870, n70871, n70872, n70873, n70874, n70875, n70876, n70877, n70878, n70879, n70880, n70881, n70882, n70883, n70884, n70885, n70886, n70887, n70888, n70889, n70890, n70891, n70892, n70893, n70894, n70895, n70896, n70897, n70898, n70899, n70900, n70901, n70902, n70903, n70904, n70905, n70906, n70907, n70908, n70909, n70910, n70911, n70912, n70913, n70914, n70915, n70916, n70917, n70918, n70919, n70920, n70921, n70922, n70923, n70924, n70925, n70926, n70927, n70928, n70929, n70930, n70931, n70932, n70933, n70934, n70935, n70936, n70937, n70938, n70939, n70940, n70941, n70942, n70943, n70944, n70945, n70946, n70947, n70948, n70949, n70950, n70951, n70952, n70953, n70954, n70955, n70956, n70957, n70958, n70959, n70960, n70961, n70962, n70963, n70964, n70965, n70966, n70967, n70968, n70969, n70970, n70971, n70972, n70973, n70974, n70975, n70976, n70977, n70978, n70979, n70980, n70981, n70982, n70983, n70984, n70985, n70986, n70987, n70988, n70989, n70990, n70991, n70992, n70993, n70994, n70995, n70996, n70997, n70998, n70999, n71000, n71001, n71002, n71003, n71004, n71005, n71006, n71007, n71008, n71009, n71010, n71011, n71012, n71013, n71014, n71015, n71016, n71017, n71018, n71019, n71020, n71021, n71022, n71023, n71024, n71025, n71026, n71027, n71028, n71029, n71030, n71031, n71032, n71033, n71034, n71035, n71036, n71037, n71038, n71039, n71040, n71041, n71042, n71043, n71044, n71045, n71046, n71047, n71048, n71049, n71050, n71051, n71052, n71053, n71054, n71055, n71056, n71057, n71058, n71059, n71060, n71061, n71062, n71063, n71064, n71065, n71066, n71067, n71068, n71069, n71070, n71071, n71072, n71073, n71074, n71075, n71076, n71077, n71078, n71079, n71080, n71081, n71082, n71083, n71084, n71085, n71086, n71087, n71088, n71089, n71090, n71091, n71092, n71093, n71094, n71095, n71096, n71097, n71098, n71099, n71100, n71101, n71102, n71103, n71104, n71105, n71106, n71107, n71108, n71109, n71110, n71111, n71112, n71113, n71114, n71115, n71116, n71117, n71118, n71119, n71120, n71121, n71122, n71123, n71124, n71125, n71126, n71127, n71128, n71129, n71130, n71131, n71132, n71133, n71134, n71135, n71136, n71137, n71138, n71139, n71140, n71141, n71142, n71143, n71144, n71145, n71146, n71147, n71148, n71149, n71150, n71151, n71152, n71153, n71154, n71155, n71156, n71157, n71158, n71159, n71160, n71161, n71162, n71163, n71164, n71165, n71166, n71167, n71168, n71169, n71170, n71171, n71172, n71173, n71174, n71175, n71176, n71177, n71178, n71179, n71180, n71181, n71182, n71183, n71184, n71185, n71186, n71187, n71188, n71189, n71190, n71191, n71192, n71193, n71194, n71195, n71196, n71197, n71198, n71199, n71200, n71201, n71202, n71203, n71204, n71205, n71206, n71207, n71208, n71209, n71210, n71211, n71212, n71213, n71214, n71215, n71216, n71217, n71218, n71219, n71220, n71221, n71222, n71223, n71224, n71225, n71226, n71227, n71228, n71229, n71230, n71231, n71232, n71233, n71234, n71235, n71236, n71237, n71238, n71239, n71240, n71241, n71242, n71243, n71244, n71245, n71246, n71247, n71248, n71249, n71250, n71251, n71252, n71253, n71254, n71255, n71256, n71257, n71258, n71259, n71260, n71261, n71262, n71263, n71264, n71265, n71266, n71267, n71268, n71269, n71270, n71271, n71272, n71273, n71274, n71275, n71276, n71277, n71278, n71279, n71280, n71281, n71282, n71283, n71284, n71285, n71286, n71287, n71288, n71289, n71290, n71291, n71292, n71293, n71294, n71295, n71296, n71297, n71298, n71299, n71300, n71301, n71302, n71303, n71304, n71305, n71306, n71307, n71308, n71309, n71310, n71311, n71312, n71313, n71314, n71315, n71316, n71317, n71318, n71319, n71320, n71321, n71322, n71323, n71324, n71325, n71326, n71327, n71328, n71329, n71330, n71331, n71332, n71333, n71334, n71335, n71336, n71337, n71338, n71339, n71340, n71341, n71342, n71343, n71344, n71345, n71346, n71347, n71348, n71349, n71350, n71351, n71352, n71353, n71354, n71355, n71356, n71357, n71358, n71359, n71360, n71361, n71362, n71363, n71364, n71365, n71366, n71367, n71368, n71369, n71370, n71371, n71372, n71373, n71374, n71375, n71376, n71377, n71378, n71379, n71380, n71381, n71382, n71383, n71384, n71385, n71386, n71387, n71388, n71389, n71390, n71391, n71392, n71393, n71394, n71395, n71396, n71397, n71398, n71399, n71400, n71401, n71402, n71403, n71404, n71405, n71406, n71407, n71408, n71409, n71410, n71411, n71412, n71413, n71414, n71415, n71416, n71417, n71418, n71419, n71420, n71421, n71422, n71423, n71424, n71425, n71426, n71427, n71428, n71429, n71430, n71431, n71432, n71433, n71434, n71435, n71436, n71437, n71438, n71439, n71440, n71441, n71442, n71443, n71444, n71445, n71446, n71447, n71448, n71449, n71450, n71451, n71452, n71453, n71454, n71455, n71456, n71457, n71458, n71459, n71460, n71461, n71462, n71463, n71464, n71465, n71466, n71467, n71468, n71469, n71470, n71471, n71472, n71473, n71474, n71475, n71476, n71477, n71478, n71479, n71480, n71481, n71482, n71483, n71484, n71485, n71486, n71487, n71488, n71489, n71490, n71491, n71492, n71493, n71494, n71495, n71496, n71497, n71498, n71499, n71500, n71501, n71502, n71503, n71504, n71505, n71506, n71507, n71508, n71509, n71510, n71511, n71512, n71513, n71514, n71515, n71516, n71517, n71518, n71519, n71520, n71521, n71522, n71523, n71524, n71525, n71526, n71527, n71528, n71529, n71530, n71531, n71532, n71533, n71534, n71535, n71536, n71537, n71538, n71539, n71540, n71541, n71542, n71543, n71544, n71545, n71546, n71547, n71548, n71549, n71550, n71551, n71552, n71553, n71554, n71555, n71556, n71557, n71558, n71559, n71560, n71561, n71562, n71563, n71564, n71565, n71566, n71567, n71568, n71569, n71570, n71571, n71572, n71573, n71574, n71575, n71576, n71577, n71578, n71579, n71580, n71581, n71582, n71583, n71584, n71585, n71586, n71587, n71588, n71589, n71590, n71591, n71592, n71593, n71594, n71595, n71596, n71597, n71598, n71599, n71600, n71601, n71602, n71603, n71604, n71605, n71606, n71607, n71608, n71609, n71610, n71611, n71612, n71613, n71614, n71615, n71616, n71617, n71618, n71619, n71620, n71621, n71622, n71623, n71624, n71625, n71626, n71627, n71628, n71629, n71630, n71631, n71632, n71633, n71634, n71635, n71636, n71637, n71638, n71639, n71640, n71641, n71642, n71643, n71644, n71645, n71646, n71647, n71648, n71649, n71650, n71651, n71652, n71653, n71654, n71655, n71656, n71657, n71658, n71659, n71660, n71661, n71662, n71663, n71664, n71665, n71666, n71667, n71668, n71669, n71670, n71671, n71672, n71673, n71674, n71675, n71676, n71677, n71678, n71679, n71680, n71681, n71682, n71683, n71684, n71685, n71686, n71687, n71688, n71689, n71690, n71691, n71692, n71693, n71694, n71695, n71696, n71697, n71698, n71699, n71700, n71701, n71702, n71703, n71704, n71705, n71706, n71707, n71708, n71709, n71710, n71711, n71712, n71713, n71714, n71715, n71716, n71717, n71718, n71719, n71720, n71721, n71722, n71723, n71724, n71725, n71726, n71727, n71728, n71729, n71730, n71731, n71732, n71733, n71734, n71735, n71736, n71737, n71738, n71739, n71740, n71741, n71742, n71743, n71744, n71745, n71746, n71747, n71748, n71749, n71750, n71751, n71752, n71753, n71754, n71755, n71756, n71757, n71758, n71759, n71760, n71761, n71762, n71763, n71764, n71765, n71766, n71767, n71768, n71769, n71770, n71771, n71772, n71773, n71774, n71775, n71776, n71777, n71778, n71779, n71780, n71781, n71782, n71783, n71784, n71785, n71786, n71787, n71788, n71789, n71790, n71791, n71792, n71793, n71794, n71795, n71796, n71797, n71798, n71799, n71800, n71801, n71802, n71803, n71804, n71805, n71806, n71807, n71808, n71809, n71810, n71811, n71812, n71813, n71814, n71815, n71816, n71817, n71818, n71819, n71820, n71821, n71822, n71823, n71824, n71825, n71826, n71827, n71828, n71829, n71830, n71831, n71832, n71833, n71834, n71835, n71836, n71837, n71838, n71839, n71840, n71841, n71842, n71843, n71844, n71845, n71846, n71847, n71848, n71849, n71850, n71851, n71852, n71853, n71854, n71855, n71856, n71857, n71858, n71859, n71860, n71861, n71862, n71863, n71864, n71865, n71866, n71867, n71868, n71869, n71870, n71871, n71872, n71873, n71874, n71875, n71876, n71877, n71878, n71879, n71880, n71881, n71882, n71883, n71884, n71885, n71886, n71887, n71888, n71889, n71890, n71891, n71892, n71893, n71894, n71895, n71896, n71897, n71898, n71899, n71900, n71901, n71902, n71903, n71904, n71905, n71906, n71907, n71908, n71909, n71910, n71911, n71912, n71913, n71914, n71915, n71916, n71917, n71918, n71919, n71920, n71921, n71922, n71923, n71924, n71925, n71926, n71927, n71928, n71929, n71930, n71931, n71932, n71933, n71934, n71935, n71936, n71937, n71938, n71939, n71940, n71941, n71942, n71943, n71944, n71945, n71946, n71947, n71948, n71949, n71950, n71951, n71952, n71953, n71954, n71955, n71956, n71957, n71958, n71959, n71960, n71961, n71962, n71963, n71964, n71965, n71966, n71967, n71968, n71969, n71970, n71971, n71972, n71973, n71974, n71975, n71976, n71977, n71978, n71979, n71980, n71981, n71982, n71983, n71984, n71985, n71986, n71987, n71988, n71989, n71990, n71991, n71992, n71993, n71994, n71995, n71996, n71997, n71998, n71999, n72000, n72001, n72002, n72003, n72004, n72005, n72006, n72007, n72008, n72009, n72010, n72011, n72012, n72013, n72014, n72015, n72016, n72017, n72018, n72019, n72020, n72021, n72022, n72023, n72024, n72025, n72026, n72027, n72028, n72029, n72030, n72031, n72032, n72033, n72034, n72035, n72036, n72037, n72038, n72039, n72040, n72041, n72042, n72043, n72044, n72045, n72046, n72047, n72048, n72049, n72050, n72051, n72052, n72053, n72054, n72055, n72056, n72057, n72058, n72059, n72060, n72061, n72062, n72063, n72064, n72065, n72066, n72067, n72068, n72069, n72070, n72071, n72072, n72073, n72074, n72075, n72076, n72077, n72078, n72079, n72080, n72081, n72082, n72083, n72084, n72085, n72086, n72087, n72088, n72089, n72090, n72091, n72092, n72093, n72094, n72095, n72096, n72097, n72098, n72099, n72100, n72101, n72102, n72103, n72104, n72105, n72106, n72107, n72108, n72109, n72110, n72111, n72112, n72113, n72114, n72115, n72116, n72117, n72118, n72119, n72120, n72121, n72122, n72123, n72124, n72125, n72126, n72127, n72128, n72129, n72130, n72131, n72132, n72133, n72134, n72135, n72136, n72137, n72138, n72139, n72140, n72141, n72142, n72143, n72144, n72145, n72146, n72147, n72148, n72149, n72150, n72151, n72152, n72153, n72154, n72155, n72156, n72157, n72158, n72159, n72160, n72161, n72162, n72163, n72164, n72165, n72166, n72167, n72168, n72169, n72170, n72171, n72172, n72173, n72174, n72175, n72176, n72177, n72178, n72179, n72180, n72181, n72182, n72183, n72184, n72185, n72186, n72187, n72188, n72189, n72190, n72191, n72192, n72193, n72194, n72195, n72196, n72197, n72198, n72199, n72200, n72201, n72202, n72203, n72204, n72205, n72206, n72207, n72208, n72209, n72210, n72211, n72212, n72213, n72214, n72215, n72216, n72217, n72218, n72219, n72220, n72221, n72222, n72223, n72224, n72225, n72226, n72227, n72228, n72229, n72230, n72231, n72232, n72233, n72234, n72235, n72236, n72237, n72238, n72239, n72240, n72241, n72242, n72243, n72244, n72245, n72246, n72247, n72248, n72249, n72250, n72251, n72252, n72253, n72254, n72255, n72256, n72257, n72258, n72259, n72260, n72261, n72262, n72263, n72264, n72265, n72266, n72267, n72268, n72269, n72270, n72271, n72272, n72273, n72274, n72275, n72276, n72277, n72278, n72279, n72280, n72281, n72282, n72283, n72284, n72285, n72286, n72287, n72288, n72289, n72290, n72291, n72292, n72293, n72294, n72295, n72296, n72297, n72298, n72299, n72300, n72301, n72302, n72303, n72304, n72305, n72306, n72307, n72308, n72309, n72310, n72311, n72312, n72313, n72314, n72315, n72316, n72317, n72318, n72319, n72320, n72321, n72322, n72323, n72324, n72325, n72326, n72327, n72328, n72329, n72330, n72331, n72332, n72333, n72334, n72335, n72336, n72337, n72338, n72339, n72340, n72341, n72342, n72343, n72344, n72345, n72346, n72347, n72348, n72349, n72350, n72351, n72352, n72353, n72354, n72355, n72356, n72357, n72358, n72359, n72360, n72361, n72362, n72363, n72364, n72365, n72366, n72367, n72368, n72369, n72370, n72371, n72372, n72373, n72374, n72375, n72376, n72377, n72378, n72379, n72380, n72381, n72382, n72383, n72384, n72385, n72386, n72387, n72388, n72389, n72390, n72391, n72392, n72393, n72394, n72395, n72396, n72397, n72398, n72399, n72400, n72401, n72402, n72403, n72404, n72405, n72406, n72407, n72408, n72409, n72410, n72411, n72412, n72413, n72414, n72415, n72416, n72417, n72418, n72419, n72420, n72421, n72422, n72423, n72424, n72425, n72426, n72427, n72428, n72429, n72430, n72431, n72432, n72433, n72434, n72435, n72436, n72437, n72438, n72439, n72440, n72441, n72442, n72443, n72444, n72445, n72446, n72447, n72448, n72449, n72450, n72451, n72452, n72453, n72454, n72455, n72456, n72457, n72458, n72459, n72460, n72461, n72462, n72463, n72464, n72465, n72466, n72467, n72468, n72469, n72470, n72471, n72472, n72473, n72474, n72475, n72476, n72477, n72478, n72479, n72480, n72481, n72482, n72483, n72484, n72485, n72486, n72487, n72488, n72489, n72490, n72491, n72492, n72493, n72494, n72495, n72496, n72497, n72498, n72499, n72500, n72501, n72502, n72503, n72504, n72505, n72506, n72507, n72508, n72509, n72510, n72511, n72512, n72513, n72514, n72515, n72516, n72517, n72518, n72519, n72520, n72521, n72522, n72523, n72524, n72525, n72526, n72527, n72528, n72529, n72530, n72531, n72532, n72533, n72534, n72535, n72536, n72537, n72538, n72539, n72540, n72541, n72542, n72543, n72544, n72545, n72546, n72547, n72548, n72549, n72550, n72551, n72552, n72553, n72554, n72555, n72556, n72557, n72558, n72559, n72560, n72561, n72562, n72563, n72564, n72565, n72566, n72567, n72568, n72569, n72570, n72571, n72572, n72573, n72574, n72575, n72576, n72577, n72578, n72579, n72580, n72581, n72582, n72583, n72584, n72585, n72586, n72587, n72588, n72589, n72590, n72591, n72592, n72593, n72594, n72595, n72596, n72597, n72598, n72599, n72600, n72601, n72602, n72603, n72604, n72605, n72606, n72607, n72608, n72609, n72610, n72611, n72612, n72613, n72614, n72615, n72616, n72617, n72618, n72619, n72620, n72621, n72622, n72623, n72624, n72625, n72626, n72627, n72628, n72629, n72630, n72631, n72632, n72633, n72634, n72635, n72636, n72637, n72638, n72639, n72640, n72641, n72642, n72643, n72644, n72645, n72646, n72647, n72648, n72649, n72650, n72651, n72652, n72653, n72654, n72655, n72656, n72657, n72658, n72659, n72660, n72661, n72662, n72663, n72664, n72665, n72666, n72667, n72668, n72669, n72670, n72671, n72672, n72673, n72674, n72675, n72676, n72677, n72678, n72679, n72680, n72681, n72682, n72683, n72684, n72685, n72686, n72687, n72688, n72689, n72690, n72691, n72692, n72693, n72694, n72695, n72696, n72697, n72698, n72699, n72700, n72701, n72702, n72703, n72704, n72705, n72706, n72707, n72708, n72709, n72710, n72711, n72712, n72713, n72714, n72715, n72716, n72717, n72718, n72719, n72720, n72721, n72722, n72723, n72724, n72725, n72726, n72727, n72728, n72729, n72730, n72731, n72732, n72733, n72734, n72735, n72736, n72737, n72738, n72739, n72740, n72741, n72742, n72743, n72744, n72745, n72746, n72747, n72748, n72749, n72750, n72751, n72752, n72753, n72754, n72755, n72756, n72757, n72758, n72759, n72760, n72761, n72762, n72763, n72764, n72765, n72766, n72767, n72768, n72769, n72770, n72771, n72772, n72773, n72774, n72775, n72776, n72777, n72778, n72779, n72780, n72781, n72782, n72783, n72784, n72785, n72786, n72787, n72788, n72789, n72790, n72791, n72792, n72793, n72794, n72795, n72796, n72797, n72798, n72799, n72800, n72801, n72802, n72803, n72804, n72805, n72806, n72807, n72808, n72809, n72810, n72811, n72812, n72813, n72814, n72815, n72816, n72817, n72818, n72819, n72820, n72821, n72822, n72823, n72824, n72825, n72826, n72827, n72828, n72829, n72830, n72831, n72832, n72833, n72834, n72835, n72836, n72837, n72838, n72839, n72840, n72841, n72842, n72843, n72844, n72845, n72846, n72847, n72848, n72849, n72850, n72851, n72852, n72853, n72854, n72855, n72856, n72857, n72858, n72859, n72860, n72861, n72862, n72863, n72864, n72865, n72866, n72867, n72868, n72869, n72870, n72871, n72872, n72873, n72874, n72875, n72876, n72877, n72878, n72879, n72880, n72881, n72882, n72883, n72884, n72885, n72886, n72887, n72888, n72889, n72890, n72891, n72892, n72893, n72894, n72895, n72896, n72897, n72898, n72899, n72900, n72901, n72902, n72903, n72904, n72905, n72906, n72907, n72908, n72909, n72910, n72911, n72912, n72913, n72914, n72915, n72916, n72917, n72918, n72919, n72920, n72921, n72922, n72923, n72924, n72925, n72926, n72927, n72928, n72929, n72930, n72931, n72932, n72933, n72934, n72935, n72936, n72937, n72938, n72939, n72940, n72941, n72942, n72943, n72944, n72945, n72946, n72947, n72948, n72949, n72950, n72951, n72952, n72953, n72954, n72955, n72956, n72957, n72958, n72959, n72960, n72961, n72962, n72963, n72964, n72965, n72966, n72967, n72968, n72969, n72970, n72971, n72972, n72973, n72974, n72975, n72976, n72977, n72978, n72979, n72980, n72981, n72982, n72983, n72984, n72985, n72986, n72987, n72988, n72989, n72990, n72991, n72992, n72993, n72994, n72995, n72996, n72997, n72998, n72999, n73000, n73001, n73002, n73003, n73004, n73005, n73006, n73007, n73008, n73009, n73010, n73011, n73012, n73013, n73014, n73015, n73016, n73017, n73018, n73019, n73020, n73021, n73022, n73023, n73024, n73025, n73026, n73027, n73028, n73029, n73030, n73031, n73032, n73033, n73034, n73035, n73036, n73037, n73038, n73039, n73040, n73041, n73042, n73043, n73044, n73045, n73046, n73047, n73048, n73049, n73050, n73051, n73052, n73053, n73054, n73055, n73056, n73057, n73058, n73059, n73060, n73061, n73062, n73063, n73064, n73065, n73066, n73067, n73068, n73069, n73070, n73071, n73072, n73073, n73074, n73075, n73076, n73077, n73078, n73079, n73080, n73081, n73082, n73083, n73084, n73085, n73086, n73087, n73088, n73089, n73090, n73091, n73092, n73093, n73094, n73095, n73096, n73097, n73098, n73099, n73100, n73101, n73102, n73103, n73104, n73105, n73106, n73107, n73108, n73109, n73110, n73111, n73112, n73113, n73114, n73115, n73116, n73117, n73118, n73119, n73120, n73121, n73122, n73123, n73124, n73125, n73126, n73127, n73128, n73129, n73130, n73131, n73132, n73133, n73134, n73135, n73136, n73137, n73138, n73139, n73140, n73141, n73142, n73143, n73144, n73145, n73146, n73147, n73148, n73149, n73150, n73151, n73152, n73153, n73154, n73155, n73156, n73157, n73158, n73159, n73160, n73161, n73162, n73163, n73164, n73165, n73166, n73167, n73168, n73169, n73170, n73171, n73172, n73173, n73174, n73175, n73176, n73177, n73178, n73179, n73180, n73181, n73182, n73183, n73184, n73185, n73186, n73187, n73188, n73189, n73190, n73191, n73192, n73193, n73194, n73195, n73196, n73197, n73198, n73199, n73200, n73201, n73202, n73203, n73204, n73205, n73206, n73207, n73208, n73209, n73210, n73211, n73212, n73213, n73214, n73215, n73216, n73217, n73218, n73219, n73220, n73221, n73222, n73223, n73224, n73225, n73226, n73227, n73228, n73229, n73230, n73231, n73232, n73233, n73234, n73235, n73236, n73237, n73238, n73239, n73240, n73241, n73242, n73243, n73244, n73245, n73246, n73247, n73248, n73249, n73250, n73251, n73252, n73253, n73254, n73255, n73256, n73257, n73258, n73259, n73260, n73261, n73262, n73263, n73264, n73265, n73266, n73267, n73268, n73269, n73270, n73271, n73272, n73273, n73274, n73275, n73276, n73277, n73278, n73279, n73280, n73281, n73282, n73283, n73284, n73285, n73286, n73287, n73288, n73289, n73290, n73291, n73292, n73293, n73294, n73295, n73296, n73297, n73298, n73299, n73300, n73301, n73302, n73303, n73304, n73305, n73306, n73307, n73308, n73309, n73310, n73311, n73312, n73313, n73314, n73315, n73316, n73317, n73318, n73319, n73320, n73321, n73322, n73323, n73324, n73325, n73326, n73327, n73328, n73329, n73330, n73331, n73332, n73333, n73334, n73335, n73336, n73337, n73338, n73339, n73340, n73341, n73342, n73343, n73344, n73345, n73346, n73347, n73348, n73349, n73350, n73351, n73352, n73353, n73354, n73355, n73356, n73357, n73358, n73359, n73360, n73361, n73362, n73363, n73364, n73365, n73366, n73367, n73368, n73369, n73370, n73371, n73372, n73373, n73374, n73375, n73376, n73377, n73378, n73379, n73380, n73381, n73382, n73383, n73384, n73385, n73386, n73387, n73388, n73389, n73390, n73391, n73392, n73393, n73394, n73395, n73396, n73397, n73398, n73399, n73400, n73401, n73402, n73403, n73404, n73405, n73406, n73407, n73408, n73409, n73410, n73411, n73412, n73413, n73414, n73415, n73416, n73417, n73418, n73419, n73420, n73421, n73422, n73423, n73424, n73425, n73426, n73427, n73428, n73429, n73430, n73431, n73432, n73433, n73434, n73435, n73436, n73437, n73438, n73439, n73440, n73441, n73442, n73443, n73444, n73445, n73446, n73447, n73448, n73449, n73450, n73451, n73452, n73453, n73454, n73455, n73456, n73457, n73458, n73459, n73460, n73461, n73462, n73463, n73464, n73465, n73466, n73467, n73468, n73469, n73470, n73471, n73472, n73473, n73474, n73475, n73476, n73477, n73478, n73479, n73480, n73481, n73482, n73483, n73484, n73485, n73486, n73487, n73488, n73489, n73490, n73491, n73492, n73493, n73494, n73495, n73496, n73497, n73498, n73499, n73500, n73501, n73502, n73503, n73504, n73505, n73506, n73507, n73508, n73509, n73510, n73511, n73512, n73513, n73514, n73515, n73516, n73517, n73518, n73519, n73520, n73521, n73522, n73523, n73524, n73525, n73526, n73527, n73528, n73529, n73530, n73531, n73532, n73533, n73534, n73535, n73536, n73537, n73538, n73539, n73540, n73541, n73542, n73543, n73544, n73545, n73546, n73547, n73548, n73549, n73550, n73551, n73552, n73553, n73554, n73555, n73556, n73557, n73558, n73559, n73560, n73561, n73562, n73563, n73564, n73565, n73566, n73567, n73568, n73569, n73570, n73571, n73572, n73573, n73574, n73575, n73576, n73577, n73578, n73579, n73580, n73581, n73582, n73583, n73584, n73585, n73586, n73587, n73588, n73589, n73590, n73591, n73592, n73593, n73594, n73595, n73596, n73597, n73598, n73599, n73600, n73601, n73602, n73603, n73604, n73605, n73606, n73607, n73608, n73609, n73610, n73611, n73612, n73613, n73614, n73615, n73616, n73617, n73618, n73619, n73620, n73621, n73622, n73623, n73624, n73625, n73626, n73627, n73628, n73629, n73630, n73631, n73632, n73633, n73634, n73635, n73636, n73637, n73638, n73639, n73640, n73641, n73642, n73643, n73644, n73645, n73646, n73647, n73648, n73649, n73650, n73651, n73652, n73653, n73654, n73655, n73656, n73657, n73658, n73659, n73660, n73661, n73662, n73663, n73664, n73665, n73666, n73667, n73668, n73669, n73670, n73671, n73672, n73673, n73674, n73675, n73676, n73677, n73678, n73679, n73680, n73681, n73682, n73683, n73684, n73685, n73686, n73687, n73688, n73689, n73690, n73691, n73692, n73693, n73694, n73695, n73696, n73697, n73698, n73699, n73700, n73701, n73702, n73703, n73704, n73705, n73706, n73707, n73708, n73709, n73710, n73711, n73712, n73713, n73714, n73715, n73716, n73717, n73718, n73719, n73720, n73721, n73722, n73723, n73724, n73725, n73726, n73727, n73728, n73729, n73730, n73731, n73732, n73733, n73734, n73735, n73736, n73737, n73738, n73739, n73740, n73741, n73742, n73743, n73744, n73745, n73746, n73747, n73748, n73749, n73750, n73751, n73752, n73753, n73754, n73755, n73756, n73757, n73758, n73759, n73760, n73761, n73762, n73763, n73764, n73765, n73766, n73767, n73768, n73769, n73770, n73771, n73772, n73773, n73774, n73775, n73776, n73777, n73778, n73779, n73780, n73781, n73782, n73783, n73784, n73785, n73786, n73787, n73788, n73789, n73790, n73791, n73792, n73793, n73794, n73795, n73796, n73797, n73798, n73799, n73800, n73801, n73802, n73803, n73804, n73805, n73806, n73807, n73808, n73809, n73810, n73811, n73812, n73813, n73814, n73815, n73816, n73817, n73818, n73819, n73820, n73821, n73822, n73823, n73824, n73825, n73826, n73827, n73828, n73829, n73830, n73831, n73832, n73833, n73834, n73835, n73836, n73837, n73838, n73839, n73840, n73841, n73842, n73843, n73844, n73845, n73846, n73847, n73848, n73849, n73850, n73851, n73852, n73853, n73854, n73855, n73856, n73857, n73858, n73859, n73860, n73861, n73862, n73863, n73864, n73865, n73866, n73867, n73868, n73869, n73870, n73871, n73872, n73873, n73874, n73875, n73876, n73877, n73878, n73879, n73880, n73881, n73882, n73883, n73884, n73885, n73886, n73887, n73888, n73889, n73890, n73891, n73892, n73893, n73894, n73895, n73896, n73897, n73898, n73899, n73900, n73901, n73902, n73903, n73904, n73905, n73906, n73907, n73908, n73909, n73910, n73911, n73912, n73913, n73914, n73915, n73916, n73917, n73918, n73919, n73920, n73921, n73922, n73923, n73924, n73925, n73926, n73927, n73928, n73929, n73930, n73931, n73932, n73933, n73934, n73935, n73936, n73937, n73938, n73939, n73940, n73941, n73942, n73943, n73944, n73945, n73946, n73947, n73948, n73949, n73950, n73951, n73952, n73953, n73954, n73955, n73956, n73957, n73958, n73959, n73960, n73961, n73962, n73963, n73964, n73965, n73966, n73967, n73968, n73969, n73970, n73971, n73972, n73973, n73974, n73975, n73976, n73977, n73978, n73979, n73980, n73981, n73982, n73983, n73984, n73985, n73986, n73987, n73988, n73989, n73990, n73991, n73992, n73993, n73994, n73995, n73996, n73997, n73998, n73999, n74000, n74001, n74002, n74003, n74004, n74005, n74006, n74007, n74008, n74009, n74010, n74011, n74012, n74013, n74014, n74015, n74016, n74017, n74018, n74019, n74020, n74021, n74022, n74023, n74024, n74025, n74026, n74027, n74028, n74029, n74030, n74031, n74032, n74033, n74034, n74035, n74036, n74037, n74038, n74039, n74040, n74041, n74042, n74043, n74044, n74045, n74046, n74047, n74048, n74049, n74050, n74051, n74052, n74053, n74054, n74055, n74056, n74057, n74058, n74059, n74060, n74061, n74062, n74063, n74064, n74065, n74066, n74067, n74068, n74069, n74070, n74071, n74072, n74073, n74074, n74075, n74076, n74077, n74078, n74079, n74080, n74081, n74082, n74083, n74084, n74085, n74086, n74087, n74088, n74089, n74090, n74091, n74092, n74093, n74094, n74095, n74096, n74097, n74098, n74099, n74100, n74101, n74102, n74103, n74104, n74105, n74106, n74107, n74108, n74109, n74110, n74111, n74112, n74113, n74114, n74115, n74116, n74117, n74118, n74119, n74120, n74121, n74122, n74123, n74124, n74125, n74126, n74127, n74128, n74129, n74130, n74131, n74132, n74133, n74134, n74135, n74136, n74137, n74138, n74139, n74140, n74141, n74142, n74143, n74144, n74145, n74146, n74147, n74148, n74149, n74150, n74151, n74152, n74153, n74154, n74155, n74156, n74157, n74158, n74159, n74160, n74161, n74162, n74163, n74164, n74165, n74166, n74167, n74168, n74169, n74170, n74171, n74172, n74173, n74174, n74175, n74176, n74177, n74178, n74179, n74180, n74181, n74182, n74183, n74184, n74185, n74186, n74187, n74188, n74189, n74190, n74191, n74192, n74193, n74194, n74195, n74196, n74197, n74198, n74199, n74200, n74201, n74202, n74203, n74204, n74205, n74206, n74207, n74208, n74209, n74210, n74211, n74212, n74213, n74214, n74215, n74216, n74217, n74218, n74219, n74220, n74221, n74222, n74223, n74224, n74225, n74226, n74227, n74228, n74229, n74230, n74231, n74232, n74233, n74234, n74235, n74236, n74237, n74238, n74239, n74240, n74241, n74242, n74243, n74244, n74245, n74246, n74247, n74248, n74249, n74250, n74251, n74252, n74253, n74254, n74255, n74256, n74257, n74258, n74259, n74260, n74261, n74262, n74263, n74264, n74265, n74266, n74267, n74268, n74269, n74270, n74271, n74272, n74273, n74274, n74275, n74276, n74277, n74278, n74279, n74280, n74281, n74282, n74283, n74284, n74285, n74286, n74287, n74288, n74289, n74290, n74291, n74292, n74293, n74294, n74295, n74296, n74297, n74298, n74299, n74300, n74301, n74302, n74303, n74304, n74305, n74306, n74307, n74308, n74309, n74310, n74311, n74312, n74313, n74314, n74315, n74316, n74317, n74318, n74319, n74320, n74321, n74322, n74323, n74324, n74325, n74326, n74327, n74328, n74329, n74330, n74331, n74332, n74333, n74334, n74335, n74336, n74337, n74338, n74339, n74340, n74341, n74342, n74343, n74344, n74345, n74346, n74347, n74348, n74349, n74350, n74351, n74352, n74353, n74354, n74355, n74356, n74357, n74358, n74359, n74360, n74361, n74362, n74363, n74364, n74365, n74366, n74367, n74368, n74369, n74370, n74371, n74372, n74373, n74374, n74375, n74376, n74377, n74378, n74379, n74380, n74381, n74382, n74383, n74384, n74385, n74386, n74387, n74388, n74389, n74390, n74391, n74392, n74393, n74394, n74395, n74396, n74397, n74398, n74399, n74400, n74401, n74402, n74403, n74404, n74405, n74406, n74407, n74408, n74409, n74410, n74411, n74412, n74413, n74414, n74415, n74416, n74417, n74418, n74419, n74420, n74421, n74422, n74423, n74424, n74425, n74426, n74427, n74428, n74429, n74430, n74431, n74432, n74433, n74434, n74435, n74436, n74437, n74438, n74439, n74440, n74441, n74442, n74443, n74444, n74445, n74446, n74447, n74448, n74449, n74450, n74451, n74452, n74453, n74454, n74455, n74456, n74457, n74458, n74459, n74460, n74461, n74462, n74463, n74464, n74465, n74466, n74467, n74468, n74469, n74470, n74471, n74472, n74473, n74474, n74475, n74476, n74477, n74478, n74479, n74480, n74481, n74482, n74483, n74484, n74485, n74486, n74487, n74488, n74489, n74490, n74491, n74492, n74493, n74494, n74495, n74496, n74497, n74498, n74499, n74500, n74501, n74502, n74503, n74504, n74505, n74506, n74507, n74508, n74509, n74510, n74511, n74512, n74513, n74514, n74515, n74516, n74517, n74518, n74519, n74520, n74521, n74522, n74523, n74524, n74525, n74526, n74527, n74528, n74529, n74530, n74531, n74532, n74533, n74534, n74535, n74536, n74537, n74538, n74539, n74540, n74541, n74542, n74543, n74544, n74545, n74546, n74547, n74548, n74549, n74550, n74551, n74552, n74553, n74554, n74555, n74556, n74557, n74558, n74559, n74560, n74561, n74562, n74563, n74564, n74565, n74566, n74567, n74568, n74569, n74570, n74571, n74572, n74573, n74574, n74575, n74576, n74577, n74578, n74579, n74580, n74581, n74582, n74583, n74584, n74585, n74586, n74587, n74588, n74589, n74590, n74591, n74592, n74593, n74594, n74595, n74596, n74597, n74598, n74599, n74600, n74601, n74602, n74603, n74604, n74605, n74606, n74607, n74608, n74609, n74610, n74611, n74612, n74613, n74614, n74615, n74616, n74617, n74618, n74619, n74620, n74621, n74622, n74623, n74624, n74625, n74626, n74627, n74628, n74629, n74630, n74631, n74632, n74633, n74634, n74635, n74636, n74637, n74638, n74639, n74640, n74641, n74642, n74643, n74644, n74645, n74646, n74647, n74648, n74649, n74650, n74651, n74652, n74653, n74654, n74655, n74656, n74657, n74658, n74659, n74660, n74661, n74662, n74663, n74664, n74665, n74666, n74667, n74668, n74669, n74670, n74671, n74672, n74673, n74674, n74675, n74676, n74677, n74678, n74679, n74680, n74681, n74682, n74683, n74684, n74685, n74686, n74687, n74688, n74689, n74690, n74691, n74692, n74693, n74694, n74695, n74696, n74697, n74698, n74699, n74700, n74701, n74702, n74703, n74704, n74705, n74706, n74707, n74708, n74709, n74710, n74711, n74712, n74713, n74714, n74715, n74716, n74717, n74718, n74719, n74720, n74721, n74722, n74723, n74724, n74725, n74726, n74727, n74728, n74729, n74730, n74731, n74732, n74733, n74734, n74735, n74736, n74737, n74738, n74739, n74740, n74741, n74742, n74743, n74744, n74745, n74746, n74747, n74748, n74749, n74750, n74751, n74752, n74753, n74754, n74755, n74756, n74757, n74758, n74759, n74760, n74761, n74762, n74763, n74764, n74765, n74766, n74767, n74768, n74769, n74770, n74771, n74772, n74773, n74774, n74775, n74776, n74777, n74778, n74779, n74780, n74781, n74782, n74783, n74784, n74785, n74786, n74787, n74788, n74789, n74790, n74791, n74792, n74793, n74794, n74795, n74796, n74797, n74798, n74799, n74800, n74801, n74802, n74803, n74804, n74805, n74806, n74807, n74808, n74809, n74810, n74811, n74812, n74813, n74814, n74815, n74816, n74817, n74818, n74819, n74820, n74821, n74822, n74823, n74824, n74825, n74826, n74827, n74828, n74829, n74830, n74831, n74832, n74833, n74834, n74835, n74836, n74837, n74838, n74839, n74840, n74841, n74842, n74843, n74844, n74845, n74846, n74847, n74848, n74849, n74850, n74851, n74852, n74853, n74854, n74855, n74856, n74857, n74858, n74859, n74860, n74861, n74862, n74863, n74864, n74865, n74866, n74867, n74868, n74869, n74870, n74871, n74872, n74873, n74874, n74875, n74876, n74877, n74878, n74879, n74880, n74881, n74882, n74883, n74884, n74885, n74886, n74887, n74888, n74889, n74890, n74891, n74892, n74893, n74894, n74895, n74896, n74897, n74898, n74899, n74900, n74901, n74902, n74903, n74904, n74905, n74906, n74907, n74908, n74909, n74910, n74911, n74912, n74913, n74914, n74915, n74916, n74917, n74918, n74919, n74920, n74921, n74922, n74923, n74924, n74925, n74926, n74927, n74928, n74929, n74930, n74931, n74932, n74933, n74934, n74935, n74936, n74937, n74938, n74939, n74940, n74941, n74942, n74943, n74944, n74945, n74946, n74947, n74948, n74949, n74950, n74951, n74952, n74953, n74954, n74955, n74956, n74957, n74958, n74959, n74960, n74961, n74962, n74963, n74964, n74965, n74966, n74967, n74968, n74969, n74970, n74971, n74972, n74973, n74974, n74975, n74976, n74977, n74978, n74979, n74980, n74981, n74982, n74983, n74984, n74985, n74986, n74987, n74988, n74989, n74990, n74991, n74992, n74993, n74994, n74995, n74996, n74997, n74998, n74999, n75000, n75001, n75002, n75003, n75004, n75005, n75006, n75007, n75008, n75009, n75010, n75011, n75012, n75013, n75014, n75015, n75016, n75017, n75018, n75019, n75020, n75021, n75022, n75023, n75024, n75025, n75026, n75027, n75028, n75029, n75030, n75031, n75032, n75033, n75034, n75035, n75036, n75037, n75038, n75039, n75040, n75041, n75042, n75043, n75044, n75045, n75046, n75047, n75048, n75049, n75050, n75051, n75052, n75053, n75054, n75055, n75056, n75057, n75058, n75059, n75060, n75061, n75062, n75063, n75064, n75065, n75066, n75067, n75068, n75069, n75070, n75071, n75072, n75073, n75074, n75075, n75076, n75077, n75078, n75079, n75080, n75081, n75082, n75083, n75084, n75085, n75086, n75087, n75088, n75089, n75090, n75091, n75092, n75093, n75094, n75095, n75096, n75097, n75098, n75099, n75100, n75101, n75102, n75103, n75104, n75105, n75106, n75107, n75108, n75109, n75110, n75111, n75112, n75113, n75114, n75115, n75116, n75117, n75118, n75119, n75120, n75121, n75122, n75123, n75124, n75125, n75126, n75127, n75128, n75129, n75130, n75131, n75132, n75133, n75134, n75135, n75136, n75137, n75138, n75139, n75140, n75141, n75142, n75143, n75144, n75145, n75146, n75147, n75148, n75149, n75150, n75151, n75152, n75153, n75154, n75155, n75156, n75157, n75158, n75159, n75160, n75161, n75162, n75163, n75164, n75165, n75166, n75167, n75168, n75169, n75170, n75171, n75172, n75173, n75174, n75175, n75176, n75177, n75178, n75179, n75180, n75181, n75182, n75183, n75184, n75185, n75186, n75187, n75188, n75189, n75190, n75191, n75192, n75193, n75194, n75195, n75196, n75197, n75198, n75199, n75200, n75201, n75202, n75203, n75204, n75205, n75206, n75207, n75208, n75209, n75210, n75211, n75212, n75213, n75214, n75215, n75216, n75217, n75218, n75219, n75220, n75221, n75222, n75223, n75224, n75225, n75226, n75227, n75228, n75229, n75230, n75231, n75232, n75233, n75234, n75235, n75236, n75237, n75238, n75239, n75240, n75241, n75242, n75243, n75244, n75245, n75246, n75247, n75248, n75249, n75250, n75251, n75252, n75253, n75254, n75255, n75256, n75257, n75258, n75259, n75260, n75261, n75262, n75263, n75264, n75265, n75266, n75267, n75268, n75269, n75270, n75271, n75272, n75273, n75274, n75275, n75276, n75277, n75278, n75279, n75280, n75281, n75282, n75283, n75284, n75285, n75286, n75287, n75288, n75289, n75290, n75291, n75292, n75293, n75294, n75295, n75296, n75297, n75298, n75299, n75300, n75301, n75302, n75303, n75304, n75305, n75306, n75307, n75308, n75309, n75310, n75311, n75312, n75313, n75314, n75315, n75316, n75317, n75318, n75319, n75320, n75321, n75322, n75323, n75324, n75325, n75326, n75327, n75328, n75329, n75330, n75331, n75332, n75333, n75334, n75335, n75336, n75337, n75338, n75339, n75340, n75341, n75342, n75343, n75344, n75345, n75346, n75347, n75348, n75349, n75350, n75351, n75352, n75353, n75354, n75355, n75356, n75357, n75358, n75359, n75360, n75361, n75362, n75363, n75364, n75365, n75366, n75367, n75368, n75369, n75370, n75371, n75372, n75373, n75374, n75375, n75376, n75377, n75378, n75379, n75380, n75381, n75382, n75383, n75384, n75385, n75386, n75387, n75388, n75389, n75390, n75391, n75392, n75393, n75394, n75395, n75396, n75397, n75398, n75399, n75400, n75401, n75402, n75403, n75404, n75405, n75406, n75407, n75408, n75409, n75410, n75411, n75412, n75413, n75414, n75415, n75416, n75417, n75418, n75419, n75420, n75421, n75422, n75423, n75424, n75425, n75426, n75427, n75428, n75429, n75430, n75431, n75432, n75433, n75434, n75435, n75436, n75437, n75438, n75439, n75440, n75441, n75442, n75443, n75444, n75445, n75446, n75447, n75448, n75449, n75450, n75451, n75452, n75453, n75454, n75455, n75456, n75457, n75458, n75459, n75460, n75461, n75462, n75463, n75464, n75465, n75466, n75467, n75468, n75469, n75470, n75471, n75472, n75473, n75474, n75475, n75476, n75477, n75478, n75479, n75480, n75481, n75482, n75483, n75484, n75485, n75486, n75487, n75488, n75489, n75490, n75491, n75492, n75493, n75494, n75495, n75496, n75497, n75498, n75499, n75500, n75501, n75502, n75503, n75504, n75505, n75506, n75507, n75508, n75509, n75510, n75511, n75512, n75513, n75514, n75515, n75516, n75517, n75518, n75519, n75520, n75521, n75522, n75523, n75524, n75525, n75526, n75527, n75528, n75529, n75530, n75531, n75532, n75533, n75534, n75535, n75536, n75537, n75538, n75539, n75540, n75541, n75542, n75543, n75544, n75545, n75546, n75547, n75548, n75549, n75550, n75551, n75552, n75553, n75554, n75555, n75556, n75557, n75558, n75559, n75560, n75561, n75562, n75563, n75564, n75565, n75566, n75567, n75568, n75569, n75570, n75571, n75572, n75573, n75574, n75575, n75576, n75577, n75578, n75579, n75580, n75581, n75582, n75583, n75584, n75585, n75586, n75587, n75588, n75589, n75590, n75591, n75592, n75593, n75594, n75595, n75596, n75597, n75598, n75599, n75600, n75601, n75602, n75603, n75604, n75605, n75606, n75607, n75608, n75609, n75610, n75611, n75612, n75613, n75614, n75615, n75616, n75617, n75618, n75619, n75620, n75621, n75622, n75623, n75624, n75625, n75626, n75627, n75628, n75629, n75630, n75631, n75632, n75633, n75634, n75635, n75636, n75637, n75638, n75639, n75640, n75641, n75642, n75643, n75644, n75645, n75646, n75647, n75648, n75649, n75650, n75651, n75652, n75653, n75654, n75655, n75656, n75657, n75658, n75659, n75660, n75661, n75662, n75663, n75664, n75665, n75666, n75667, n75668, n75669, n75670, n75671, n75672, n75673, n75674, n75675, n75676, n75677, n75678, n75679, n75680, n75681, n75682, n75683, n75684, n75685, n75686, n75687, n75688, n75689, n75690, n75691, n75692, n75693, n75694, n75695, n75696, n75697, n75698, n75699, n75700, n75701, n75702, n75703, n75704, n75705, n75706, n75707, n75708, n75709, n75710, n75711, n75712, n75713, n75714, n75715, n75716, n75717, n75718, n75719, n75720, n75721, n75722, n75723, n75724, n75725, n75726, n75727, n75728, n75729, n75730, n75731, n75732, n75733, n75734, n75735, n75736, n75737, n75738, n75739, n75740, n75741, n75742, n75743, n75744, n75745, n75746, n75747, n75748, n75749, n75750, n75751, n75752, n75753, n75754, n75755, n75756, n75757, n75758, n75759, n75760, n75761, n75762, n75763, n75764, n75765, n75766, n75767, n75768, n75769, n75770, n75771, n75772, n75773, n75774, n75775, n75776, n75777, n75778, n75779, n75780, n75781, n75782, n75783, n75784, n75785, n75786, n75787, n75788, n75789, n75790, n75791, n75792, n75793, n75794, n75795, n75796, n75797, n75798, n75799, n75800, n75801, n75802, n75803, n75804, n75805, n75806, n75807, n75808, n75809, n75810, n75811, n75812, n75813, n75814, n75815, n75816, n75817, n75818, n75819, n75820, n75821, n75822, n75823, n75824, n75825, n75826, n75827, n75828, n75829, n75830, n75831, n75832, n75833, n75834, n75835, n75836, n75837, n75838, n75839, n75840, n75841, n75842, n75843, n75844, n75845, n75846, n75847, n75848, n75849, n75850, n75851, n75852, n75853, n75854, n75855, n75856, n75857, n75858, n75859, n75860, n75861, n75862, n75863, n75864, n75865, n75866, n75867, n75868, n75869, n75870, n75871, n75872, n75873, n75874, n75875, n75876, n75877, n75878, n75879, n75880, n75881, n75882, n75883, n75884, n75885, n75886, n75887, n75888, n75889, n75890, n75891, n75892, n75893, n75894, n75895, n75896, n75897, n75898, n75899, n75900, n75901, n75902, n75903, n75904, n75905, n75906, n75907, n75908, n75909, n75910, n75911, n75912, n75913, n75914, n75915, n75916, n75917, n75918, n75919, n75920, n75921, n75922, n75923, n75924, n75925, n75926, n75927, n75928, n75929, n75930, n75931, n75932, n75933, n75934, n75935, n75936, n75937, n75938, n75939, n75940, n75941, n75942, n75943, n75944, n75945, n75946, n75947, n75948, n75949, n75950, n75951, n75952, n75953, n75954, n75955, n75956, n75957, n75958, n75959, n75960, n75961, n75962, n75963, n75964, n75965, n75966, n75967, n75968, n75969, n75970, n75971, n75972, n75973, n75974, n75975, n75976, n75977, n75978, n75979, n75980, n75981, n75982, n75983, n75984, n75985, n75986, n75987, n75988, n75989, n75990, n75991, n75992, n75993, n75994, n75995, n75996, n75997, n75998, n75999, n76000, n76001, n76002, n76003, n76004, n76005, n76006, n76007, n76008, n76009, n76010, n76011, n76012, n76013, n76014, n76015, n76016, n76017, n76018, n76019, n76020, n76021, n76022, n76023, n76024, n76025, n76026, n76027, n76028, n76029, n76030, n76031, n76032, n76033, n76034, n76035, n76036, n76037, n76038, n76039, n76040, n76041, n76042, n76043, n76044, n76045, n76046, n76047, n76048, n76049, n76050, n76051, n76052, n76053, n76054, n76055, n76056, n76057, n76058, n76059, n76060, n76061, n76062, n76063, n76064, n76065, n76066, n76067, n76068, n76069, n76070, n76071, n76072, n76073, n76074, n76075, n76076, n76077, n76078, n76079, n76080, n76081, n76082, n76083, n76084, n76085, n76086, n76087, n76088, n76089, n76090, n76091, n76092, n76093, n76094, n76095, n76096, n76097, n76098, n76099, n76100, n76101, n76102, n76103, n76104, n76105, n76106, n76107, n76108, n76109, n76110, n76111, n76112, n76113, n76114, n76115, n76116, n76117, n76118, n76119, n76120, n76121, n76122, n76123, n76124, n76125, n76126, n76127, n76128, n76129, n76130, n76131, n76132, n76133, n76134, n76135, n76136, n76137, n76138, n76139, n76140, n76141, n76142, n76143, n76144, n76145, n76146, n76147, n76148, n76149, n76150, n76151, n76152, n76153, n76154, n76155, n76156, n76157, n76158, n76159, n76160, n76161, n76162, n76163, n76164, n76165, n76166, n76167, n76168, n76169, n76170, n76171, n76172, n76173, n76174, n76175, n76176, n76177, n76178, n76179, n76180, n76181, n76182, n76183, n76184, n76185, n76186, n76187, n76188, n76189, n76190, n76191, n76192, n76193, n76194, n76195, n76196, n76197, n76198, n76199, n76200, n76201, n76202, n76203, n76204, n76205, n76206, n76207, n76208, n76209, n76210, n76211, n76212, n76213, n76214, n76215, n76216, n76217, n76218, n76219, n76220, n76221, n76222, n76223, n76224, n76225, n76226, n76227, n76228, n76229, n76230, n76231, n76232, n76233, n76234, n76235, n76236, n76237, n76238, n76239, n76240, n76241, n76242, n76243, n76244, n76245, n76246, n76247, n76248, n76249, n76250, n76251, n76252, n76253, n76254, n76255, n76256, n76257, n76258, n76259, n76260, n76261, n76262, n76263, n76264, n76265, n76266, n76267, n76268, n76269, n76270, n76271, n76272, n76273, n76274, n76275, n76276, n76277, n76278, n76279, n76280, n76281, n76282, n76283, n76284, n76285, n76286, n76287, n76288, n76289, n76290, n76291, n76292, n76293, n76294, n76295, n76296, n76297, n76298, n76299, n76300, n76301, n76302, n76303, n76304, n76305, n76306, n76307, n76308, n76309, n76310, n76311, n76312, n76313, n76314, n76315, n76316, n76317, n76318, n76319, n76320, n76321, n76322, n76323, n76324, n76325, n76326, n76327, n76328, n76329, n76330, n76331, n76332, n76333, n76334, n76335, n76336, n76337, n76338, n76339, n76340, n76341, n76342, n76343, n76344, n76345, n76346, n76347, n76348, n76349, n76350, n76351, n76352, n76353, n76354, n76355, n76356, n76357, n76358, n76359, n76360, n76361, n76362, n76363, n76364, n76365, n76366, n76367, n76368, n76369, n76370, n76371, n76372, n76373, n76374, n76375, n76376, n76377, n76378, n76379, n76380, n76381, n76382, n76383, n76384, n76385, n76386, n76387, n76388, n76389, n76390, n76391, n76392, n76393, n76394, n76395, n76396, n76397, n76398, n76399, n76400, n76401, n76402, n76403, n76404, n76405, n76406, n76407, n76408, n76409, n76410, n76411, n76412, n76413, n76414, n76415, n76416, n76417, n76418, n76419, n76420, n76421, n76422, n76423, n76424, n76425, n76426, n76427, n76428, n76429, n76430, n76431, n76432, n76433, n76434, n76435, n76436, n76437, n76438, n76439, n76440, n76441, n76442, n76443, n76444, n76445, n76446, n76447, n76448, n76449, n76450, n76451, n76452, n76453, n76454, n76455, n76456, n76457, n76458, n76459, n76460, n76461, n76462, n76463, n76464, n76465, n76466, n76467, n76468, n76469, n76470, n76471, n76472, n76473, n76474, n76475, n76476, n76477, n76478, n76479, n76480, n76481, n76482, n76483, n76484, n76485, n76486, n76487, n76488, n76489, n76490, n76491, n76492, n76493, n76494, n76495, n76496, n76497, n76498, n76499, n76500, n76501, n76502, n76503, n76504, n76505, n76506, n76507, n76508, n76509, n76510, n76511, n76512, n76513, n76514, n76515, n76516, n76517, n76518, n76519, n76520, n76521, n76522, n76523, n76524, n76525, n76526, n76527, n76528, n76529, n76530, n76531, n76532, n76533, n76534, n76535, n76536, n76537, n76538, n76539, n76540, n76541, n76542, n76543, n76544, n76545, n76546, n76547, n76548, n76549, n76550, n76551, n76552, n76553, n76554, n76555, n76556, n76557, n76558, n76559, n76560, n76561, n76562, n76563, n76564, n76565, n76566, n76567, n76568, n76569, n76570, n76571, n76572, n76573, n76574, n76575, n76576, n76577, n76578, n76579, n76580, n76581, n76582, n76583, n76584, n76585, n76586, n76587, n76588, n76589, n76590, n76591, n76592, n76593, n76594, n76595, n76596, n76597, n76598, n76599, n76600, n76601, n76602, n76603, n76604, n76605, n76606, n76607, n76608, n76609, n76610, n76611, n76612, n76613, n76614, n76615, n76616, n76617, n76618, n76619, n76620, n76621, n76622, n76623, n76624, n76625, n76626, n76627, n76628, n76629, n76630, n76631, n76632, n76633, n76634, n76635, n76636, n76637, n76638, n76639, n76640, n76641, n76642, n76643, n76644, n76645, n76646, n76647, n76648, n76649, n76650, n76651, n76652, n76653, n76654, n76655, n76656, n76657, n76658, n76659, n76660, n76661, n76662, n76663, n76664, n76665, n76666, n76667, n76668, n76669, n76670, n76671, n76672, n76673, n76674, n76675, n76676, n76677, n76678, n76679, n76680, n76681, n76682, n76683, n76684, n76685, n76686, n76687, n76688, n76689, n76690, n76691, n76692, n76693, n76694, n76695, n76696, n76697, n76698, n76699, n76700, n76701, n76702, n76703, n76704, n76705, n76706, n76707, n76708, n76709, n76710, n76711, n76712, n76713, n76714, n76715, n76716, n76717, n76718, n76719, n76720, n76721, n76722, n76723, n76724, n76725, n76726, n76727, n76728, n76729, n76730, n76731, n76732, n76733, n76734, n76735, n76736, n76737, n76738, n76739, n76740, n76741, n76742, n76743, n76744, n76745, n76746, n76747, n76748, n76749, n76750, n76751, n76752, n76753, n76754, n76755, n76756, n76757, n76758, n76759, n76760, n76761, n76762, n76763, n76764, n76765, n76766, n76767, n76768, n76769, n76770, n76771, n76772, n76773, n76774, n76775, n76776, n76777, n76778, n76779, n76780, n76781, n76782, n76783, n76784, n76785, n76786, n76787, n76788, n76789, n76790, n76791, n76792, n76793, n76794, n76795, n76796, n76797, n76798, n76799, n76800, n76801, n76802, n76803, n76804, n76805, n76806, n76807, n76808, n76809, n76810, n76811, n76812, n76813, n76814, n76815, n76816, n76817, n76818, n76819, n76820, n76821, n76822, n76823, n76824, n76825, n76826, n76827, n76828, n76829, n76830, n76831, n76832, n76833, n76834, n76835, n76836, n76837, n76838, n76839, n76840, n76841, n76842, n76843, n76844, n76845, n76846, n76847, n76848, n76849, n76850, n76851, n76852, n76853, n76854, n76855, n76856, n76857, n76858, n76859, n76860, n76861, n76862, n76863, n76864, n76865, n76866, n76867, n76868, n76869, n76870, n76871, n76872, n76873, n76874, n76875, n76876, n76877, n76878, n76879, n76880, n76881, n76882, n76883, n76884, n76885, n76886, n76887, n76888, n76889, n76890, n76891, n76892, n76893, n76894, n76895, n76896, n76897, n76898, n76899, n76900, n76901, n76902, n76903, n76904, n76905, n76906, n76907, n76908, n76909, n76910, n76911, n76912, n76913, n76914, n76915, n76916, n76917, n76918, n76919, n76920, n76921, n76922, n76923, n76924, n76925, n76926, n76927, n76928, n76929, n76930, n76931, n76932, n76933, n76934, n76935, n76936, n76937, n76938, n76939, n76940, n76941, n76942, n76943, n76944, n76945, n76946, n76947, n76948, n76949, n76950, n76951, n76952, n76953, n76954, n76955, n76956, n76957, n76958, n76959, n76960, n76961, n76962, n76963, n76964, n76965, n76966, n76967, n76968, n76969, n76970, n76971, n76972, n76973, n76974, n76975, n76976, n76977, n76978, n76979, n76980, n76981, n76982, n76983, n76984, n76985, n76986, n76987, n76988, n76989, n76990, n76991, n76992, n76993, n76994, n76995, n76996, n76997, n76998, n76999, n77000, n77001, n77002, n77003, n77004, n77005, n77006, n77007, n77008, n77009, n77010, n77011, n77012, n77013, n77014, n77015, n77016, n77017, n77018, n77019, n77020, n77021, n77022, n77023, n77024, n77025, n77026, n77027, n77028, n77029, n77030, n77031, n77032, n77033, n77034, n77035, n77036, n77037, n77038, n77039, n77040, n77041, n77042, n77043, n77044, n77045, n77046, n77047, n77048, n77049, n77050, n77051, n77052, n77053, n77054, n77055, n77056, n77057, n77058, n77059, n77060, n77061, n77062, n77063, n77064, n77065, n77066, n77067, n77068, n77069, n77070, n77071, n77072, n77073, n77074, n77075, n77076, n77077, n77078, n77079, n77080, n77081, n77082, n77083, n77084, n77085, n77086, n77087, n77088, n77089, n77090, n77091, n77092, n77093, n77094, n77095, n77096, n77097, n77098, n77099, n77100, n77101, n77102, n77103, n77104, n77105, n77106, n77107, n77108, n77109, n77110, n77111, n77112, n77113, n77114, n77115, n77116, n77117, n77118, n77119, n77120, n77121, n77122, n77123, n77124, n77125, n77126, n77127, n77128, n77129, n77130, n77131, n77132, n77133, n77134, n77135, n77136, n77137, n77138, n77139, n77140, n77141, n77142, n77143, n77144, n77145, n77146, n77147, n77148, n77149, n77150, n77151, n77152, n77153, n77154, n77155, n77156, n77157, n77158, n77159, n77160, n77161, n77162, n77163, n77164, n77165, n77166, n77167, n77168, n77169, n77170, n77171, n77172, n77173, n77174, n77175, n77176, n77177, n77178, n77179, n77180, n77181, n77182, n77183, n77184, n77185, n77186, n77187, n77188, n77189, n77190, n77191, n77192, n77193, n77194, n77195, n77196, n77197, n77198, n77199, n77200, n77201, n77202, n77203, n77204, n77205, n77206, n77207, n77208, n77209, n77210, n77211, n77212, n77213, n77214, n77215, n77216, n77217, n77218, n77219, n77220, n77221, n77222, n77223, n77224, n77225, n77226, n77227, n77228, n77229, n77230, n77231, n77232, n77233, n77234, n77235, n77236, n77237, n77238, n77239, n77240, n77241, n77242, n77243, n77244, n77245, n77246, n77247, n77248, n77249, n77250, n77251, n77252, n77253, n77254, n77255, n77256, n77257, n77258, n77259, n77260, n77261, n77262, n77263, n77264, n77265, n77266, n77267, n77268, n77269, n77270, n77271, n77272, n77273, n77274, n77275, n77276, n77277, n77278, n77279, n77280, n77281, n77282, n77283, n77284, n77285, n77286, n77287, n77288, n77289, n77290, n77291, n77292, n77293, n77294, n77295, n77296, n77297, n77298, n77299, n77300, n77301, n77302, n77303, n77304, n77305, n77306, n77307, n77308, n77309, n77310, n77311, n77312, n77313, n77314, n77315, n77316, n77317, n77318, n77319, n77320, n77321, n77322, n77323, n77324, n77325, n77326, n77327, n77328, n77329, n77330, n77331, n77332, n77333, n77334, n77335, n77336, n77337, n77338, n77339, n77340, n77341, n77342, n77343, n77344, n77345, n77346, n77347, n77348, n77349, n77350, n77351, n77352, n77353, n77354, n77355, n77356, n77357, n77358, n77359, n77360, n77361, n77362, n77363, n77364, n77365, n77366, n77367, n77368, n77369, n77370, n77371, n77372, n77373, n77374, n77375, n77376, n77377, n77378, n77379, n77380, n77381, n77382, n77383, n77384, n77385, n77386, n77387, n77388, n77389, n77390, n77391, n77392, n77393, n77394, n77395, n77396, n77397, n77398, n77399, n77400, n77401, n77402, n77403, n77404, n77405, n77406, n77407, n77408, n77409, n77410, n77411, n77412, n77413, n77414, n77415, n77416, n77417, n77418, n77419, n77420, n77421, n77422, n77423, n77424, n77425, n77426, n77427, n77428, n77429, n77430, n77431, n77432, n77433, n77434, n77435, n77436, n77437, n77438, n77439, n77440, n77441, n77442, n77443, n77444, n77445, n77446, n77447, n77448, n77449, n77450, n77451, n77452, n77453, n77454, n77455, n77456, n77457, n77458, n77459, n77460, n77461, n77462, n77463, n77464, n77465, n77466, n77467, n77468, n77469, n77470, n77471, n77472, n77473, n77474, n77475, n77476, n77477, n77478, n77479, n77480, n77481, n77482, n77483, n77484, n77485, n77486, n77487, n77488, n77489, n77490, n77491, n77492, n77493, n77494, n77495, n77496, n77497, n77498, n77499, n77500, n77501, n77502, n77503, n77504, n77505, n77506, n77507, n77508, n77509, n77510, n77511, n77512, n77513, n77514, n77515, n77516, n77517, n77518, n77519, n77520, n77521, n77522, n77523, n77524, n77525, n77526, n77527, n77528, n77529, n77530, n77531, n77532, n77533, n77534, n77535, n77536, n77537, n77538, n77539, n77540, n77541, n77542, n77543, n77544, n77545, n77546, n77547, n77548, n77549, n77550, n77551, n77552, n77553, n77554, n77555, n77556, n77557, n77558, n77559, n77560, n77561, n77562, n77563, n77564, n77565, n77566, n77567, n77568, n77569, n77570, n77571, n77572, n77573, n77574, n77575, n77576, n77577, n77578, n77579, n77580, n77581, n77582, n77583, n77584, n77585, n77586, n77587, n77588, n77589, n77590, n77591, n77592, n77593, n77594, n77595, n77596, n77597, n77598, n77599, n77600, n77601, n77602, n77603, n77604, n77605, n77606, n77607, n77608, n77609, n77610, n77611, n77612, n77613, n77614, n77615, n77616, n77617, n77618, n77619, n77620, n77621, n77622, n77623, n77624, n77625, n77626, n77627, n77628, n77629, n77630, n77631, n77632, n77633, n77634, n77635, n77636, n77637, n77638, n77639, n77640, n77641, n77642, n77643, n77644, n77645, n77646, n77647, n77648, n77649, n77650, n77651, n77652, n77653, n77654, n77655, n77656, n77657, n77658, n77659, n77660, n77661, n77662, n77663, n77664, n77665, n77666, n77667, n77668, n77669, n77670, n77671, n77672, n77673, n77674, n77675, n77676, n77677, n77678, n77679, n77680, n77681, n77682, n77683, n77684, n77685, n77686, n77687, n77688, n77689, n77690, n77691, n77692, n77693, n77694, n77695, n77696, n77697, n77698, n77699, n77700, n77701, n77702, n77703, n77704, n77705, n77706, n77707, n77708, n77709, n77710, n77711, n77712, n77713, n77714, n77715, n77716, n77717, n77718, n77719, n77720, n77721, n77722, n77723, n77724, n77725, n77726, n77727, n77728, n77729, n77730, n77731, n77732, n77733, n77734, n77735, n77736, n77737, n77738, n77739, n77740, n77741, n77742, n77743, n77744, n77745, n77746, n77747, n77748, n77749, n77750, n77751, n77752, n77753, n77754, n77755, n77756, n77757, n77758, n77759, n77760, n77761, n77762, n77763, n77764, n77765, n77766, n77767, n77768, n77769, n77770, n77771, n77772, n77773, n77774, n77775, n77776, n77777, n77778, n77779, n77780, n77781, n77782, n77783, n77784, n77785, n77786, n77787, n77788, n77789, n77790, n77791, n77792, n77793, n77794, n77795, n77796, n77797, n77798, n77799, n77800, n77801, n77802, n77803, n77804, n77805, n77806, n77807, n77808, n77809, n77810, n77811, n77812, n77813, n77814, n77815, n77816, n77817, n77818, n77819, n77820, n77821, n77822, n77823, n77824, n77825, n77826, n77827, n77828, n77829, n77830, n77831, n77832, n77833, n77834, n77835, n77836, n77837, n77838, n77839, n77840, n77841, n77842, n77843, n77844, n77845, n77846, n77847, n77848, n77849, n77850, n77851, n77852, n77853, n77854, n77855, n77856, n77857, n77858, n77859, n77860, n77861, n77862, n77863, n77864, n77865, n77866, n77867, n77868, n77869, n77870, n77871, n77872, n77873, n77874, n77875, n77876, n77877, n77878, n77879, n77880, n77881, n77882, n77883, n77884, n77885, n77886, n77887, n77888, n77889, n77890, n77891, n77892, n77893, n77894, n77895, n77896, n77897, n77898, n77899, n77900, n77901, n77902, n77903, n77904, n77905, n77906, n77907, n77908, n77909, n77910, n77911, n77912, n77913, n77914, n77915, n77916, n77917, n77918, n77919, n77920, n77921, n77922, n77923, n77924, n77925, n77926, n77927, n77928, n77929, n77930, n77931, n77932, n77933, n77934, n77935, n77936, n77937, n77938, n77939, n77940, n77941, n77942, n77943, n77944, n77945, n77946, n77947, n77948, n77949, n77950, n77951, n77952, n77953, n77954, n77955, n77956, n77957, n77958, n77959, n77960, n77961, n77962, n77963, n77964, n77965, n77966, n77967, n77968, n77969, n77970, n77971, n77972, n77973, n77974, n77975, n77976, n77977, n77978, n77979, n77980, n77981, n77982, n77983, n77984, n77985, n77986, n77987, n77988, n77989, n77990, n77991, n77992, n77993, n77994, n77995, n77996, n77997, n77998, n77999, n78000, n78001, n78002, n78003, n78004, n78005, n78006, n78007, n78008, n78009, n78010, n78011, n78012, n78013, n78014, n78015, n78016, n78017, n78018, n78019, n78020, n78021, n78022, n78023, n78024, n78025, n78026, n78027, n78028, n78029, n78030, n78031, n78032, n78033, n78034, n78035, n78036, n78037, n78038, n78039, n78040, n78041, n78042, n78043, n78044, n78045, n78046, n78047, n78048, n78049, n78050, n78051, n78052, n78053, n78054, n78055, n78056, n78057, n78058, n78059, n78060, n78061, n78062, n78063, n78064, n78065, n78066, n78067, n78068, n78069, n78070, n78071, n78072, n78073, n78074, n78075, n78076, n78077, n78078, n78079, n78080, n78081, n78082, n78083, n78084, n78085, n78086, n78087, n78088, n78089, n78090, n78091, n78092, n78093, n78094, n78095, n78096, n78097, n78098, n78099, n78100, n78101, n78102, n78103, n78104, n78105, n78106, n78107, n78108, n78109, n78110, n78111, n78112, n78113, n78114, n78115, n78116, n78117, n78118, n78119, n78120, n78121, n78122, n78123, n78124, n78125, n78126, n78127, n78128, n78129, n78130, n78131, n78132, n78133, n78134, n78135, n78136, n78137, n78138, n78139, n78140, n78141, n78142, n78143, n78144, n78145, n78146, n78147, n78148, n78149, n78150, n78151, n78152, n78153, n78154, n78155, n78156, n78157, n78158, n78159, n78160, n78161, n78162, n78163, n78164, n78165, n78166, n78167, n78168, n78169, n78170, n78171, n78172, n78173, n78174, n78175, n78176, n78177, n78178, n78179, n78180, n78181, n78182, n78183, n78184, n78185, n78186, n78187, n78188, n78189, n78190, n78191, n78192, n78193, n78194, n78195, n78196, n78197, n78198, n78199, n78200, n78201, n78202, n78203, n78204, n78205, n78206, n78207, n78208, n78209, n78210, n78211, n78212, n78213, n78214, n78215, n78216, n78217, n78218, n78219, n78220, n78221, n78222, n78223, n78224, n78225, n78226, n78227, n78228, n78229, n78230, n78231, n78232, n78233, n78234, n78235, n78236, n78237, n78238, n78239, n78240, n78241, n78242, n78243, n78244;
  assign n10199 = ~n273;
  assign n8554 = ~n197;
  assign n3384 = ~n66;
  assign n11822 = ~n41;
  assign n3229 = ~n78;
  assign n7342 = ~n219;
  assign n17111 = ~n160;
  assign n4032 = ~n370;
  assign n10917 = ~n61;
  assign n13481 = ~n324;
  assign n15109 = ~n415;
  assign n20271 = ~n18;
  assign n21353 = ~n2;
  assign n15486 = ~n392;
  assign n15399 = ~n406;
  assign n3342 = ~n65;
  assign n9753 = ~n485;
  assign n20341 = ~n20;
  assign n11437 = ~n260;
  assign n11500 = ~n52;
  assign n7047 = ~n430;
  assign n5391 = ~n148;
  assign n5602 = ~n137;
  assign n17141 = ~n473;
  assign n2896 = ~n86;
  assign n18263 = ~n462;
  assign n14752 = ~n101;
  assign n12343 = ~n35;
  assign n16051 = ~n190;
  assign n18294 = ~n463;
  assign n14988 = ~n412;
  assign n7900 = ~n212;
  assign n8851 = ~n510;
  assign n15473 = ~n407;
  assign n20920 = ~n13;
  assign n14200 = ~n119;
  assign n14245 = ~n104;
  assign n5793 = ~n442;
  assign n18788 = ~n253;
  assign n9219 = ~n503;
  assign n3578 = ~n378;
  assign n8128 = ~n202;
  assign n12900 = ~n341;
  assign n1703 = ~n298;
  assign n12057 = ~n47;
  assign n18051 = ~n456;
  assign n10065 = ~n286;
  assign n19414 = ~n236;
  assign n18899 = ~n240;
  assign n1678 = ~n297;
  assign n10723 = ~n268;
  assign n1118 = ~n319;
  assign n15638 = ~n185;
  assign n15157 = ~n400;
  assign n20137 = ~n31;
  assign n3280 = ~n79;
  assign n10398 = ~n278;
  assign n2975 = ~n72;
  assign n16911 = ~n172;
  assign n12610 = ~n38;
  assign n14600 = ~n97;
  assign n16277 = ~n177;
  assign n2139 = ~n91;
  assign n17578 = ~n166;
  assign n11934 = ~n44;
  assign n9976 = ~n284;
  assign n17182 = ~n161;
  assign n10140 = ~n272;
  assign n12996 = ~n343;
  assign n16739 = ~n168;
  assign n17352 = ~n476;
  assign n7252 = ~n218;
  assign n6467 = ~n132;
  assign n1423 = ~n308;
  assign n11173 = ~n48;
  assign n17956 = ~n470;
  assign n13293 = ~n335;
  assign n7930 = ~n213;
  assign n11976 = ~n45;
  assign n7981 = ~n214;
  assign n19971 = ~n27;
  assign n14879 = ~n409;
  assign n1797 = ~n300;
  assign n21237 = ~n1;
  assign n4506 = ~n365;
  assign n14678 = ~n99;
  assign n10627 = ~n267;
  assign n6815 = ~n424;
  assign n11752 = ~n40;
  assign n13365 = ~n321;
  assign n19641 = ~n226;
  assign n5509 = ~n151;
  assign n19179 = ~n246;
  assign n16311 = ~n387;
  assign n15296 = ~n403;
  assign n3502 = ~n377;
  assign n20442 = ~n22;
  assign n8981 = ~n497;
  assign n3315 = ~n64;
  assign n20485 = ~n23;
  assign n20775 = ~n11;
  assign n2910 = ~n87;
  assign n1764 = ~n299;
  assign n3911 = ~n383;
  assign n7794 = ~n210;
  assign n10976 = ~n271;
  assign n8944 = ~n496;
  assign n9407 = ~n491;
  assign n20295 = ~n19;
  assign n10703 = ~n58;
  assign n12021 = ~n46;
  assign n8745 = ~n508;
  assign n840 = ~n315;
  assign n1201 = ~n305;
  assign n6432 = ~n434;
  assign n13964 = ~n113;
  assign n5464 = ~n150;
  assign n11154 = ~n257;
  assign n19695 = ~n227;
  assign n3604 = ~n69;
  assign n15327 = ~n404;
  assign n3056 = ~n74;
  assign n14942 = ~n411;
  assign n9791 = ~n486;
  assign n13918 = ~n112;
  assign n13017 = ~n328;
  assign n19881 = ~n25;
  assign n19197 = ~n247;
  assign n3736 = ~n380;
  assign n19742 = ~n229;
  assign n9421 = ~n492;
  assign n1450 = ~n309;
  assign n12647 = ~n336;
  assign n13411 = ~n322;
  assign n16246 = ~n386;
  assign n18693 = ~n251;
  assign n4257 = ~n375;
  assign n3849 = ~n382;
  assign n9304 = ~n489;
  assign n8495 = ~n196;
  assign n14316 = ~n106;
  assign n8167 = ~n203;
  assign n5544 = ~n136;
  assign n13253 = ~n334;
  assign n10044 = ~n285;
  assign n4169 = ~n373;
  assign n4928 = ~n358;
  assign n11658 = ~n54;
  assign n3182 = ~n77;
  assign n15251 = ~n402;
  assign n7122 = ~n416;
  assign n13583 = ~n121;
  assign n18124 = ~n458;
  assign n7015 = ~n429;
  assign n14171 = ~n118;
  assign n7384 = ~n221;
  assign n5708 = ~n441;
  assign n9577 = ~n480;
  assign n13745 = ~n124;
  assign n12231 = ~n34;
  assign n11352 = ~n50;
  assign n15572 = ~n394;
  assign n10522 = ~n265;
  assign n13543 = ~n325;
  assign n901 = ~n316;
  assign n15056 = ~n413;
  assign n9544 = ~n495;
  assign n7559 = ~n223;
  assign n16633 = ~n182;
  assign n9015 = ~n498;
  assign n4376 = ~n362;
  assign n8239 = ~n205;
  assign n2766 = ~n83;
  assign n2323 = ~n93;
  assign n4471 = ~n364;
  assign n792 = ~n314;
  assign n17487 = ~n165;
  assign n8358 = ~n192;
  assign n8107 = ~n201;
  assign n6144 = ~n446;
  assign n15732 = ~n396;
  assign n4067 = ~n371;
  assign n12352 = ~n348;
  assign n15067 = ~n414;
  assign n19533 = ~n239;
  assign n8392 = ~n193;
  assign n19809 = ~n230;
  assign n9908 = ~n282;
  assign n18199 = ~n460;
  assign n20607 = ~n9;
  assign n17901 = ~n469;
  assign n8617 = ~n198;
  assign n20542 = ~n8;
  assign n13171 = ~n331;
  assign n17859 = ~n468;
  assign n13098 = ~n330;
  assign n18888 = ~n255;
  assign n13622 = ~n122;
  assign n4683 = ~n353;
  assign n1922 = ~n303;
  assign n9697 = ~n483;
  assign n19596 = ~n225;
  assign n1356 = ~n307;
  assign n5179 = ~n159;
  assign n5088 = ~n157;
  assign n5311 = ~n146;
  assign n10269 = ~n275;
  assign n6286 = ~n130;
  assign n13222 = ~n333;
  assign n7437 = ~n420;
  assign n4120 = ~n372;
  assign n2109 = ~n290;
  assign n21168 = ~n0;
  assign n10788 = ~n59;
  assign n13776 = ~n125;
  assign n8425 = ~n194;
  assign n18144 = ~n459;
  assign n12199 = ~n346;
  assign n18335 = ~n448;
  assign n5130 = ~n158;
  assign n7609 = ~n422;
  assign n13593 = ~n326;
  assign n9721 = ~n484;
  assign n3990 = ~n369;
  assign n17983 = ~n471;
  assign n18218 = ~n461;
  assign n17816 = ~n467;
  assign n3431 = ~n67;
  assign n6678 = ~n438;
  assign n17421 = ~n164;
  assign n5626 = ~n138;
  assign n19360 = ~n235;
  assign n14061 = ~n115;
  assign n78244 = ~n7;
  assign n12170 = ~n33;
  assign n18450 = ~n451;
  assign n14563 = ~n96;
  assign n18059 = ~n457;
  assign n6633 = ~n134;
  assign n15813 = ~n397;
  assign n11429 = ~n51;
  assign n10589 = ~n266;
  assign n7117 = ~n431;
  assign n16437 = ~n179;
  assign n13319 = ~n320;
  assign n18650 = ~n454;
  assign n6920 = ~n427;
  assign n10372 = ~n277;
  assign n2009 = ~n288;
  assign n17004 = ~n174;
  assign n9936 = ~n283;
  assign n16551 = ~n389;
  assign n1286 = ~n306;
  assign n9262 = ~n488;
  assign n6946 = ~n428;
  assign n15210 = ~n401;
  assign n2069 = ~n289;
  assign n1874 = ~n302;
  assign n12118 = ~n32;
  assign n12503 = ~n350;
  assign n14640 = ~n98;
  assign n8583 = ~n505;
  assign n9619 = ~n481;
  assign n18624 = ~n250;
  assign n9190 = ~n502;
  assign n10418 = ~n279;
  assign n4295 = ~n360;
  assign n9098 = ~n500;
  assign n3787 = ~n381;
  assign n1618 = ~n296;
  assign n17431 = ~n477;
  assign n13196 = ~n332;
  assign n9510 = ~n494;
  assign n21468 = ~n4;
  assign n4762 = ~n355;
  assign n18839 = ~n254;
  assign n5860 = ~n443;
  assign n5959 = ~n142;
  assign n18500 = ~n452;
  assign n7523 = ~n421;
  assign n6709 = ~n439;
  assign n16715 = ~n183;
  assign n7845 = ~n211;
  assign n4867 = ~n357;
  assign n8797 = ~n509;
  assign n8015 = ~n215;
  assign n6508 = ~n435;
  assign n18389 = ~n449;
  assign n13075 = ~n329;
  assign n8665 = ~n507;
  assign n16558 = ~n181;
  assign n15860 = ~n188;
  assign n1168 = ~n304;
  assign n4727 = ~n354;
  assign n17333 = ~n163;
  assign n4334 = ~n361;
  assign n1559 = ~n311;
  assign n6577 = ~n436;
  assign n13696 = ~n123;
  assign n15671 = ~n186;
  assign n14072 = ~n116;
  assign n3634 = ~n379;
  assign n9459 = ~n493;
  assign n12940 = ~n342;
  assign n9663 = ~n482;
  assign n1025 = ~n318;
  assign n3147 = ~n76;
  assign n14810 = ~n102;
  assign n19279 = ~n233;
  assign n16510 = ~n180;
  assign n1851 = ~n301;
  assign n17696 = ~n465;
  assign n5423 = ~n149;
  assign n20204 = ~n16;
  assign n7536 = ~n222;
  assign n21721 = ~n6;
  assign n4635 = ~n352;
  assign n19483 = ~n238;
  assign n11263 = ~n49;
  assign n9138 = ~n501;
  assign n12313 = ~n347;
  assign n19125 = ~n245;
  assign n17044 = ~n175;
  assign n8895 = ~n511;
  assign n11085 = ~n256;
  assign n16646 = ~n390;
  assign n7333 = ~n419;
  assign n2783 = ~n84;
  assign n4556 = ~n366;
  assign n16378 = ~n178;
  assign n12533 = ~n37;
  assign n17570 = ~n479;
  assign n12419 = ~n36;
  assign n8067 = ~n200;
  assign n1507 = ~n310;
  assign n15354 = ~n405;
  assign n5010 = ~n155;
  assign n3685 = ~n70;
  assign n14111 = ~n117;
  assign n14710 = ~n100;
  assign n15897 = ~n398;
  assign n5352 = ~n147;
  assign n12617 = ~n351;
  assign n10623 = ~n57;
  assign n12734 = ~n337;
  assign n14279 = ~n105;
  assign n12147 = ~n345;
  assign n16859 = ~n170;
  assign n2621 = ~n81;
  assign n10216 = ~n274;
  assign n11627 = ~n262;
  assign n20052 = ~n29;
  assign n746 = ~n313;
  assign n16793 = ~n169;
  assign n6316 = ~n433;
  assign n2210 = ~n291;
  assign n3965 = ~n368;
  assign n17666 = ~n464;
  assign n10873 = ~n60;
  assign n10470 = ~n264;
  assign n2826 = ~n85;
  assign n11714 = ~n55;
  assign n18542 = ~n453;
  assign n17747 = ~n466;
  assign n4987 = ~n154;
  assign n21407 = ~n3;
  assign n16072 = ~n384;
  assign n19316 = ~n234;
  assign n12767 = ~n338;
  assign n19255 = ~n232;
  assign n3021 = ~n73;
  assign n20212 = ~n17;
  assign n17249 = ~n162;
  assign n11867 = ~n42;
  assign n2082 = ~n90;
  assign n9053 = ~n499;
  assign n19565 = ~n224;
  assign n16229 = ~n176;
  assign n2338 = ~n292;
  assign n9894 = ~n281;
  assign n10097 = ~n287;
  assign n20006 = ~n28;
  assign n2673 = ~n82;
  assign n2545 = ~n294;
  assign n3531 = ~n68;
  assign n12444 = ~n349;
  assign n7185 = ~n217;
  assign n18956 = ~n241;
  assign n14517 = ~n111;
  assign n7273 = ~n418;
  assign n12857 = ~n340;
  assign n5694 = ~n139;
  assign n18410 = ~n450;
  assign n14910 = ~n410;
  assign n8227 = ~n204;
  assign n15529 = ~n393;
  assign n4218 = ~n374;
  assign n21670 = ~n5;
  assign n6045 = ~n143;
  assign n5747 = ~n140;
  assign n18560 = ~n249;
  assign n6372 = ~n131;
  assign n7227 = ~n417;
  assign n14377 = ~n107;
  assign n6535 = ~n133;
  assign n19000 = ~n242;
  assign n2483 = ~n95;
  assign n17477 = ~n478;
  assign n2593 = ~n80;
  assign n8317 = ~n207;
  assign n11895 = ~n43;
  assign n7684 = ~n208;
  assign n2430 = ~n293;
  assign n16138 = ~n385;
  assign n20379 = ~n21;
  assign n6018 = ~n445;
  assign n6214 = ~n129;
  assign n20836 = ~n12;
  assign n2398 = ~n94;
  assign n16960 = ~n173;
  assign n5852 = ~n141;
  assign n14397 = ~n108;
  assign n16084 = ~n191;
  assign n10999 = ~n62;
  assign n11134 = ~n63;
  assign n8474 = ~n195;
  assign n12818 = ~n339;
  assign n15662 = ~n395;
  assign n4946 = ~n153;
  assign n7739 = ~n209;
  assign n2029 = ~n89;
  assign n14444 = ~n109;
  assign n13832 = ~n126;
  assign n11582 = ~n53;
  assign n18712 = ~n252;
  assign n16887 = ~n171;
  assign n10896 = ~n270;
  assign n4592 = ~n367;
  assign n15777 = ~n187;
  assign n6878 = ~n426;
  assign n7394 = ~n220;
  assign n15951 = ~n189;
  assign n20683 = ~n10;
  assign n17168 = ~n474;
  assign n6136 = ~n128;
  assign n11492 = ~n261;
  assign n5261 = ~n145;
  assign n4824 = ~n356;
  assign n17233 = ~n475;
  assign n16413 = ~n388;
  assign n19082 = ~n244;
  assign n9340 = ~n490;
  assign n13439 = ~n323;
  assign n21044 = ~n15;
  assign n10806 = ~n269;
  assign n2217 = ~n92;
  assign n970 = ~n317;
  assign n8278 = ~n206;
  assign n20098 = ~n30;
  assign n14006 = ~n114;
  assign n13893 = ~n127;
  assign n5208 = ~n144;
  assign n3117 = ~n75;
  assign n15958 = ~n399;
  assign n6292 = ~n432;
  assign n6844 = ~n425;
  assign n5043 = ~n156;
  assign n14497 = ~n110;
  assign n6169 = ~n447;
  assign n5930 = ~n444;
  assign n10334 = ~n276;
  assign n8632 = ~n506;
  assign n19432 = ~n237;
  assign n11226 = ~n258;
  assign n6625 = ~n437;
  assign n19716 = ~n228;
  assign n4427 = ~n363;
  assign n11347 = ~n259;
  assign n20935 = ~n14;
  assign n19943 = ~n26;
  assign n19042 = ~n243;
  assign n78243 = n78244 & n21721;
  assign n78242 = n78243 & n21670;
  assign n78056 = ~n78243;
  assign n78054 = n78242 ^ n21468;
  assign n78241 = n78242 & n21468;
  assign n78064 = n5 ^ n78056;
  assign n78240 = n78241 ^ n21407;
  assign n78239 = n78241 & n21407;
  assign n78053 = ~n78054;
  assign n78060 = ~n78064;
  assign n78235 = n78239 ^ n21353;
  assign n78051 = n78240 & n78054;
  assign n78238 = ~n78240;
  assign n78236 = n78239 & n21353;
  assign n78230 = n78051 & n78235;
  assign n78233 = n78236 ^ n21237;
  assign n78232 = n78236 & n21237;
  assign n78237 = n78238 & n78053;
  assign n78034 = ~n78051;
  assign n78234 = ~n78235;
  assign n78227 = n0 ^ n78232;
  assign n78226 = n78230 & n78233;
  assign n78016 = n78051 ^ n78234;
  assign n78229 = n78232 & n21168;
  assign n78231 = ~n78233;
  assign n78036 = ~n78237;
  assign n77977 = n78226 ^ n78227;
  assign n78223 = n15 ^ n78229;
  assign n78004 = n78230 ^ n78231;
  assign n78225 = n78229 & n21044;
  assign n78228 = ~n78226;
  assign n77979 = ~n77977;
  assign n78220 = n14 ^ n78225;
  assign n78002 = ~n78004;
  assign n78224 = n78225 & n20935;
  assign n78222 = n78228 & n78227;
  assign n77965 = n78222 ^ n78223;
  assign n78215 = n78224 ^ n20920;
  assign n78221 = n78224 & n20920;
  assign n78219 = n78222 & n78223;
  assign n77943 = n78219 ^ n78220;
  assign n78211 = n12 ^ n78221;
  assign n78217 = n78219 & n78220;
  assign n78218 = ~n78215;
  assign n78216 = n78221 & n20836;
  assign n77959 = ~n77965;
  assign n78208 = n11 ^ n78216;
  assign n77931 = n78217 ^ n78218;
  assign n78213 = n78216 & n20775;
  assign n77945 = ~n77943;
  assign n78214 = ~n78217;
  assign n78205 = n78213 ^ n20683;
  assign n77928 = ~n77931;
  assign n78209 = n78213 & n20683;
  assign n78210 = n78214 & n78215;
  assign n77866 = n9 ^ n78209;
  assign n78206 = n78209 & n20607;
  assign n77907 = n78210 ^ n78211;
  assign n78202 = ~n78205;
  assign n78212 = ~n78210;
  assign n78197 = n78206 ^ n20542;
  assign n78203 = n78206 & n20542;
  assign n78207 = n78212 & n78211;
  assign n78190 = n23 ^ n78203;
  assign n78200 = n78203 & n20485;
  assign n78194 = ~n78197;
  assign n77892 = n78207 ^ n78208;
  assign n78201 = n78207 & n78208;
  assign n78187 = n78200 ^ n20442;
  assign n78198 = n78200 & n20442;
  assign n77882 = n78201 ^ n78202;
  assign n77902 = ~n77892;
  assign n78204 = ~n78201;
  assign n78180 = n21 ^ n78198;
  assign n78184 = ~n78187;
  assign n78195 = n78198 & n20379;
  assign n77880 = ~n77882;
  assign n77849 = n78204 & n78205;
  assign n78176 = n78195 ^ n20341;
  assign n78192 = n78195 & n20341;
  assign n78199 = ~n77849;
  assign n78170 = n19 ^ n78192;
  assign n78188 = n78192 & n20295;
  assign n78174 = ~n78176;
  assign n78193 = n78199 & n77866;
  assign n78164 = n78188 ^ n20271;
  assign n78185 = n78188 & n20271;
  assign n77853 = n78193 ^ n78194;
  assign n78196 = ~n78193;
  assign n78161 = n78185 ^ n20212;
  assign n78182 = n78185 & n20212;
  assign n78167 = ~n78164;
  assign n78189 = n78196 & n78197;
  assign n78156 = n16 ^ n78182;
  assign n78160 = ~n78161;
  assign n78178 = n78182 & n20204;
  assign n77837 = n78189 ^ n78190;
  assign n78191 = ~n78189;
  assign n78152 = n78178 ^ n20137;
  assign n78177 = n78178 & n20137;
  assign n78183 = n78191 & n78190;
  assign n78150 = n78177 ^ n20098;
  assign n78172 = n78177 & n20098;
  assign n78154 = ~n78152;
  assign n77829 = n78183 ^ n78184;
  assign n78186 = ~n78183;
  assign n78147 = n78172 ^ n20052;
  assign n78168 = n78172 & n20052;
  assign n78149 = ~n78150;
  assign n78179 = n78186 & n78187;
  assign n78143 = n28 ^ n78168;
  assign n78146 = ~n78147;
  assign n78165 = n78168 & n20006;
  assign n77818 = n78179 ^ n78180;
  assign n78181 = ~n78179;
  assign n78137 = n78165 ^ n19971;
  assign n78162 = n78165 & n19971;
  assign n78173 = n78181 & n78180;
  assign n78130 = n26 ^ n78162;
  assign n78158 = n78162 & n19943;
  assign n78140 = ~n78137;
  assign n77811 = n78173 ^ n78174;
  assign n78175 = ~n78173;
  assign n78123 = n25 ^ n78158;
  assign n78099 = n78158 & n19881;
  assign n78169 = n78175 & n78176;
  assign n78118 = ~n78123;
  assign n77796 = n78169 ^ n78170;
  assign n78171 = ~n78169;
  assign n78166 = n78171 & n78170;
  assign n77788 = n78166 ^ n78167;
  assign n78163 = ~n78166;
  assign n77782 = ~n77788;
  assign n78159 = n78163 & n78164;
  assign n77766 = n78159 ^ n78160;
  assign n78157 = n78159 & n78161;
  assign n77740 = n78157 ^ n78156;
  assign n77764 = ~n77766;
  assign n78155 = ~n78157;
  assign n78153 = n78155 & n78156;
  assign n77732 = n78153 ^ n78154;
  assign n78151 = ~n78153;
  assign n78148 = n78151 & n78152;
  assign n76199 = n78148 ^ n78149;
  assign n78145 = n78148 & n78150;
  assign n77230 = n39 ^ n76199;
  assign n78141 = n78145 ^ n78146;
  assign n78142 = n78145 & n78147;
  assign n76204 = ~n76199;
  assign n76103 = n78141 ^ n76199;
  assign n78138 = n78142 ^ n78143;
  assign n78134 = n78141 & n76199;
  assign n77999 = ~n77230;
  assign n78113 = n76204 & n39;
  assign n78144 = ~n78142;
  assign n76009 = n78134 ^ n78138;
  assign n78133 = n76103 & n38;
  assign n76115 = ~n76103;
  assign n78135 = ~n78138;
  assign n78139 = n78144 & n78143;
  assign n78110 = ~n78133;
  assign n76085 = ~n76009;
  assign n78132 = n76115 & n12610;
  assign n78128 = n78134 & n78135;
  assign n78127 = n78139 ^ n78140;
  assign n78136 = ~n78139;
  assign n78095 = n76115 ^ n76085;
  assign n78079 = n76085 & n76103;
  assign n75948 = n78128 ^ n78127;
  assign n78125 = ~n78132;
  assign n78126 = ~n78128;
  assign n78129 = n78136 & n78137;
  assign n78119 = n78079 & n36;
  assign n78112 = n78125 & n78110;
  assign n78124 = n78125 & n78113;
  assign n76006 = ~n75948;
  assign n78114 = ~n78079;
  assign n78115 = n78126 & n78127;
  assign n78116 = n78129 ^ n78130;
  assign n78131 = ~n78129;
  assign n77207 = n78112 ^ n78113;
  assign n78111 = n78114 & n12419;
  assign n75861 = n78115 ^ n78116;
  assign n78067 = ~n78119;
  assign n78109 = ~n78124;
  assign n78121 = ~n78116;
  assign n78120 = ~n78115;
  assign n78122 = n78131 & n78130;
  assign n78058 = n78079 ^ n75861;
  assign n78093 = n75861 & n78079;
  assign n77980 = ~n77207;
  assign n78102 = n78109 & n78110;
  assign n75942 = ~n75861;
  assign n78076 = ~n78111;
  assign n78106 = n78120 & n78121;
  assign n78107 = n78122 ^ n78123;
  assign n78117 = ~n78122;
  assign n78097 = n78058 & n12343;
  assign n78098 = ~n78058;
  assign n78094 = n78102 ^ n78095;
  assign n78103 = n78102 & n12533;
  assign n75836 = n78106 ^ n78107;
  assign n78104 = ~n78102;
  assign n78108 = ~n78107;
  assign n78105 = n78117 & n78118;
  assign n78084 = n37 ^ n78094;
  assign n78045 = ~n78097;
  assign n78091 = n78098 & n35;
  assign n75834 = ~n75836;
  assign n78096 = ~n78103;
  assign n78101 = n78104 & n37;
  assign n78100 = n24 ^ n78105;
  assign n78089 = n78106 & n78108;
  assign n77961 = n78084 ^ n77980;
  assign n78048 = n78084 & n77980;
  assign n78039 = ~n78091;
  assign n78086 = n78093 ^ n75834;
  assign n78092 = n78095 & n78096;
  assign n78080 = n75834 & n78093;
  assign n78090 = n78099 ^ n78100;
  assign n78088 = ~n78101;
  assign n77165 = ~n77961;
  assign n78047 = ~n78048;
  assign n78085 = n78086 & n12231;
  assign n75703 = n78089 ^ n78090;
  assign n78025 = ~n78086;
  assign n78082 = n78089 & n78090;
  assign n78087 = ~n78092;
  assign n77992 = n78080 ^ n75703;
  assign n75627 = n7 ^ n78082;
  assign n77948 = n75703 & n78080;
  assign n78081 = n78025 & n34;
  assign n75757 = ~n75703;
  assign n78029 = ~n78085;
  assign n78077 = n78082 & n7;
  assign n78083 = ~n78082;
  assign n78078 = n78087 & n78088;
  assign n78068 = n77992 & n12170;
  assign n78070 = ~n77992;
  assign n78071 = n77948 & n32;
  assign n75683 = ~n75627;
  assign n78072 = n78077 & n6;
  assign n78069 = n78078 ^ n78079;
  assign n78040 = ~n77948;
  assign n78009 = ~n78081;
  assign n78073 = n78083 & n7;
  assign n78075 = ~n78078;
  assign n77997 = ~n78068;
  assign n78049 = n36 ^ n78069;
  assign n78061 = n78070 & n33;
  assign n77936 = ~n78071;
  assign n78065 = n78040 & n12118;
  assign n78063 = ~n78072;
  assign n78059 = n78073 & n21721;
  assign n78074 = n78075 & n78076;
  assign n77159 = n78048 ^ n78049;
  assign n78046 = ~n78049;
  assign n75466 = n78059 ^ n78060;
  assign n77973 = ~n78061;
  assign n78052 = n78059 & n78064;
  assign n77954 = ~n78065;
  assign n78062 = ~n78059;
  assign n78066 = ~n78074;
  assign n77946 = ~n77159;
  assign n78031 = n78046 & n78047;
  assign n75387 = n78052 ^ n78053;
  assign n75525 = ~n75466;
  assign n78050 = ~n78052;
  assign n78055 = n78062 & n78063;
  assign n78057 = n78066 & n78067;
  assign n78023 = ~n78031;
  assign n75451 = ~n75387;
  assign n78042 = n78050 & n78051;
  assign n78043 = n78050 & n78054;
  assign n75545 = n78055 & n78056;
  assign n78037 = n78057 ^ n78058;
  assign n78044 = ~n78057;
  assign n78032 = n35 ^ n78037;
  assign n77918 = n77948 ^ n75545;
  assign n78018 = ~n78042;
  assign n75613 = ~n75545;
  assign n78035 = ~n78043;
  assign n78041 = n78044 & n78045;
  assign n77926 = n78031 ^ n78032;
  assign n78030 = n77918 & n47;
  assign n78026 = ~n77918;
  assign n78022 = ~n78032;
  assign n78033 = n78035 & n78036;
  assign n78027 = n75613 & n78040;
  assign n78038 = ~n78041;
  assign n77933 = ~n77926;
  assign n77989 = n78022 & n78023;
  assign n78021 = n78026 & n12057;
  assign n77876 = n78027 ^ n75466;
  assign n77901 = ~n78030;
  assign n78020 = n78027 & n75466;
  assign n78015 = n78033 & n78034;
  assign n78024 = n78038 & n78039;
  assign n75225 = n78015 ^ n78016;
  assign n78011 = n77876 & n46;
  assign n77994 = ~n77989;
  assign n78013 = n78020 & n75451;
  assign n78012 = ~n77876;
  assign n77923 = ~n78021;
  assign n78010 = n78024 ^ n78025;
  assign n78017 = ~n78015;
  assign n78014 = ~n78020;
  assign n78028 = ~n78024;
  assign n78006 = n75225 & n77230;
  assign n77990 = n34 ^ n78010;
  assign n75275 = ~n75225;
  assign n77863 = ~n78011;
  assign n78007 = n78012 & n12021;
  assign n78005 = ~n78013;
  assign n77987 = n78014 & n75387;
  assign n78003 = n78017 & n78016;
  assign n75303 = n78017 & n78018;
  assign n78019 = n78028 & n78029;
  assign n77975 = n77987 ^ n75275;
  assign n77090 = n77989 ^ n77990;
  assign n77988 = n75275 & n77999;
  assign n75163 = n78003 ^ n78004;
  assign n77983 = n77987 & n75275;
  assign n77228 = ~n78006;
  assign n77822 = n44 ^ n77987;
  assign n78000 = n77987 & n44;
  assign n77884 = ~n78007;
  assign n77993 = ~n77990;
  assign n77998 = ~n77987;
  assign n78001 = ~n78003;
  assign n75357 = ~n75303;
  assign n78008 = ~n78019;
  assign n77971 = n77975 & n11895;
  assign n77749 = n77983 ^ n75163;
  assign n77981 = n75163 & n77207;
  assign n77912 = ~n77090;
  assign n77786 = ~n77975;
  assign n77215 = ~n77988;
  assign n75215 = ~n75163;
  assign n77982 = ~n77983;
  assign n77956 = n77993 & n77994;
  assign n77995 = n77998 & n11934;
  assign n77809 = ~n78000;
  assign n77976 = n78001 & n78002;
  assign n77986 = n77998 & n78005;
  assign n77991 = n78008 & n78009;
  assign n77963 = n77749 & n42;
  assign n77784 = ~n77971;
  assign n77968 = n77786 & n43;
  assign n77966 = ~n77749;
  assign n75140 = n77976 ^ n77977;
  assign n77970 = n75215 & n77980;
  assign n77204 = ~n77981;
  assign n77967 = n75215 & n77982;
  assign n77952 = ~n77956;
  assign n77984 = n77986 & n11976;
  assign n77848 = ~n77986;
  assign n77978 = ~n77976;
  assign n77974 = n77991 ^ n77992;
  assign n77820 = ~n77995;
  assign n77996 = ~n77991;
  assign n77728 = ~n77963;
  assign n77950 = n77966 & n11867;
  assign n77962 = n75140 & n77165;
  assign n77768 = ~n77968;
  assign n77960 = ~n77967;
  assign n75154 = ~n75140;
  assign n77193 = ~n77970;
  assign n77957 = n33 ^ n77974;
  assign n77964 = n77978 & n77979;
  assign n77969 = n77848 & n45;
  assign n77846 = ~n77984;
  assign n77985 = n77996 & n77997;
  assign n77747 = ~n77950;
  assign n77085 = n77956 ^ n77957;
  assign n77701 = n77960 & n75140;
  assign n77955 = n75154 & n77961;
  assign n77168 = ~n77962;
  assign n75046 = n77964 ^ n77965;
  assign n77949 = n77967 & n75154;
  assign n77951 = ~n77957;
  assign n77833 = ~n77969;
  assign n77958 = ~n77964;
  assign n77972 = ~n77985;
  assign n77941 = n77701 & n40;
  assign n77897 = ~n77085;
  assign n77939 = n75046 & n77946;
  assign n75078 = ~n75046;
  assign n77940 = ~n77949;
  assign n77920 = n77951 & n77952;
  assign n77932 = ~n77701;
  assign n77178 = ~n77955;
  assign n77942 = n77958 & n77959;
  assign n77947 = n77972 & n77973;
  assign n77157 = ~n77939;
  assign n77937 = n77932 & n11752;
  assign n77929 = n77932 & n77940;
  assign n77693 = ~n77941;
  assign n77938 = n75078 & n77159;
  assign n74986 = n77942 ^ n77943;
  assign n77930 = n77942 & n77945;
  assign n77916 = ~n77920;
  assign n77934 = n77947 ^ n77948;
  assign n77953 = ~n77947;
  assign n77687 = n77701 ^ n74986;
  assign n77924 = n77929 & n11822;
  assign n74963 = n77930 ^ n77931;
  assign n77911 = n74986 & n77932;
  assign n77925 = n74986 & n77933;
  assign n77921 = n32 ^ n77934;
  assign n75050 = ~n74986;
  assign n77720 = ~n77929;
  assign n77697 = ~n77937;
  assign n77149 = ~n77938;
  assign n77927 = ~n77930;
  assign n77944 = n77953 & n77954;
  assign n77904 = n77687 & n11714;
  assign n77669 = n77911 ^ n74963;
  assign n77909 = n74963 & n77090;
  assign n77905 = ~n77687;
  assign n77039 = n77920 ^ n77921;
  assign n75009 = ~n74963;
  assign n77914 = n77720 & n41;
  assign n77718 = ~n77924;
  assign n77910 = ~n77911;
  assign n77118 = ~n77925;
  assign n77919 = n75050 & n77926;
  assign n77906 = n77927 & n77928;
  assign n77915 = ~n77921;
  assign n77935 = ~n77944;
  assign n77894 = n77669 & n54;
  assign n77890 = ~n77669;
  assign n77685 = ~n77904;
  assign n77899 = n77905 & n55;
  assign n74899 = n77906 ^ n77907;
  assign n77093 = ~n77909;
  assign n77889 = n77910 & n74963;
  assign n77903 = n75009 & n77912;
  assign n77870 = ~n77039;
  assign n77709 = ~n77914;
  assign n77877 = n77915 & n77916;
  assign n77136 = ~n77919;
  assign n77908 = ~n77906;
  assign n77917 = n77935 & n77936;
  assign n77886 = n77890 & n11658;
  assign n77664 = ~n77894;
  assign n77893 = n74899 & n77897;
  assign n77678 = ~n77899;
  assign n74956 = ~n74899;
  assign n77895 = ~n77889;
  assign n77108 = ~n77903;
  assign n77898 = n77118 & n77136;
  assign n77885 = ~n77877;
  assign n77891 = n77908 & n77907;
  assign n77896 = n77917 ^ n77918;
  assign n77922 = ~n77917;
  assign n77674 = ~n77886;
  assign n77887 = n74956 & n77085;
  assign n77888 = n77889 & n74956;
  assign n74857 = n77891 ^ n77892;
  assign n77069 = ~n77893;
  assign n77858 = n77895 & n74899;
  assign n77878 = n47 ^ n77896;
  assign n77132 = ~n77898;
  assign n77881 = n77891 & n77902;
  assign n77913 = n77922 & n77923;
  assign n77639 = n52 ^ n77858;
  assign n77874 = n74857 & n77039;
  assign n77006 = n77877 ^ n77878;
  assign n74838 = n77881 ^ n77882;
  assign n77872 = n77858 & n11500;
  assign n74916 = ~n74857;
  assign n77841 = n77878 & n77885;
  assign n77082 = ~n77887;
  assign n77869 = ~n77858;
  assign n77873 = ~n77888;
  assign n77879 = ~n77881;
  assign n77900 = ~n77913;
  assign n77631 = n77858 ^ n74838;
  assign n77860 = n74838 & n77006;
  assign n77831 = n77869 & n74838;
  assign n77861 = ~n77006;
  assign n77867 = n74916 & n77870;
  assign n77654 = ~n77872;
  assign n77868 = n77869 & n52;
  assign n77859 = n77869 & n77873;
  assign n74846 = ~n74838;
  assign n77036 = ~n77874;
  assign n77865 = n77879 & n77880;
  assign n77875 = n77900 & n77901;
  assign n77844 = n77631 & n51;
  assign n77843 = ~n77631;
  assign n77855 = n77859 & n53;
  assign n77001 = ~n77860;
  assign n77856 = n74846 & n77861;
  assign n77850 = n77865 ^ n77866;
  assign n77062 = ~n77867;
  assign n77852 = n77865 & n77866;
  assign n77644 = ~n77868;
  assign n77857 = ~n77859;
  assign n77864 = n77875 ^ n77876;
  assign n77883 = ~n77875;
  assign n77840 = n77843 & n11429;
  assign n77626 = ~n77844;
  assign n74769 = n77849 ^ n77850;
  assign n74729 = n77852 ^ n77853;
  assign n77637 = ~n77855;
  assign n77021 = ~n77856;
  assign n77851 = n77857 & n11582;
  assign n77842 = n46 ^ n77864;
  assign n77854 = ~n77852;
  assign n77871 = n77883 & n77884;
  assign n77618 = n77831 ^ n74769;
  assign n74833 = ~n74769;
  assign n77629 = ~n77840;
  assign n76974 = n77841 ^ n77842;
  assign n74794 = ~n74729;
  assign n77660 = ~n77851;
  assign n77836 = n77854 & n77853;
  assign n77814 = n77842 & n77841;
  assign n77862 = ~n77871;
  assign n77825 = n77618 & n50;
  assign n77823 = ~n77618;
  assign n77826 = n77831 & n74833;
  assign n74688 = n77836 ^ n77837;
  assign n77835 = n74769 & n76974;
  assign n77828 = n77836 & n77837;
  assign n77834 = ~n76974;
  assign n77838 = n77660 & n77637;
  assign n77847 = n77862 & n77863;
  assign n77813 = n77823 & n11352;
  assign n77612 = ~n77825;
  assign n77824 = n77826 & n74794;
  assign n74649 = n77828 ^ n77829;
  assign n77816 = ~n77826;
  assign n77827 = n74833 & n77834;
  assign n77817 = n77828 & n77829;
  assign n74731 = ~n74688;
  assign n76992 = ~n77835;
  assign n77658 = ~n77838;
  assign n77830 = n77847 ^ n77848;
  assign n77845 = ~n77847;
  assign n77623 = ~n77813;
  assign n77800 = n77816 & n74729;
  assign n74606 = n77817 ^ n77818;
  assign n77799 = ~n77824;
  assign n74712 = ~n74649;
  assign n77810 = n77817 & n77818;
  assign n76972 = ~n77827;
  assign n77815 = n45 ^ n77830;
  assign n77839 = n77845 & n77846;
  assign n77583 = n48 ^ n77800;
  assign n77793 = n77800 ^ n74712;
  assign n77791 = n74712 & n77800;
  assign n74571 = n77810 ^ n77811;
  assign n77807 = n77800 & n11173;
  assign n74657 = ~n74606;
  assign n77798 = ~n77800;
  assign n77795 = n77810 & n77811;
  assign n76956 = n77814 ^ n77815;
  assign n77805 = n77815 & n77814;
  assign n77832 = ~n77839;
  assign n77773 = n77791 ^ n74657;
  assign n77777 = n77793 & n63;
  assign n77778 = ~n77793;
  assign n77772 = n77791 & n74657;
  assign n74529 = n77795 ^ n77796;
  assign n77792 = n77798 & n77799;
  assign n74618 = ~n74571;
  assign n77794 = n77798 & n48;
  assign n77787 = n77795 & n77796;
  assign n77601 = ~n77807;
  assign n77801 = n76956 & n74794;
  assign n77802 = ~n76956;
  assign n77804 = ~n77805;
  assign n77821 = n77832 & n77833;
  assign n77760 = n77772 ^ n74618;
  assign n77769 = n77773 & n62;
  assign n77545 = ~n77777;
  assign n77771 = n77778 & n11134;
  assign n77770 = ~n77773;
  assign n74474 = n77787 ^ n77788;
  assign n77757 = n74618 & n77772;
  assign n77789 = n77792 & n49;
  assign n74577 = ~n74529;
  assign n77586 = ~n77794;
  assign n77780 = ~n77792;
  assign n77781 = ~n77787;
  assign n76960 = ~n77801;
  assign n77797 = n77802 & n74729;
  assign n77806 = n77821 ^ n77822;
  assign n77819 = ~n77821;
  assign n77753 = n77760 & n61;
  assign n77756 = ~n77760;
  assign n77511 = ~n77769;
  assign n77761 = n77770 & n10999;
  assign n77759 = n77757 & n10873;
  assign n77569 = ~n77771;
  assign n74510 = ~n74474;
  assign n77758 = ~n77757;
  assign n77776 = n77780 & n11263;
  assign n77765 = n77781 & n77782;
  assign n77576 = ~n77789;
  assign n76933 = ~n77797;
  assign n76919 = n77805 ^ n77806;
  assign n77803 = ~n77806;
  assign n77812 = n77819 & n77820;
  assign n77459 = ~n77753;
  assign n77751 = n77756 & n10917;
  assign n77741 = n77757 ^ n74510;
  assign n77738 = n77758 & n74474;
  assign n77558 = ~n77759;
  assign n77529 = ~n77761;
  assign n77754 = n77569 & n77545;
  assign n77755 = n77758 & n60;
  assign n74421 = n77765 ^ n77766;
  assign n77763 = ~n77765;
  assign n77606 = ~n77776;
  assign n77779 = n76919 & n74731;
  assign n77790 = ~n76919;
  assign n77742 = n77803 & n77804;
  assign n77808 = ~n77812;
  assign n77408 = n77738 ^ n74421;
  assign n77737 = n77741 & n10788;
  assign n77440 = ~n77741;
  assign n77744 = n77529 & n77511;
  assign n77491 = ~n77751;
  assign n77567 = ~n77754;
  assign n74488 = ~n74421;
  assign n77474 = ~n77755;
  assign n77745 = ~n77738;
  assign n77752 = n77606 & n77576;
  assign n77739 = n77763 & n77764;
  assign n76890 = ~n77779;
  assign n77775 = n77790 & n74688;
  assign n77750 = ~n77742;
  assign n77785 = n77808 & n77809;
  assign n77729 = n77408 & n58;
  assign n77723 = ~n77408;
  assign n77733 = n77440 & n59;
  assign n77734 = n77491 & n77459;
  assign n77444 = ~n77737;
  assign n74379 = n77739 ^ n77740;
  assign n77542 = ~n77744;
  assign n77724 = n74488 & n77745;
  assign n77735 = n77474 & n77558;
  assign n77731 = n77739 & n77740;
  assign n77608 = ~n77752;
  assign n76915 = ~n77775;
  assign n77762 = n77785 ^ n77786;
  assign n77783 = ~n77785;
  assign n77722 = n77723 & n10703;
  assign n77370 = n77724 ^ n74379;
  assign n77386 = ~n77729;
  assign n74423 = n77731 ^ n77732;
  assign n77422 = ~n77733;
  assign n77507 = ~n77734;
  assign n74448 = ~n74379;
  assign n77470 = ~n77735;
  assign n77743 = n43 ^ n77762;
  assign n77774 = n77783 & n77784;
  assign n77712 = n77370 & n10623;
  assign n77713 = ~n77370;
  assign n77399 = ~n77722;
  assign n77714 = n74448 & n77724;
  assign n76830 = n77742 ^ n77743;
  assign n77715 = n77743 & n77750;
  assign n77767 = ~n77774;
  assign n77372 = ~n77712;
  assign n77711 = n77713 & n57;
  assign n77334 = n56 ^ n77714;
  assign n77725 = n76830 & n74712;
  assign n77726 = ~n76830;
  assign n77748 = n77767 & n77768;
  assign n77351 = ~n77711;
  assign n76835 = ~n77725;
  assign n77721 = n77726 & n74649;
  assign n77730 = n77748 ^ n77749;
  assign n77746 = ~n77748;
  assign n76858 = ~n77721;
  assign n77716 = n42 ^ n77730;
  assign n77736 = n77746 & n77747;
  assign n76808 = n77715 ^ n77716;
  assign n77702 = n77716 & n77715;
  assign n77727 = ~n77736;
  assign n77705 = n76808 & n74606;
  assign n77707 = ~n76808;
  assign n77699 = ~n77702;
  assign n77719 = n77727 & n77728;
  assign n76805 = ~n77705;
  assign n77704 = n77707 & n74657;
  assign n77706 = n77719 ^ n77720;
  assign n77717 = ~n77719;
  assign n76784 = ~n77704;
  assign n77703 = n41 ^ n77706;
  assign n77710 = n77717 & n77718;
  assign n76753 = n77702 ^ n77703;
  assign n77698 = ~n77703;
  assign n77708 = ~n77710;
  assign n77690 = n76753 & n74618;
  assign n77694 = ~n76753;
  assign n77682 = n77698 & n77699;
  assign n77700 = n77708 & n77709;
  assign n76729 = ~n77690;
  assign n77689 = n77694 & n74571;
  assign n77688 = ~n77682;
  assign n77691 = n77700 ^ n77701;
  assign n77696 = ~n77700;
  assign n76748 = ~n77689;
  assign n77683 = n40 ^ n77691;
  assign n77695 = n77696 & n77697;
  assign n76702 = n77682 ^ n77683;
  assign n77671 = n77683 & n77688;
  assign n77692 = ~n77695;
  assign n77679 = n76702 & n74577;
  assign n77680 = ~n76702;
  assign n77686 = n77692 & n77693;
  assign n76669 = ~n77679;
  assign n77675 = n77680 & n74529;
  assign n77676 = n77686 ^ n77687;
  assign n77684 = ~n77686;
  assign n76698 = ~n77675;
  assign n77672 = n55 ^ n77676;
  assign n77681 = n77684 & n77685;
  assign n76618 = n77671 ^ n77672;
  assign n77670 = ~n77672;
  assign n77677 = ~n77681;
  assign n77665 = n76618 & n74474;
  assign n77662 = ~n76618;
  assign n77655 = n77670 & n77671;
  assign n77668 = n77677 & n77678;
  assign n77661 = n77662 & n74510;
  assign n76612 = ~n77665;
  assign n77666 = n77668 ^ n77669;
  assign n77673 = ~n77668;
  assign n76638 = ~n77661;
  assign n77656 = n54 ^ n77666;
  assign n77667 = n77673 & n77674;
  assign n76584 = n77655 ^ n77656;
  assign n77646 = n77656 & n77655;
  assign n77663 = ~n77667;
  assign n77652 = n76584 & n74421;
  assign n77648 = ~n76584;
  assign n77657 = n77663 & n77664;
  assign n77645 = n77648 & n74488;
  assign n76588 = ~n77652;
  assign n77647 = n77657 ^ n77658;
  assign n77659 = ~n77657;
  assign n76563 = ~n77645;
  assign n76531 = n77646 ^ n77647;
  assign n77650 = ~n77647;
  assign n77653 = n77659 & n77660;
  assign n77641 = n76531 & n74448;
  assign n77642 = ~n76531;
  assign n77640 = n77650 & n77646;
  assign n77651 = n77653 & n77654;
  assign n77649 = ~n77653;
  assign n77633 = n77640 ^ n74423;
  assign n76497 = ~n77641;
  assign n77635 = n77642 & n74379;
  assign n77634 = ~n77640;
  assign n77638 = n77649 & n77637;
  assign n77643 = ~n77651;
  assign n76523 = ~n77635;
  assign n77632 = n77638 ^ n77639;
  assign n77636 = n77643 & n77644;
  assign n76470 = n77632 ^ n77633;
  assign n77619 = n77632 & n77634;
  assign n77630 = n77636 & n77637;
  assign n77624 = n77630 ^ n77631;
  assign n77628 = ~n77630;
  assign n77620 = n51 ^ n77624;
  assign n77627 = n77628 & n77629;
  assign n77614 = n77619 ^ n77620;
  assign n77621 = ~n77620;
  assign n77625 = ~n77627;
  assign n74445 = n76199 ^ n77614;
  assign n77613 = ~n77614;
  assign n77602 = n77621 & n77619;
  assign n77617 = n77625 & n77626;
  assign n77564 = n77613 & n76204;
  assign n77609 = n77613 & n76199;
  assign n77615 = n77617 ^ n77618;
  assign n77622 = ~n77617;
  assign n76193 = n71 ^ n77609;
  assign n77610 = ~n77609;
  assign n77603 = n50 ^ n77615;
  assign n77616 = n77622 & n77623;
  assign n77086 = ~n76193;
  assign n77599 = n77602 ^ n77603;
  assign n77543 = n77610 & n71;
  assign n77604 = ~n77603;
  assign n77611 = ~n77616;
  assign n77598 = n77599 & n76115;
  assign n77591 = n77543 & n70;
  assign n77589 = ~n77543;
  assign n77595 = ~n77599;
  assign n77596 = n77604 & n77602;
  assign n77607 = n77611 & n77612;
  assign n77588 = n77589 & n3685;
  assign n77524 = ~n77591;
  assign n77587 = n77595 & n76103;
  assign n77579 = ~n77598;
  assign n77594 = ~n77596;
  assign n77597 = n77607 ^ n77608;
  assign n77605 = ~n77607;
  assign n77581 = n77579 & n77564;
  assign n77574 = ~n77587;
  assign n77540 = ~n77588;
  assign n77548 = n77596 ^ n77597;
  assign n77593 = ~n77597;
  assign n77600 = n77605 & n77606;
  assign n77577 = n77579 & n77574;
  assign n77573 = ~n77581;
  assign n77584 = n77548 & n76009;
  assign n77580 = ~n77548;
  assign n77571 = n77593 & n77594;
  assign n77590 = n77600 & n77601;
  assign n77592 = ~n77600;
  assign n77561 = n77573 & n77574;
  assign n77565 = ~n77577;
  assign n77578 = n77580 & n76085;
  assign n77562 = ~n77584;
  assign n77585 = ~n77590;
  assign n77582 = n77592 & n77576;
  assign n77549 = n77561 ^ n76009;
  assign n74366 = n77564 ^ n77565;
  assign n77563 = ~n77561;
  assign n77547 = ~n77578;
  assign n77572 = n77582 ^ n77583;
  assign n77575 = n77585 & n77586;
  assign n74305 = n77548 ^ n77549;
  assign n74359 = ~n74366;
  assign n77560 = n77562 & n77563;
  assign n77512 = n77571 ^ n77572;
  assign n77566 = n77575 & n77576;
  assign n77570 = ~n77572;
  assign n74325 = ~n74305;
  assign n77517 = n74359 & n76103;
  assign n77546 = ~n77560;
  assign n77559 = n77512 & n75948;
  assign n77552 = n77566 ^ n77567;
  assign n77556 = ~n77512;
  assign n77551 = n77570 & n77571;
  assign n77568 = ~n77566;
  assign n77516 = n74325 & n76085;
  assign n77526 = n77543 ^ n77517;
  assign n77515 = ~n77517;
  assign n77534 = n77546 & n77547;
  assign n77500 = n77551 ^ n77552;
  assign n77550 = n77556 & n76006;
  assign n77519 = ~n77559;
  assign n77555 = ~n77551;
  assign n77557 = n77568 & n77569;
  assign n77493 = n77516 ^ n77517;
  assign n77503 = n70 ^ n77526;
  assign n77514 = ~n77516;
  assign n77513 = n77534 ^ n75948;
  assign n77533 = n77515 & n77540;
  assign n77532 = ~n77534;
  assign n77539 = n77500 & n75942;
  assign n77538 = ~n77500;
  assign n77531 = ~n77550;
  assign n77521 = n77552 & n77555;
  assign n77554 = n77557 & n77558;
  assign n77553 = ~n77557;
  assign n76127 = n77503 ^ n76193;
  assign n77460 = n77503 & n76193;
  assign n77488 = ~n77493;
  assign n74270 = n77512 ^ n77513;
  assign n77478 = n77514 & n77515;
  assign n77527 = n77531 & n77532;
  assign n77523 = ~n77533;
  assign n77530 = n77538 & n75861;
  assign n77496 = ~n77539;
  assign n77541 = n77553 & n77545;
  assign n77544 = ~n77554;
  assign n77051 = ~n76127;
  assign n77467 = ~n77460;
  assign n74288 = ~n74270;
  assign n77492 = n77523 & n77524;
  assign n77518 = ~n77527;
  assign n77481 = ~n77530;
  assign n77522 = n77541 ^ n77542;
  assign n77537 = n77544 & n77545;
  assign n77536 = ~n77541;
  assign n77479 = n74288 & n76006;
  assign n77475 = n77492 ^ n77493;
  assign n77508 = n77492 & n3604;
  assign n77509 = ~n77492;
  assign n77499 = n77518 & n77519;
  assign n77435 = n77521 ^ n77522;
  assign n77484 = n77522 & n77521;
  assign n77535 = n77536 & n77529;
  assign n77528 = ~n77537;
  assign n77461 = n69 ^ n77475;
  assign n77453 = n77478 ^ n77479;
  assign n77455 = n77479 & n77478;
  assign n77476 = n77499 ^ n77500;
  assign n77489 = ~n77508;
  assign n77497 = n77509 & n69;
  assign n77501 = n77435 & n75834;
  assign n77495 = ~n77499;
  assign n77502 = ~n77435;
  assign n77520 = n77528 & n77529;
  assign n77525 = ~n77535;
  assign n76072 = n77460 ^ n77461;
  assign n77417 = n77461 & n77467;
  assign n77438 = ~n77453;
  assign n74247 = n77476 ^ n75942;
  assign n77477 = ~n77476;
  assign n77483 = n77488 & n77489;
  assign n77487 = n77495 & n77496;
  assign n77472 = ~n77497;
  assign n77442 = ~n77501;
  assign n77498 = n77502 & n75836;
  assign n77510 = ~n77520;
  assign n77506 = n77525 & n77511;
  assign n77024 = ~n76072;
  assign n77420 = ~n77417;
  assign n74236 = ~n74247;
  assign n77456 = n77477 & n75861;
  assign n77471 = ~n77483;
  assign n77480 = ~n77487;
  assign n77463 = ~n77498;
  assign n77485 = n77506 ^ n77507;
  assign n77504 = n77510 & n77511;
  assign n77505 = ~n77506;
  assign n77392 = n77455 ^ n77456;
  assign n77465 = ~n77456;
  assign n77452 = n77471 & n77472;
  assign n77464 = n77480 & n77481;
  assign n77411 = n77484 ^ n77485;
  assign n77448 = n77485 & n77484;
  assign n77490 = ~n77504;
  assign n77494 = n77505 & n77491;
  assign n77433 = n77452 ^ n77453;
  assign n77450 = n77452 & n3531;
  assign n77436 = n77464 ^ n75836;
  assign n77414 = n77465 & n77455;
  assign n77451 = ~n77452;
  assign n77468 = n77411 & n75703;
  assign n77462 = ~n77464;
  assign n77466 = ~n77411;
  assign n77447 = ~n77448;
  assign n77482 = n77490 & n77491;
  assign n77486 = ~n77494;
  assign n77418 = n68 ^ n77433;
  assign n74193 = n77435 ^ n77436;
  assign n77437 = ~n77450;
  assign n77445 = n77451 & n68;
  assign n77454 = n77462 & n77463;
  assign n77457 = n77466 & n75757;
  assign n77410 = ~n77468;
  assign n77473 = ~n77482;
  assign n77469 = n77486 & n77459;
  assign n76022 = n77417 ^ n77418;
  assign n77415 = n74193 & n75834;
  assign n77419 = ~n77418;
  assign n74202 = ~n74193;
  assign n77434 = n77437 & n77438;
  assign n77425 = ~n77445;
  assign n77441 = ~n77454;
  assign n77427 = ~n77457;
  assign n77449 = n77469 ^ n77470;
  assign n77458 = n77473 & n77474;
  assign n76988 = ~n76022;
  assign n77359 = n77414 ^ n77415;
  assign n77361 = n77419 & n77420;
  assign n77413 = ~n77415;
  assign n77424 = ~n77434;
  assign n77429 = n77441 & n77442;
  assign n77383 = n77448 ^ n77449;
  assign n77439 = n77458 & n77459;
  assign n77446 = ~n77449;
  assign n77393 = n77359 & n66;
  assign n77395 = ~n77359;
  assign n77363 = n77413 & n77414;
  assign n77401 = n77424 & n77425;
  assign n77412 = n77429 ^ n75703;
  assign n77426 = ~n77429;
  assign n77431 = n77383 & n75683;
  assign n77430 = ~n77383;
  assign n77423 = n77439 ^ n77440;
  assign n77404 = n77446 & n77447;
  assign n77443 = ~n77439;
  assign n77338 = ~n77393;
  assign n77387 = n77395 & n3384;
  assign n77391 = n67 ^ n77401;
  assign n74151 = n77411 ^ n77412;
  assign n77400 = n77401 & n3431;
  assign n77406 = ~n77401;
  assign n77405 = n59 ^ n77423;
  assign n77416 = n77426 & n77427;
  assign n77428 = n77430 & n75627;
  assign n77390 = ~n77431;
  assign n77403 = ~n77404;
  assign n77432 = n77443 & n77444;
  assign n77356 = ~n77387;
  assign n77362 = n77391 ^ n77392;
  assign n74158 = ~n74151;
  assign n77394 = ~n77400;
  assign n77344 = n77404 ^ n77405;
  assign n77397 = n77406 & n67;
  assign n77409 = ~n77416;
  assign n77402 = ~n77405;
  assign n77366 = ~n77428;
  assign n77421 = ~n77432;
  assign n75958 = n77361 ^ n77362;
  assign n77316 = n77362 & n77361;
  assign n77364 = n74158 & n75703;
  assign n77384 = n77394 & n77392;
  assign n77381 = n77344 & n75613;
  assign n77388 = ~n77344;
  assign n77377 = ~n77397;
  assign n77373 = n77402 & n77403;
  assign n77382 = n77409 & n77410;
  assign n77407 = n77421 & n77422;
  assign n76957 = ~n75958;
  assign n77321 = n77363 ^ n77364;
  assign n77323 = ~n77316;
  assign n77368 = ~n77364;
  assign n77327 = ~n77381;
  assign n77367 = n77382 ^ n77383;
  assign n77376 = ~n77384;
  assign n77379 = n77388 & n75545;
  assign n77375 = ~n77373;
  assign n77389 = ~n77382;
  assign n77380 = n77407 ^ n77408;
  assign n77398 = ~n77407;
  assign n77353 = n77321 & n65;
  assign n77345 = ~n77321;
  assign n74118 = n77367 ^ n75683;
  assign n77348 = n77368 & n77363;
  assign n77349 = n77367 & n75683;
  assign n77358 = n77376 & n77377;
  assign n77355 = ~n77379;
  assign n77374 = n58 ^ n77380;
  assign n77378 = n77389 & n77390;
  assign n77396 = n77398 & n77399;
  assign n77341 = n77345 & n3342;
  assign n77287 = n77348 ^ n77349;
  assign n77300 = ~n77353;
  assign n77309 = n77349 & n77348;
  assign n77336 = n77358 ^ n77359;
  assign n74103 = ~n74118;
  assign n77357 = ~n77358;
  assign n77296 = n77373 ^ n77374;
  assign n77329 = n77374 & n77375;
  assign n77365 = ~n77378;
  assign n77385 = ~n77396;
  assign n77317 = n66 ^ n77336;
  assign n77325 = n77287 & n3315;
  assign n77332 = ~n77287;
  assign n77318 = ~n77341;
  assign n77313 = ~n77309;
  assign n77342 = n77296 & n75466;
  assign n77347 = n77356 & n77357;
  assign n77352 = ~n77296;
  assign n77343 = n77365 & n77366;
  assign n77369 = n77385 & n77386;
  assign n75892 = n77316 ^ n77317;
  assign n77283 = ~n77325;
  assign n77322 = ~n77317;
  assign n77324 = n77332 & n64;
  assign n77295 = ~n77342;
  assign n77335 = n77343 ^ n77344;
  assign n77337 = ~n77347;
  assign n77340 = n77352 & n75525;
  assign n77354 = ~n77343;
  assign n77346 = n77369 ^ n77370;
  assign n77371 = ~n77369;
  assign n76922 = ~n75892;
  assign n77284 = n77322 & n77323;
  assign n77276 = ~n77324;
  assign n74096 = n77335 ^ n75613;
  assign n77320 = n77337 & n77338;
  assign n77308 = ~n77340;
  assign n77330 = ~n77335;
  assign n77331 = n57 ^ n77346;
  assign n77339 = n77354 & n77355;
  assign n77360 = n77371 & n77372;
  assign n77288 = ~n77284;
  assign n77301 = n77320 ^ n77321;
  assign n74067 = ~n74096;
  assign n77310 = n77330 & n75545;
  assign n77271 = n77329 ^ n77331;
  assign n77319 = ~n77320;
  assign n77326 = ~n77339;
  assign n77328 = ~n77331;
  assign n77350 = ~n77360;
  assign n77285 = n65 ^ n77301;
  assign n77251 = n77309 ^ n77310;
  assign n77311 = n77271 & n75387;
  assign n77314 = n77318 & n77319;
  assign n77312 = ~n77310;
  assign n77315 = ~n77271;
  assign n77306 = n77326 & n77327;
  assign n77304 = n77328 & n77329;
  assign n77333 = n77350 & n77351;
  assign n75819 = n77284 ^ n77285;
  assign n77262 = n77285 & n77288;
  assign n77293 = n77251 & n79;
  assign n77298 = ~n77251;
  assign n77297 = n77306 ^ n75466;
  assign n77270 = ~n77311;
  assign n77268 = n77312 & n77313;
  assign n77299 = ~n77314;
  assign n77303 = n77315 & n75451;
  assign n77307 = ~n77306;
  assign n77305 = n77333 ^ n77334;
  assign n76865 = ~n75819;
  assign n77249 = ~n77293;
  assign n74024 = n77296 ^ n77297;
  assign n77289 = n77298 & n3280;
  assign n77286 = n77299 & n77300;
  assign n77279 = ~n77303;
  assign n77259 = n77304 ^ n77305;
  assign n77302 = n77307 & n77308;
  assign n77274 = n77286 ^ n77287;
  assign n77265 = ~n77289;
  assign n74051 = ~n74024;
  assign n77282 = ~n77286;
  assign n77291 = n77259 & n75357;
  assign n77294 = ~n77302;
  assign n77292 = ~n77259;
  assign n77263 = n64 ^ n77274;
  assign n77273 = n74051 & n75525;
  assign n77280 = n77282 & n77283;
  assign n77241 = ~n77291;
  assign n77290 = n77292 & n75303;
  assign n77281 = n77294 & n77295;
  assign n76818 = n77262 ^ n77263;
  assign n77233 = n77268 ^ n77273;
  assign n77261 = ~n77263;
  assign n77267 = ~n77273;
  assign n77275 = ~n77280;
  assign n77272 = n77281 ^ n75387;
  assign n77278 = ~n77281;
  assign n77255 = ~n77290;
  assign n76806 = ~n76818;
  assign n77257 = n77233 & n3229;
  assign n77236 = n77261 & n77262;
  assign n77256 = ~n77233;
  assign n77246 = n77267 & n77268;
  assign n73988 = n77271 ^ n77272;
  assign n77266 = n77275 & n77276;
  assign n77277 = n77278 & n77279;
  assign n77252 = n77256 & n78;
  assign n77239 = ~n77257;
  assign n77235 = ~n77236;
  assign n77250 = n79 ^ n77266;
  assign n73990 = ~n73988;
  assign n77243 = ~n77246;
  assign n77264 = ~n77266;
  assign n77269 = ~n77277;
  assign n77237 = n77250 ^ n77251;
  assign n77220 = ~n77252;
  assign n77247 = n73990 & n75387;
  assign n77260 = n77264 & n77265;
  assign n77258 = n77269 & n77270;
  assign n75717 = n77236 ^ n77237;
  assign n77213 = n77246 ^ n77247;
  assign n77234 = ~n77237;
  assign n77242 = ~n77247;
  assign n77244 = n77258 ^ n77259;
  assign n77248 = ~n77260;
  assign n77254 = ~n77258;
  assign n76771 = ~n75717;
  assign n77225 = n77213 & n3182;
  assign n77210 = n77234 & n77235;
  assign n77226 = ~n77213;
  assign n77223 = n77242 & n77243;
  assign n73985 = n77244 ^ n75357;
  assign n77232 = n77248 & n77249;
  assign n77245 = ~n77244;
  assign n77253 = n77254 & n77255;
  assign n77209 = ~n77225;
  assign n77222 = n77226 & n77;
  assign n77218 = n77232 ^ n77233;
  assign n73936 = ~n73985;
  assign n77238 = ~n77232;
  assign n77224 = n77245 & n75303;
  assign n77240 = ~n77253;
  assign n77211 = n78 ^ n77218;
  assign n77197 = ~n77222;
  assign n77187 = n77223 ^ n77224;
  assign n77200 = n77224 & n77223;
  assign n77231 = n77238 & n77239;
  assign n77229 = n77240 & n77241;
  assign n75656 = n77210 ^ n77211;
  assign n77180 = n77211 & n77210;
  assign n77175 = ~n77187;
  assign n77216 = n77229 ^ n77230;
  assign n77219 = ~n77231;
  assign n77227 = ~n77229;
  assign n76711 = ~n75656;
  assign n73898 = n77216 ^ n75225;
  assign n77212 = n77219 & n77220;
  assign n77217 = ~n77216;
  assign n77221 = n77227 & n77228;
  assign n77198 = n77212 ^ n77213;
  assign n73938 = ~n73898;
  assign n77208 = ~n77212;
  assign n77201 = n77217 & n75275;
  assign n77214 = ~n77221;
  assign n77181 = n77 ^ n77198;
  assign n77155 = n77200 ^ n77201;
  assign n77205 = n77208 & n77209;
  assign n77202 = ~n77201;
  assign n77206 = n77214 & n77215;
  assign n75554 = n77180 ^ n77181;
  assign n77160 = n77181 & n77180;
  assign n77191 = n77155 & n75;
  assign n77195 = ~n77155;
  assign n77184 = n77202 & n77200;
  assign n77196 = ~n77205;
  assign n77194 = n77206 ^ n77207;
  assign n77203 = ~n77206;
  assign n76654 = ~n75554;
  assign n77141 = ~n77191;
  assign n73855 = n75163 ^ n77194;
  assign n77190 = n77195 & n3117;
  assign n77186 = n77196 & n77197;
  assign n77185 = n77194 & n75163;
  assign n77189 = ~n77184;
  assign n77199 = n77203 & n77204;
  assign n77127 = n77184 ^ n77185;
  assign n77170 = n77186 ^ n77187;
  assign n77182 = n77186 & n3147;
  assign n77153 = ~n77190;
  assign n73895 = ~n73855;
  assign n77183 = ~n77186;
  assign n77188 = ~n77185;
  assign n77192 = ~n77199;
  assign n77161 = n76 ^ n77170;
  assign n77172 = n77127 & n74;
  assign n77171 = ~n77127;
  assign n77174 = ~n77182;
  assign n77179 = n77183 & n76;
  assign n77142 = n77188 & n77189;
  assign n77176 = n77192 & n77193;
  assign n75515 = n77160 ^ n77161;
  assign n77128 = n77161 & n77160;
  assign n77164 = n77171 & n3056;
  assign n77114 = ~n77172;
  assign n77169 = n77174 & n77175;
  assign n77166 = n77176 ^ n75140;
  assign n77146 = ~n77142;
  assign n77163 = ~n77179;
  assign n77177 = ~n77176;
  assign n76598 = ~n75515;
  assign n77130 = ~n77128;
  assign n77123 = ~n77164;
  assign n73815 = n77165 ^ n77166;
  assign n77162 = ~n77169;
  assign n77173 = n77177 & n77178;
  assign n77154 = n77162 & n77163;
  assign n73810 = ~n73815;
  assign n77167 = ~n77173;
  assign n77139 = n77154 ^ n77155;
  assign n77143 = n73810 & n75140;
  assign n77152 = ~n77154;
  assign n77158 = n77167 & n77168;
  assign n77129 = n75 ^ n77139;
  assign n77100 = n77142 ^ n77143;
  assign n77145 = ~n77143;
  assign n77150 = n77152 & n77153;
  assign n77144 = n77158 ^ n77159;
  assign n77156 = ~n77158;
  assign n75398 = n77128 ^ n77129;
  assign n77101 = n77129 & n77130;
  assign n77138 = n77100 & n3021;
  assign n77137 = ~n77100;
  assign n73825 = n77144 ^ n75078;
  assign n77133 = n77145 & n77146;
  assign n77140 = ~n77150;
  assign n77147 = ~n77144;
  assign n77151 = n77156 & n77157;
  assign n76550 = ~n75398;
  assign n77124 = n77137 & n73;
  assign n77105 = ~n77138;
  assign n73761 = ~n73825;
  assign n77126 = n77140 & n77141;
  assign n77134 = n77147 & n75046;
  assign n77148 = ~n77151;
  assign n77089 = ~n77124;
  assign n77116 = n77126 ^ n77127;
  assign n77077 = n77133 ^ n77134;
  assign n77111 = n77134 & n77133;
  assign n77122 = ~n77126;
  assign n77131 = n77148 & n77149;
  assign n77102 = n74 ^ n77116;
  assign n77119 = n77077 & n2975;
  assign n77121 = n77122 & n77123;
  assign n77120 = ~n77077;
  assign n73701 = n77131 ^ n77132;
  assign n77110 = ~n77111;
  assign n77135 = ~n77131;
  assign n75339 = n77101 ^ n77102;
  assign n76443 = n77102 & n77101;
  assign n77075 = ~n77119;
  assign n77115 = n77120 & n72;
  assign n77113 = ~n77121;
  assign n77112 = n73701 & n75050;
  assign n73798 = ~n73701;
  assign n77125 = n77135 & n77136;
  assign n76468 = ~n75339;
  assign n77098 = n77111 ^ n77112;
  assign n77099 = n77113 & n77114;
  assign n77064 = ~n77115;
  assign n77109 = ~n77112;
  assign n77117 = ~n77125;
  assign n77095 = n77098 & n87;
  assign n77087 = n77099 ^ n77100;
  assign n77097 = ~n77098;
  assign n77104 = ~n77099;
  assign n77071 = n77109 & n77110;
  assign n77106 = n77117 & n77118;
  assign n76417 = n73 ^ n77087;
  assign n77033 = ~n77095;
  assign n77094 = n77097 & n2910;
  assign n77096 = n77104 & n77105;
  assign n77091 = n77106 ^ n74963;
  assign n77067 = ~n77071;
  assign n77107 = ~n77106;
  assign n77078 = ~n76417;
  assign n73663 = n77090 ^ n77091;
  assign n77050 = ~n77094;
  assign n77088 = ~n77096;
  assign n77103 = n77107 & n77108;
  assign n77043 = n77078 & n76443;
  assign n77083 = n73663 & n77086;
  assign n77045 = n77050 & n77033;
  assign n77076 = n77088 & n77089;
  assign n73744 = ~n73663;
  assign n77092 = ~n77103;
  assign n77057 = ~n77043;
  assign n77065 = n77076 ^ n77077;
  assign n76189 = ~n77083;
  assign n77079 = n73744 & n76193;
  assign n77072 = n73744 & n74963;
  assign n77074 = ~n77076;
  assign n77084 = n77092 & n77093;
  assign n77044 = n72 ^ n77065;
  assign n77012 = n77071 ^ n77072;
  assign n77073 = n77074 & n77075;
  assign n76168 = ~n77079;
  assign n77066 = ~n77072;
  assign n77070 = n77084 ^ n77085;
  assign n77081 = ~n77084;
  assign n77026 = n77043 ^ n77044;
  assign n77027 = n77044 & n77057;
  assign n77060 = n77012 & n2896;
  assign n77053 = ~n77012;
  assign n77055 = n77066 & n77067;
  assign n73648 = n77070 ^ n74956;
  assign n77063 = ~n77073;
  assign n77056 = n77070 & n74956;
  assign n77080 = n77081 & n77082;
  assign n73380 = n77026 ^ n74445;
  assign n77034 = n77026 & n74445;
  assign n77030 = ~n77026;
  assign n77042 = n77053 & n86;
  assign n76981 = n77055 ^ n77056;
  assign n77019 = ~n77060;
  assign n77054 = n73648 & n76127;
  assign n77046 = n77063 & n77064;
  assign n77059 = ~n77055;
  assign n73626 = ~n73648;
  assign n77058 = ~n77056;
  assign n77068 = ~n77080;
  assign n77014 = n73380 & n76204;
  assign n73382 = ~n73380;
  assign n76984 = n77030 & n74445;
  assign n77003 = ~n77034;
  assign n77038 = n76981 & n85;
  assign n76998 = ~n77042;
  assign n77037 = ~n76981;
  assign n77028 = n77045 ^ n77046;
  assign n77047 = n73626 & n77051;
  assign n76148 = ~n77054;
  assign n77005 = n77058 & n77059;
  assign n77049 = ~n77046;
  assign n77052 = n77068 & n77069;
  assign n77002 = ~n77014;
  assign n77023 = n77027 ^ n77028;
  assign n77029 = n77037 & n2826;
  assign n76965 = ~n77038;
  assign n77031 = ~n77028;
  assign n77009 = ~n77005;
  assign n76124 = ~n77047;
  assign n77041 = n77049 & n77050;
  assign n77040 = n77052 ^ n74857;
  assign n77061 = ~n77052;
  assign n76924 = n77002 & n77003;
  assign n77016 = n77023 & n74366;
  assign n77017 = ~n77023;
  assign n76979 = ~n77029;
  assign n76986 = n77031 & n77027;
  assign n73593 = n77039 ^ n77040;
  assign n77032 = ~n77041;
  assign n77048 = n77061 & n77062;
  assign n74872 = n103 ^ n76924;
  assign n76852 = n76924 & n103;
  assign n76928 = ~n76924;
  assign n76995 = ~n77016;
  assign n77008 = n77017 & n74359;
  assign n77022 = n73593 & n76072;
  assign n73660 = ~n73593;
  assign n77011 = n77032 & n77033;
  assign n77035 = ~n77048;
  assign n75865 = ~n74872;
  assign n76996 = n76995 & n76984;
  assign n76990 = ~n77008;
  assign n76999 = n77011 ^ n77012;
  assign n76098 = ~n77022;
  assign n77015 = n73660 & n77024;
  assign n77004 = n73660 & n74916;
  assign n77018 = ~n77011;
  assign n77025 = n77035 & n77036;
  assign n76983 = n76995 & n76990;
  assign n76989 = ~n76996;
  assign n76987 = n86 ^ n76999;
  assign n76938 = n77004 ^ n77005;
  assign n76969 = n77004 & n77009;
  assign n76064 = ~n77015;
  assign n77010 = n77018 & n77019;
  assign n77007 = n77025 ^ n74838;
  assign n77020 = ~n77025;
  assign n73273 = n76983 ^ n76984;
  assign n76954 = n76986 ^ n76987;
  assign n76982 = n76989 & n76990;
  assign n76949 = n76987 & n76986;
  assign n73550 = n77006 ^ n77007;
  assign n76997 = ~n77010;
  assign n77013 = n77020 & n77021;
  assign n76968 = n76954 & n74325;
  assign n76963 = n73273 & n74359;
  assign n73280 = ~n73273;
  assign n76967 = ~n76954;
  assign n76943 = ~n76982;
  assign n76993 = n73550 & n76022;
  assign n73552 = ~n73550;
  assign n76980 = n76997 & n76998;
  assign n77000 = ~n77013;
  assign n76947 = ~n76963;
  assign n76962 = n76967 & n74305;
  assign n76953 = n76943 ^ n74325;
  assign n76930 = ~n76968;
  assign n76961 = n73280 & n76103;
  assign n76966 = n76980 ^ n76981;
  assign n76970 = n73552 & n74838;
  assign n76985 = n73552 & n76988;
  assign n76052 = ~n76993;
  assign n76978 = ~n76980;
  assign n76994 = n77000 & n77001;
  assign n73187 = n76953 ^ n76954;
  assign n76946 = ~n76961;
  assign n76942 = ~n76962;
  assign n76950 = n76966 ^ n2826;
  assign n76868 = n76969 ^ n76970;
  assign n76973 = ~n76970;
  assign n76976 = n76978 & n76979;
  assign n76016 = ~n76985;
  assign n76975 = n76994 ^ n74769;
  assign n76991 = ~n76994;
  assign n76931 = n73187 & n74325;
  assign n73198 = ~n73187;
  assign n76940 = n76942 & n76943;
  assign n76923 = n76946 & n76947;
  assign n76884 = n76949 ^ n76950;
  assign n76895 = n76950 & n76949;
  assign n76934 = n76973 & n76969;
  assign n73483 = n76974 ^ n76975;
  assign n76964 = ~n76976;
  assign n76977 = n76991 & n76992;
  assign n76909 = n76923 ^ n76924;
  assign n76921 = n73198 & n76085;
  assign n76900 = ~n76931;
  assign n76927 = ~n76923;
  assign n76929 = ~n76940;
  assign n76958 = n73483 & n75958;
  assign n76951 = n76964 & n76965;
  assign n73581 = ~n73483;
  assign n76971 = ~n76977;
  assign n76904 = n76909 & n102;
  assign n76901 = ~n76921;
  assign n76894 = ~n76909;
  assign n76877 = n76927 & n76928;
  assign n76898 = n76929 & n76930;
  assign n76925 = n76951 ^ n76938;
  assign n76952 = n73581 & n76957;
  assign n75997 = ~n76958;
  assign n76945 = n76951 & n2783;
  assign n76935 = n73581 & n74833;
  assign n76948 = ~n76951;
  assign n76955 = n76971 & n76972;
  assign n76892 = n76894 & n14810;
  assign n76881 = n76898 ^ n76884;
  assign n76878 = n76900 & n76901;
  assign n76850 = ~n76904;
  assign n76897 = n76898 & n74270;
  assign n76905 = ~n76898;
  assign n76896 = n84 ^ n76925;
  assign n76821 = n76934 ^ n76935;
  assign n76936 = ~n76935;
  assign n76937 = ~n76945;
  assign n76941 = n76948 & n84;
  assign n75964 = ~n76952;
  assign n76939 = n76955 ^ n76956;
  assign n76959 = ~n76955;
  assign n76823 = n76877 ^ n76878;
  assign n76875 = n76881 & n74288;
  assign n76876 = ~n76878;
  assign n76863 = ~n76881;
  assign n76871 = ~n76892;
  assign n76813 = n76895 ^ n76896;
  assign n76883 = ~n76897;
  assign n76893 = n76905 & n74288;
  assign n76912 = n76821 & n82;
  assign n76903 = ~n76896;
  assign n76913 = ~n76821;
  assign n76907 = n76936 & n76934;
  assign n76926 = n76937 & n76938;
  assign n73473 = n76939 ^ n74794;
  assign n76908 = n76939 & n74794;
  assign n76917 = ~n76941;
  assign n76944 = n76959 & n76960;
  assign n76846 = n76823 & n14752;
  assign n73109 = n76863 ^ n74270;
  assign n76848 = ~n76823;
  assign n76866 = n76871 & n76852;
  assign n76827 = ~n76875;
  assign n76851 = n76871 & n76850;
  assign n76803 = n76876 & n76877;
  assign n76873 = n76883 & n76884;
  assign n76872 = n76813 & n74247;
  assign n76870 = ~n76813;
  assign n76856 = ~n76893;
  assign n76832 = n76903 & n76895;
  assign n76769 = n76907 ^ n76908;
  assign n76796 = ~n76912;
  assign n76902 = n76913 & n2673;
  assign n76920 = n73473 & n76922;
  assign n73466 = ~n73473;
  assign n76911 = ~n76907;
  assign n76916 = ~n76926;
  assign n76910 = ~n76908;
  assign n76932 = ~n76944;
  assign n76824 = ~n76846;
  assign n76843 = n73109 & n75948;
  assign n76844 = n76848 & n101;
  assign n74791 = n76851 ^ n76852;
  assign n73104 = ~n73109;
  assign n76849 = ~n76866;
  assign n76814 = ~n76803;
  assign n76869 = n76870 & n74236;
  assign n76837 = ~n76872;
  assign n76855 = ~n76873;
  assign n76880 = n76769 & n81;
  assign n76885 = ~n76769;
  assign n76817 = ~n76902;
  assign n76906 = n73466 & n75892;
  assign n76854 = n76910 & n76911;
  assign n76887 = n76916 & n76917;
  assign n75925 = ~n76920;
  assign n76918 = n76932 & n76933;
  assign n76826 = ~n76843;
  assign n76800 = ~n76844;
  assign n74809 = ~n74791;
  assign n76822 = n76849 & n76850;
  assign n76838 = n76855 & n76856;
  assign n76810 = ~n76869;
  assign n76739 = ~n76880;
  assign n76874 = n76885 & n2621;
  assign n76859 = n76887 ^ n76868;
  assign n76891 = n76887 & n2766;
  assign n76888 = ~n76887;
  assign n76864 = ~n76854;
  assign n75889 = ~n76906;
  assign n76882 = n76918 ^ n76919;
  assign n76914 = ~n76918;
  assign n76801 = n76822 ^ n76823;
  assign n76802 = n76826 & n76827;
  assign n76812 = n76838 ^ n74236;
  assign n76825 = ~n76822;
  assign n76836 = ~n76838;
  assign n76833 = n76859 ^ n2766;
  assign n76763 = ~n76874;
  assign n73510 = n76882 ^ n74731;
  assign n76879 = n76888 & n83;
  assign n76867 = ~n76891;
  assign n76886 = ~n76882;
  assign n76899 = n76914 & n76915;
  assign n76781 = n101 ^ n76801;
  assign n76742 = n76802 ^ n76803;
  assign n73035 = n76812 ^ n76813;
  assign n76721 = n76802 & n76814;
  assign n76819 = n76824 & n76825;
  assign n76765 = n76832 ^ n76833;
  assign n76829 = n76836 & n76837;
  assign n76772 = n76833 & n76832;
  assign n76862 = n73510 & n76865;
  assign n76860 = n76867 & n76868;
  assign n73408 = ~n73510;
  assign n76842 = ~n76879;
  assign n76853 = n76886 & n74688;
  assign n76889 = ~n76899;
  assign n75766 = n76781 ^ n74791;
  assign n76788 = n73035 & n74236;
  assign n76776 = ~n76781;
  assign n73045 = ~n73035;
  assign n76727 = ~n76721;
  assign n76799 = ~n76819;
  assign n76809 = ~n76829;
  assign n76778 = ~n76772;
  assign n76686 = n76853 ^ n76854;
  assign n76841 = ~n76860;
  assign n76847 = n73408 & n75819;
  assign n75855 = ~n76862;
  assign n76791 = n76853 & n76864;
  assign n76861 = n76889 & n76890;
  assign n75756 = ~n75766;
  assign n76718 = n76776 & n74809;
  assign n76775 = n73045 & n75861;
  assign n76755 = ~n76788;
  assign n76782 = n76799 & n76800;
  assign n76789 = n76809 & n76810;
  assign n76820 = n76841 & n76842;
  assign n76840 = n76686 & n80;
  assign n75823 = ~n76847;
  assign n76839 = ~n76686;
  assign n76794 = ~n76791;
  assign n76831 = n76861 ^ n74649;
  assign n76857 = ~n76861;
  assign n76756 = ~n76775;
  assign n76741 = n100 ^ n76782;
  assign n76779 = n76782 & n14710;
  assign n76761 = n76789 ^ n76765;
  assign n76787 = n76789 & n74202;
  assign n76780 = ~n76782;
  assign n76786 = ~n76789;
  assign n76790 = n76820 ^ n76821;
  assign n73331 = n76830 ^ n76831;
  assign n76816 = ~n76820;
  assign n76828 = n76839 & n2593;
  assign n76681 = ~n76840;
  assign n76845 = n76857 & n76858;
  assign n76719 = n76741 ^ n76742;
  assign n76722 = n76755 & n76756;
  assign n76750 = n76761 & n74193;
  assign n76743 = ~n76761;
  assign n76758 = ~n76779;
  assign n76770 = n76780 & n100;
  assign n76777 = n76786 & n74193;
  assign n76764 = ~n76787;
  assign n76773 = n82 ^ n76790;
  assign n76792 = n73331 & n74649;
  assign n76811 = n76816 & n76817;
  assign n76815 = n73331 & n76818;
  assign n73366 = ~n73331;
  assign n76709 = ~n76828;
  assign n76834 = ~n76845;
  assign n74739 = n76718 ^ n76719;
  assign n76704 = n76721 ^ n76722;
  assign n76639 = n76719 & n76718;
  assign n72955 = n74193 ^ n76743;
  assign n76726 = ~n76722;
  assign n76689 = ~n76750;
  assign n76746 = n76742 & n76758;
  assign n76749 = n76764 & n76765;
  assign n76724 = ~n76770;
  assign n76678 = n76772 ^ n76773;
  assign n76734 = ~n76777;
  assign n76706 = n76773 & n76778;
  assign n76650 = n76791 ^ n76792;
  assign n76793 = ~n76792;
  assign n76798 = n73366 & n76806;
  assign n76795 = ~n76811;
  assign n75759 = ~n76815;
  assign n76807 = n76834 & n76835;
  assign n76694 = n76704 & n99;
  assign n75667 = ~n74739;
  assign n76642 = ~n76639;
  assign n76705 = ~n76704;
  assign n76663 = n76726 & n76727;
  assign n73005 = ~n72955;
  assign n76732 = n76678 & n74158;
  assign n76723 = ~n76746;
  assign n76733 = ~n76749;
  assign n76736 = ~n76678;
  assign n76713 = ~n76706;
  assign n76767 = n76650 & n95;
  assign n76766 = ~n76650;
  assign n76759 = n76793 & n76794;
  assign n76768 = n76795 & n76796;
  assign n75789 = ~n76798;
  assign n76785 = n76807 ^ n76808;
  assign n76804 = ~n76807;
  assign n76635 = ~n76694;
  assign n76687 = n76705 & n14678;
  assign n76716 = n73005 & n75834;
  assign n76703 = n76723 & n76724;
  assign n76683 = ~n76732;
  assign n76710 = n76733 & n76734;
  assign n76720 = n76736 & n74151;
  assign n76754 = n76766 & n2483;
  assign n76627 = ~n76767;
  assign n76737 = n76768 ^ n76769;
  assign n73257 = n74606 ^ n76785;
  assign n75791 = n75759 & n75789;
  assign n76762 = ~n76768;
  assign n76760 = n76785 & n74606;
  assign n76797 = n76804 & n76805;
  assign n76671 = ~n76687;
  assign n76673 = n76703 ^ n76704;
  assign n76679 = n76710 ^ n74151;
  assign n76688 = ~n76716;
  assign n76670 = ~n76703;
  assign n76714 = ~n76720;
  assign n76715 = ~n76710;
  assign n76707 = n81 ^ n76737;
  assign n76656 = ~n76754;
  assign n76593 = n76759 ^ n76760;
  assign n76751 = n76762 & n76763;
  assign n76757 = n73257 & n76771;
  assign n73426 = ~n73257;
  assign n76774 = ~n76760;
  assign n76783 = ~n76797;
  assign n76665 = n76670 & n76671;
  assign n76640 = n99 ^ n76673;
  assign n72900 = n76678 ^ n76679;
  assign n76666 = n76688 & n76689;
  assign n76622 = n76706 ^ n76707;
  assign n76700 = n76714 & n76715;
  assign n76712 = ~n76707;
  assign n76740 = n76593 & n2398;
  assign n76735 = ~n76593;
  assign n76738 = ~n76751;
  assign n76745 = n73426 & n75717;
  assign n75715 = ~n76757;
  assign n76693 = n76774 & n76759;
  assign n76752 = n76783 & n76784;
  assign n74679 = n76639 ^ n76640;
  assign n76641 = ~n76640;
  assign n76634 = ~n76665;
  assign n76660 = n72900 & n74158;
  assign n76617 = n76663 ^ n76666;
  assign n72916 = ~n72900;
  assign n76662 = ~n76666;
  assign n76677 = n76622 & n74103;
  assign n76684 = ~n76622;
  assign n76682 = ~n76700;
  assign n76659 = n76712 & n76713;
  assign n76725 = n76735 & n94;
  assign n76717 = n76738 & n76739;
  assign n76603 = ~n76740;
  assign n75688 = ~n76745;
  assign n76730 = n76752 ^ n76753;
  assign n76747 = ~n76752;
  assign n75602 = ~n74679;
  assign n76616 = n76634 & n76635;
  assign n76554 = n76641 & n76642;
  assign n76624 = ~n76660;
  assign n76636 = n72916 & n75703;
  assign n76595 = ~n76617;
  assign n76599 = n76662 & n76663;
  assign n76630 = ~n76677;
  assign n76657 = n76682 & n76683;
  assign n76667 = n76684 & n74118;
  assign n76685 = n80 ^ n76717;
  assign n76577 = ~n76725;
  assign n73383 = n76730 ^ n74618;
  assign n76708 = ~n76717;
  assign n76731 = ~n76730;
  assign n76744 = n76747 & n76748;
  assign n76585 = n76616 ^ n76617;
  assign n76620 = n76616 & n14640;
  assign n76553 = ~n76554;
  assign n76613 = ~n76616;
  assign n76623 = ~n76636;
  assign n76621 = n76657 ^ n74103;
  assign n76653 = ~n76667;
  assign n76652 = ~n76657;
  assign n76661 = n76685 ^ n76686;
  assign n76699 = n76708 & n76709;
  assign n76696 = n73383 & n76711;
  assign n73228 = ~n73383;
  assign n76695 = n76731 & n74571;
  assign n76728 = ~n76744;
  assign n76555 = n98 ^ n76585;
  assign n76608 = n76613 & n98;
  assign n76594 = ~n76620;
  assign n72844 = n76621 ^ n76622;
  assign n76600 = n76623 & n76624;
  assign n76646 = n76652 & n76653;
  assign n76567 = n76659 ^ n76661;
  assign n76658 = ~n76661;
  assign n76546 = n76693 ^ n76695;
  assign n75645 = ~n76696;
  assign n76680 = ~n76699;
  assign n76690 = n73228 & n75656;
  assign n76692 = ~n76695;
  assign n76701 = n76728 & n76729;
  assign n74636 = n76554 ^ n76555;
  assign n76552 = ~n76555;
  assign n76581 = n76594 & n76595;
  assign n76544 = n76599 ^ n76600;
  assign n76574 = ~n76608;
  assign n76591 = n72844 & n75627;
  assign n72880 = ~n72844;
  assign n76601 = ~n76600;
  assign n76631 = n76567 & n74096;
  assign n76628 = ~n76567;
  assign n76629 = ~n76646;
  assign n76596 = n76658 & n76659;
  assign n76675 = n76546 & n2323;
  assign n76649 = n76680 & n76681;
  assign n76676 = ~n76546;
  assign n75625 = ~n76690;
  assign n76645 = n76692 & n76693;
  assign n76672 = n76701 ^ n76702;
  assign n76697 = ~n76701;
  assign n75513 = ~n74636;
  assign n76480 = n76552 & n76553;
  assign n76578 = n76544 & n14600;
  assign n76573 = ~n76581;
  assign n76568 = ~n76544;
  assign n76586 = n72880 & n74103;
  assign n76565 = ~n76591;
  assign n76549 = n76601 & n76599;
  assign n76610 = n76628 & n74067;
  assign n76607 = n76629 & n76630;
  assign n76606 = ~n76631;
  assign n76625 = n76649 ^ n76650;
  assign n76655 = ~n76649;
  assign n73335 = n76672 ^ n74577;
  assign n76542 = ~n76675;
  assign n76664 = n76676 & n93;
  assign n76651 = ~n76645;
  assign n76674 = ~n76672;
  assign n76691 = n76697 & n76698;
  assign n76561 = n76568 & n97;
  assign n76543 = n76573 & n76574;
  assign n76539 = ~n76578;
  assign n76551 = ~n76549;
  assign n76564 = ~n76586;
  assign n76566 = n76607 ^ n74067;
  assign n76570 = ~n76610;
  assign n76605 = ~n76607;
  assign n76597 = n95 ^ n76625;
  assign n76648 = n73335 & n76654;
  assign n76647 = n76655 & n76656;
  assign n76513 = ~n76664;
  assign n73171 = ~n73335;
  assign n76644 = n76674 & n74529;
  assign n76668 = ~n76691;
  assign n76504 = n76543 ^ n76544;
  assign n76503 = ~n76561;
  assign n76538 = ~n76543;
  assign n76548 = n76564 & n76565;
  assign n72799 = n76566 ^ n76567;
  assign n76507 = n76596 ^ n76597;
  assign n76589 = n76605 & n76606;
  assign n76604 = ~n76597;
  assign n76492 = n76644 ^ n76645;
  assign n76633 = n73171 & n75554;
  assign n76626 = ~n76647;
  assign n75590 = ~n76648;
  assign n76557 = n76644 & n76651;
  assign n76643 = n76668 & n76669;
  assign n76481 = n97 ^ n76504;
  assign n76527 = n76538 & n76539;
  assign n76460 = n76548 ^ n76549;
  assign n76540 = n72799 & n74067;
  assign n76477 = n76548 & n76551;
  assign n72808 = ~n72799;
  assign n76571 = n76507 & n74024;
  assign n76569 = ~n76589;
  assign n76572 = ~n76507;
  assign n76534 = n76604 & n76596;
  assign n76614 = n76492 & n92;
  assign n76592 = n76626 & n76627;
  assign n76615 = ~n76492;
  assign n75547 = ~n76633;
  assign n76619 = n76643 ^ n74474;
  assign n76637 = ~n76643;
  assign n74596 = n76480 ^ n76481;
  assign n76487 = ~n76481;
  assign n76502 = ~n76527;
  assign n76515 = ~n76540;
  assign n76520 = n72808 & n75613;
  assign n76547 = n76569 & n76570;
  assign n76537 = ~n76571;
  assign n76559 = n76572 & n74051;
  assign n76575 = n76592 ^ n76593;
  assign n76602 = ~n76592;
  assign n76453 = ~n76614;
  assign n76609 = n76615 & n2217;
  assign n73117 = n76618 ^ n76619;
  assign n76632 = n76637 & n76638;
  assign n75439 = ~n74596;
  assign n76434 = n76487 & n76480;
  assign n76484 = n76502 & n76503;
  assign n76514 = ~n76520;
  assign n76508 = n76547 ^ n74024;
  assign n76536 = ~n76547;
  assign n76511 = ~n76559;
  assign n76535 = n94 ^ n76575;
  assign n76582 = n73117 & n76598;
  assign n76590 = n76602 & n76603;
  assign n73111 = ~n73117;
  assign n76479 = ~n76609;
  assign n76611 = ~n76632;
  assign n76451 = n76484 ^ n76460;
  assign n76485 = n76484 & n14563;
  assign n76493 = ~n76484;
  assign n72749 = n76507 ^ n76508;
  assign n76476 = n76514 & n76515;
  assign n76458 = n76534 ^ n76535;
  assign n76532 = n76536 & n76537;
  assign n76482 = n76535 & n76534;
  assign n75519 = ~n76582;
  assign n76580 = n73111 & n75515;
  assign n76558 = n73111 & n74474;
  assign n76576 = ~n76590;
  assign n76583 = n76611 & n76612;
  assign n76435 = n96 ^ n76451;
  assign n76413 = n76476 ^ n76477;
  assign n76461 = ~n76485;
  assign n76465 = n76493 & n96;
  assign n76424 = n76476 & n76477;
  assign n76486 = n72749 & n75466;
  assign n72747 = ~n72749;
  assign n76509 = n76458 & n73990;
  assign n76506 = ~n76458;
  assign n76510 = ~n76532;
  assign n76490 = ~n76482;
  assign n76429 = n76557 ^ n76558;
  assign n76545 = n76576 & n76577;
  assign n76560 = ~n76558;
  assign n75477 = ~n76580;
  assign n76556 = n76583 ^ n76584;
  assign n76587 = ~n76583;
  assign n74551 = n76434 ^ n76435;
  assign n76369 = n76435 & n76434;
  assign n76449 = n76460 & n76461;
  assign n76440 = ~n76465;
  assign n76397 = ~n76413;
  assign n76464 = n72747 & n74051;
  assign n76447 = ~n76486;
  assign n76501 = n76506 & n73988;
  assign n76455 = ~n76509;
  assign n76488 = n76510 & n76511;
  assign n76519 = n76429 & n91;
  assign n76505 = n76545 ^ n76546;
  assign n76524 = ~n76429;
  assign n73033 = n76556 ^ n74421;
  assign n76541 = ~n76545;
  assign n76528 = n76560 & n76557;
  assign n76529 = n76556 & n74421;
  assign n76579 = n76587 & n76588;
  assign n75380 = ~n74551;
  assign n76372 = ~n76369;
  assign n76439 = ~n76449;
  assign n76448 = ~n76464;
  assign n76459 = n76488 ^ n73988;
  assign n76474 = ~n76488;
  assign n76475 = ~n76501;
  assign n76483 = n93 ^ n76505;
  assign n76407 = ~n76519;
  assign n76517 = n76524 & n2139;
  assign n76378 = n76528 ^ n76529;
  assign n76533 = n76541 & n76542;
  assign n76521 = n73033 & n76550;
  assign n73210 = ~n73033;
  assign n76526 = ~n76528;
  assign n76525 = ~n76529;
  assign n76562 = ~n76579;
  assign n76412 = n76439 & n76440;
  assign n76425 = n76447 & n76448;
  assign n72710 = n76458 ^ n76459;
  assign n76463 = n76474 & n76475;
  assign n76411 = n76482 ^ n76483;
  assign n76489 = ~n76483;
  assign n76495 = n76378 & n90;
  assign n76500 = ~n76378;
  assign n76427 = ~n76517;
  assign n75436 = ~n76521;
  assign n76466 = n76525 & n76526;
  assign n76516 = n73210 & n75398;
  assign n76512 = ~n76533;
  assign n76530 = n76562 & n76563;
  assign n76393 = n76412 ^ n76413;
  assign n76415 = n76412 & n14517;
  assign n76351 = n76424 ^ n76425;
  assign n76414 = ~n76412;
  assign n76423 = n72710 & n73990;
  assign n76390 = n76425 & n76424;
  assign n72715 = ~n72710;
  assign n76457 = n76411 & n73985;
  assign n76454 = ~n76463;
  assign n76456 = ~n76411;
  assign n76430 = n76489 & n76490;
  assign n76368 = ~n76495;
  assign n76494 = n76500 & n2082;
  assign n76491 = n76512 & n76513;
  assign n75402 = ~n76516;
  assign n76499 = n76530 ^ n76531;
  assign n76522 = ~n76530;
  assign n76370 = n111 ^ n76393;
  assign n76405 = n76351 & n14497;
  assign n76400 = n76414 & n111;
  assign n76396 = ~n76415;
  assign n76403 = ~n76351;
  assign n76399 = ~n76423;
  assign n76387 = ~n76390;
  assign n76422 = n72715 & n75387;
  assign n76438 = n76454 & n76455;
  assign n76446 = n76456 & n73936;
  assign n76432 = ~n76457;
  assign n76437 = ~n76430;
  assign n76450 = n76491 ^ n76492;
  assign n76381 = ~n76494;
  assign n76478 = ~n76491;
  assign n72983 = n76499 ^ n74448;
  assign n76498 = ~n76499;
  assign n76518 = n76522 & n76523;
  assign n74511 = n76369 ^ n76370;
  assign n76313 = n76370 & n76372;
  assign n76392 = n76396 & n76397;
  assign n76374 = ~n76400;
  assign n76395 = n76403 & n110;
  assign n76354 = ~n76405;
  assign n76398 = ~n76422;
  assign n76410 = n76438 ^ n73936;
  assign n76433 = ~n76438;
  assign n76409 = ~n76446;
  assign n76431 = n92 ^ n76450;
  assign n76473 = n76478 & n76479;
  assign n76471 = n72983 & n75339;
  assign n72974 = ~n72983;
  assign n76467 = n76498 & n74379;
  assign n76496 = ~n76518;
  assign n75318 = ~n74511;
  assign n76312 = ~n76313;
  assign n76373 = ~n76392;
  assign n76332 = ~n76395;
  assign n76391 = n76398 & n76399;
  assign n72665 = n76410 ^ n76411;
  assign n76360 = n76430 ^ n76431;
  assign n76421 = n76432 & n76433;
  assign n76436 = ~n76431;
  assign n76342 = n76466 ^ n76467;
  assign n76462 = n72974 & n76468;
  assign n75351 = ~n76471;
  assign n76452 = ~n76473;
  assign n76472 = ~n76467;
  assign n76469 = n76496 & n76497;
  assign n76350 = n76373 & n76374;
  assign n76310 = n76390 ^ n76391;
  assign n76379 = n72665 & n73936;
  assign n72714 = ~n72665;
  assign n76386 = ~n76391;
  assign n76402 = n76360 & n73938;
  assign n76404 = ~n76360;
  assign n76408 = ~n76421;
  assign n76383 = n76436 & n76437;
  assign n76428 = n76452 & n76453;
  assign n76444 = n76342 & n2029;
  assign n76445 = ~n76342;
  assign n75379 = ~n76462;
  assign n73123 = n76469 ^ n76470;
  assign n76419 = n76472 & n76466;
  assign n76330 = n76350 ^ n76351;
  assign n76366 = n76310 & n109;
  assign n76355 = ~n76350;
  assign n76362 = ~n76310;
  assign n76376 = n72714 & n75357;
  assign n76356 = ~n76379;
  assign n76336 = n76386 & n76387;
  assign n76359 = ~n76402;
  assign n76394 = n76404 & n73898;
  assign n76389 = n76408 & n76409;
  assign n76401 = n76428 ^ n76429;
  assign n76416 = n76443 ^ n73123;
  assign n76340 = ~n76444;
  assign n76426 = ~n76428;
  assign n76441 = n76445 & n89;
  assign n76442 = ~n73123;
  assign n76314 = n110 ^ n76330;
  assign n76347 = n76354 & n76355;
  assign n76353 = n76362 & n14444;
  assign n76293 = ~n76366;
  assign n76349 = ~n76336;
  assign n76357 = ~n76376;
  assign n76361 = n76389 ^ n73898;
  assign n76385 = ~n76394;
  assign n76384 = ~n76389;
  assign n76388 = n91 ^ n76401;
  assign n75315 = n76416 ^ n76417;
  assign n76418 = n76426 & n76427;
  assign n76319 = ~n76441;
  assign n76420 = n76442 & n74423;
  assign n75281 = n76313 ^ n76314;
  assign n76311 = ~n76314;
  assign n76331 = ~n76347;
  assign n76317 = ~n76353;
  assign n76335 = n76356 & n76357;
  assign n72634 = n76360 ^ n76361;
  assign n76371 = n76384 & n76385;
  assign n76322 = n76383 ^ n76388;
  assign n76382 = ~n76388;
  assign n76406 = ~n76418;
  assign n76297 = n76419 ^ n76420;
  assign n76276 = n76311 & n76312;
  assign n76309 = n76331 & n76332;
  assign n76264 = n76335 ^ n76336;
  assign n76338 = n72634 & n73938;
  assign n76301 = n76335 & n76349;
  assign n72638 = ~n72634;
  assign n76364 = n76322 & n73855;
  assign n76358 = ~n76371;
  assign n76363 = ~n76322;
  assign n76343 = n76382 & n76383;
  assign n76377 = n76406 & n76407;
  assign n76291 = n76309 ^ n76310;
  assign n76316 = ~n76309;
  assign n76320 = ~n76338;
  assign n76306 = ~n76301;
  assign n76334 = n72638 & n75275;
  assign n76337 = n76358 & n76359;
  assign n76352 = n76363 & n73895;
  assign n76346 = ~n76364;
  assign n76348 = ~n76343;
  assign n76365 = n76377 ^ n76378;
  assign n76380 = ~n76377;
  assign n76277 = n109 ^ n76291;
  assign n76308 = n76316 & n76317;
  assign n76321 = ~n76334;
  assign n76323 = n76337 ^ n73855;
  assign n76345 = ~n76337;
  assign n76328 = ~n76352;
  assign n76344 = n90 ^ n76365;
  assign n76375 = n76380 & n76381;
  assign n76259 = n76276 ^ n76277;
  assign n76239 = n76277 & n76276;
  assign n76292 = ~n76308;
  assign n76302 = n76320 & n76321;
  assign n72581 = n76322 ^ n76323;
  assign n76288 = n76343 ^ n76344;
  assign n76329 = n76345 & n76346;
  assign n76299 = n76344 & n76348;
  assign n76367 = ~n76375;
  assign n72331 = n76259 ^ n73380;
  assign n76256 = n76259 & n73382;
  assign n76255 = ~n76259;
  assign n76275 = n76292 & n76293;
  assign n76230 = n76301 ^ n76302;
  assign n76298 = n72581 & n75215;
  assign n72609 = ~n72581;
  assign n76305 = ~n76302;
  assign n76326 = n76288 & n73810;
  assign n76327 = ~n76329;
  assign n76325 = ~n76288;
  assign n76307 = ~n76299;
  assign n76341 = n76367 & n76368;
  assign n76241 = ~n72331;
  assign n76174 = n76255 & n73382;
  assign n76224 = ~n76256;
  assign n76253 = n76275 ^ n76264;
  assign n76278 = n76275 & n14397;
  assign n76282 = n76230 & n107;
  assign n76273 = ~n76275;
  assign n76281 = ~n76230;
  assign n76294 = n72609 & n73895;
  assign n76287 = ~n76298;
  assign n76267 = n76305 & n76306;
  assign n76315 = n76325 & n73815;
  assign n76280 = ~n76326;
  assign n76295 = n76327 & n76328;
  assign n76324 = n76341 ^ n76342;
  assign n76339 = ~n76341;
  assign n76238 = n76241 & n74445;
  assign n76240 = n108 ^ n76253;
  assign n76271 = n76273 & n108;
  assign n76263 = ~n76278;
  assign n76272 = n76281 & n14377;
  assign n76214 = ~n76282;
  assign n76270 = ~n76267;
  assign n76286 = ~n76294;
  assign n76289 = n76295 ^ n73815;
  assign n76304 = ~n76295;
  assign n76303 = ~n76315;
  assign n76300 = n89 ^ n76324;
  assign n76333 = n76339 & n76340;
  assign n76223 = ~n76238;
  assign n76235 = n76239 ^ n76240;
  assign n76194 = n76240 & n76239;
  assign n76257 = n76263 & n76264;
  assign n76244 = ~n76271;
  assign n76228 = ~n76272;
  assign n76266 = n76286 & n76287;
  assign n72544 = n76288 ^ n76289;
  assign n76251 = n76299 ^ n76300;
  assign n76290 = n76303 & n76304;
  assign n76268 = n76300 & n76307;
  assign n76318 = ~n76333;
  assign n76198 = n76223 & n76224;
  assign n76220 = n76235 & n73280;
  assign n76221 = ~n76235;
  assign n76186 = ~n76194;
  assign n76243 = ~n76257;
  assign n76173 = n76266 ^ n76267;
  assign n76232 = n76266 & n76270;
  assign n76262 = n72544 & n73810;
  assign n72553 = ~n72544;
  assign n76284 = n76251 & n73825;
  assign n76279 = ~n76290;
  assign n76285 = ~n76251;
  assign n76296 = n76318 & n76319;
  assign n76176 = n76198 ^ n76199;
  assign n76203 = ~n76198;
  assign n76202 = ~n76220;
  assign n76217 = n76221 & n73273;
  assign n76229 = n76243 & n76244;
  assign n76237 = ~n76232;
  assign n76245 = ~n76262;
  assign n76258 = n72553 & n75140;
  assign n76265 = n76279 & n76280;
  assign n76261 = ~n76284;
  assign n76274 = n76285 & n73761;
  assign n76283 = n76296 ^ n76297;
  assign n74165 = n135 ^ n76176;
  assign n75949 = n76176 & n135;
  assign n76045 = n76203 & n76204;
  assign n76200 = n76202 & n76174;
  assign n76182 = ~n76217;
  assign n76206 = n76229 ^ n76230;
  assign n76227 = ~n76229;
  assign n76246 = ~n76258;
  assign n76250 = n76265 ^ n73761;
  assign n76249 = ~n76274;
  assign n76260 = ~n76265;
  assign n76269 = n88 ^ n76283;
  assign n74191 = ~n74165;
  assign n76181 = ~n76200;
  assign n76197 = n76182 & n76202;
  assign n76195 = n107 ^ n76206;
  assign n76219 = n76227 & n76228;
  assign n76233 = n76245 & n76246;
  assign n72496 = n76250 ^ n76251;
  assign n76254 = n76260 & n76261;
  assign n76211 = n76268 ^ n76269;
  assign n76170 = n76181 & n76182;
  assign n76171 = n76194 ^ n76195;
  assign n76175 = ~n76197;
  assign n76185 = ~n76195;
  assign n76213 = ~n76219;
  assign n76216 = n76232 ^ n76233;
  assign n76234 = n72496 & n73761;
  assign n72557 = ~n72496;
  assign n76236 = ~n76233;
  assign n76252 = n76211 & n73798;
  assign n76248 = ~n76254;
  assign n76247 = ~n76211;
  assign n76140 = n76170 ^ n76171;
  assign n76169 = n76171 & n73187;
  assign n72201 = n76174 ^ n76175;
  assign n76149 = ~n76170;
  assign n76160 = ~n76171;
  assign n76146 = n76185 & n76186;
  assign n76190 = n76213 & n76214;
  assign n76205 = n76216 & n105;
  assign n76215 = ~n76216;
  assign n76209 = ~n76234;
  assign n76222 = n72557 & n75078;
  assign n76184 = n76236 & n76237;
  assign n76242 = n76247 & n73701;
  assign n76231 = n76248 & n76249;
  assign n76226 = ~n76252;
  assign n72098 = n73187 ^ n76140;
  assign n76152 = n76140 & n73187;
  assign n76153 = n72201 & n74359;
  assign n72191 = ~n72201;
  assign n76157 = n76160 & n73198;
  assign n76129 = ~n76169;
  assign n76163 = n76190 ^ n76173;
  assign n76191 = n76190 & n14316;
  assign n76180 = ~n76190;
  assign n76106 = ~n76205;
  assign n76201 = n76215 & n14279;
  assign n76196 = ~n76184;
  assign n76210 = ~n76222;
  assign n76212 = n76231 ^ n73701;
  assign n76225 = ~n76231;
  assign n76208 = ~n76242;
  assign n76125 = n72098 & n74325;
  assign n72117 = ~n72098;
  assign n76110 = ~n76152;
  assign n76131 = ~n76153;
  assign n76142 = n72191 & n73273;
  assign n76150 = ~n76157;
  assign n76151 = n106 ^ n76163;
  assign n76177 = n76180 & n106;
  assign n76172 = ~n76191;
  assign n76134 = ~n76201;
  assign n76183 = n76209 & n76210;
  assign n72459 = n76211 ^ n76212;
  assign n76218 = n76225 & n76226;
  assign n76109 = ~n76125;
  assign n76130 = ~n76142;
  assign n76137 = n76149 & n76150;
  assign n76066 = n76146 ^ n76151;
  assign n76145 = ~n76151;
  assign n76159 = n76172 & n76173;
  assign n76155 = ~n76177;
  assign n76083 = n76183 ^ n76184;
  assign n76135 = n76134 & n76106;
  assign n76187 = n72459 & n73701;
  assign n76144 = n76183 & n76196;
  assign n72467 = ~n72459;
  assign n76207 = ~n76218;
  assign n76041 = n76109 & n76110;
  assign n76120 = n76066 & n73109;
  assign n76114 = n76130 & n76131;
  assign n76116 = ~n76066;
  assign n76128 = ~n76137;
  assign n76107 = n76145 & n76146;
  assign n76154 = ~n76159;
  assign n76166 = n76083 & n104;
  assign n76164 = ~n76083;
  assign n76162 = ~n76187;
  assign n76179 = n72467 & n74986;
  assign n76192 = n76207 & n76208;
  assign n76079 = n76041 & n76009;
  assign n76084 = ~n76041;
  assign n76104 = n76114 & n76115;
  assign n76112 = n76116 & n73104;
  assign n76102 = ~n76114;
  assign n76100 = ~n76120;
  assign n76090 = n76128 & n76129;
  assign n76113 = ~n76107;
  assign n76136 = n76154 & n76155;
  assign n76156 = n76164 & n14245;
  assign n76057 = ~n76166;
  assign n76161 = ~n76179;
  assign n76165 = n76192 ^ n76193;
  assign n76188 = ~n76192;
  assign n76037 = ~n76079;
  assign n76071 = n76084 & n76085;
  assign n76067 = n76090 ^ n73109;
  assign n76101 = n76102 & n76103;
  assign n76080 = ~n76104;
  assign n76099 = ~n76090;
  assign n76070 = ~n76112;
  assign n76108 = n76135 ^ n76136;
  assign n76133 = ~n76136;
  assign n76078 = ~n76156;
  assign n76143 = n76161 & n76162;
  assign n72387 = n73663 ^ n76165;
  assign n76158 = n76165 & n73744;
  assign n76178 = n76188 & n76189;
  assign n72029 = n76066 ^ n76067;
  assign n76011 = ~n76071;
  assign n76081 = n76080 & n76045;
  assign n76086 = n76099 & n76100;
  assign n76061 = ~n76101;
  assign n76012 = n76107 ^ n76108;
  assign n76026 = n76108 & n76113;
  assign n76117 = n76133 & n76134;
  assign n76132 = n76143 ^ n76144;
  assign n76094 = n76143 & n76144;
  assign n72487 = ~n72387;
  assign n76122 = ~n76158;
  assign n76167 = ~n76178;
  assign n76044 = n72029 & n74288;
  assign n72025 = ~n72029;
  assign n76065 = n76061 & n76080;
  assign n76060 = ~n76081;
  assign n76069 = ~n76086;
  assign n76105 = ~n76117;
  assign n76119 = n76132 & n14200;
  assign n76118 = ~n76132;
  assign n76092 = ~n76094;
  assign n76138 = n72487 & n74963;
  assign n76141 = n76167 & n76168;
  assign n76018 = ~n76044;
  assign n76036 = n72025 & n73104;
  assign n76040 = n76060 & n76061;
  assign n76046 = ~n76065;
  assign n76054 = n76069 & n76070;
  assign n76082 = n76105 & n76106;
  assign n76111 = n76118 & n119;
  assign n76033 = ~n76119;
  assign n76121 = ~n76138;
  assign n76126 = n76141 ^ n73626;
  assign n76147 = ~n76141;
  assign n76017 = ~n76036;
  assign n76008 = n76040 ^ n76041;
  assign n76034 = n76045 ^ n76046;
  assign n76013 = n76054 ^ n73035;
  assign n76038 = ~n76040;
  assign n76049 = n76054 & n73045;
  assign n76043 = ~n76054;
  assign n76058 = n76082 ^ n76083;
  assign n76077 = ~n76082;
  assign n76002 = ~n76111;
  assign n76095 = n76121 & n76122;
  assign n72364 = n76126 ^ n76127;
  assign n76139 = n76147 & n76148;
  assign n75934 = n76008 ^ n76009;
  assign n71928 = n76012 ^ n76013;
  assign n75982 = n76017 & n76018;
  assign n76014 = n76034 & n6633;
  assign n76030 = n76037 & n76038;
  assign n76021 = ~n76034;
  assign n76035 = n76043 & n73035;
  assign n76031 = ~n76049;
  assign n76027 = n104 ^ n76058;
  assign n76068 = n76077 & n76078;
  assign n75969 = n76094 ^ n76095;
  assign n76088 = n76002 & n76033;
  assign n76093 = n72364 & n73626;
  assign n76091 = ~n76095;
  assign n72450 = ~n72364;
  assign n76123 = ~n76139;
  assign n75986 = n75934 & n6535;
  assign n75998 = n71928 & n74236;
  assign n75991 = n75982 & n76006;
  assign n75985 = ~n75934;
  assign n71934 = ~n71928;
  assign n75993 = ~n75982;
  assign n75990 = ~n76014;
  assign n76007 = n76021 & n134;
  assign n75940 = n76026 ^ n76027;
  assign n76010 = ~n76030;
  assign n76024 = n76031 & n76012;
  assign n76000 = ~n76035;
  assign n76004 = n76027 & n76026;
  assign n76056 = ~n76068;
  assign n76062 = n75969 & n118;
  assign n76029 = ~n76088;
  assign n76074 = ~n75969;
  assign n76048 = n76091 & n76092;
  assign n76075 = ~n76093;
  assign n76087 = n72450 & n74899;
  assign n76096 = n76123 & n76124;
  assign n75978 = n75985 & n133;
  assign n75937 = ~n75986;
  assign n75971 = ~n75991;
  assign n75979 = n75993 & n75948;
  assign n75987 = n71934 & n73035;
  assign n75956 = ~n75998;
  assign n75989 = n75990 & n75949;
  assign n75975 = ~n76007;
  assign n75981 = n76010 & n76011;
  assign n75946 = ~n75940;
  assign n75999 = ~n76024;
  assign n76028 = n76056 & n76057;
  assign n75936 = ~n76062;
  assign n76059 = n76074 & n14171;
  assign n76076 = ~n76087;
  assign n76055 = ~n76048;
  assign n76073 = n76096 ^ n73593;
  assign n76097 = ~n76096;
  assign n75908 = ~n75978;
  assign n75932 = ~n75979;
  assign n75947 = n75981 ^ n75982;
  assign n75955 = ~n75987;
  assign n75974 = ~n75989;
  assign n75983 = n75990 & n75975;
  assign n75966 = n75999 & n76000;
  assign n75970 = ~n75981;
  assign n76005 = n76028 ^ n76029;
  assign n76032 = ~n76028;
  assign n75977 = ~n76059;
  assign n72316 = n76072 ^ n76073;
  assign n76047 = n76075 & n76076;
  assign n76089 = n76097 & n76098;
  assign n75872 = n75947 ^ n75948;
  assign n75900 = n75955 & n75956;
  assign n75941 = n75966 ^ n72955;
  assign n75951 = n75970 & n75971;
  assign n75933 = n75974 & n75975;
  assign n75950 = ~n75983;
  assign n75965 = n75966 & n73005;
  assign n75967 = ~n75966;
  assign n75847 = n76004 ^ n76005;
  assign n76003 = ~n76005;
  assign n76025 = n76032 & n76033;
  assign n75880 = n76047 ^ n76048;
  assign n75994 = n76047 & n76055;
  assign n76053 = n72316 & n74857;
  assign n72403 = ~n72316;
  assign n76063 = ~n76089;
  assign n75915 = n75872 & n132;
  assign n75903 = n75933 ^ n75934;
  assign n71828 = n75940 ^ n75941;
  assign n75916 = ~n75872;
  assign n75923 = n75900 & n75942;
  assign n75922 = ~n75900;
  assign n75919 = n75949 ^ n75950;
  assign n75931 = ~n75951;
  assign n75938 = ~n75933;
  assign n75945 = ~n75965;
  assign n75954 = n75967 & n72955;
  assign n75973 = n75847 & n72900;
  assign n75972 = ~n75847;
  assign n75909 = n76003 & n76004;
  assign n76001 = ~n76025;
  assign n76042 = n72403 & n73660;
  assign n76019 = ~n76053;
  assign n76050 = n76063 & n76064;
  assign n75863 = n133 ^ n75903;
  assign n75830 = ~n75915;
  assign n75911 = n75916 & n6467;
  assign n75682 = n75919 ^ n74191;
  assign n75906 = n71828 & n72955;
  assign n71872 = ~n71828;
  assign n75912 = n75922 & n75861;
  assign n75902 = ~n75923;
  assign n75862 = n75919 & n74191;
  assign n75899 = n75931 & n75932;
  assign n75928 = n75937 & n75938;
  assign n75943 = n75945 & n75946;
  assign n75918 = ~n75954;
  assign n75957 = n75972 & n72916;
  assign n75843 = ~n75973;
  assign n75897 = ~n75909;
  assign n75968 = n76001 & n76002;
  assign n76020 = ~n76042;
  assign n76023 = n76050 ^ n73550;
  assign n76051 = ~n76050;
  assign n74108 = n75862 ^ n75863;
  assign n75875 = ~n75863;
  assign n74143 = ~n75682;
  assign n75860 = n75899 ^ n75900;
  assign n75894 = n71872 & n74193;
  assign n75874 = ~n75906;
  assign n75868 = ~n75911;
  assign n75867 = ~n75912;
  assign n75901 = ~n75899;
  assign n75907 = ~n75928;
  assign n75917 = ~n75943;
  assign n75882 = ~n75957;
  assign n75939 = n75968 ^ n75969;
  assign n75976 = ~n75968;
  assign n75995 = n76019 & n76020;
  assign n72268 = n76022 ^ n76023;
  assign n76039 = n76051 & n76052;
  assign n75595 = ~n74108;
  assign n75799 = n75860 ^ n75861;
  assign n75802 = n75875 & n75862;
  assign n75873 = ~n75894;
  assign n75890 = n75901 & n75902;
  assign n75871 = n75907 & n75908;
  assign n75884 = n75917 & n75918;
  assign n75910 = n118 ^ n75939;
  assign n75960 = n75976 & n75977;
  assign n75808 = n75994 ^ n75995;
  assign n75920 = n75995 & n75994;
  assign n75992 = n72268 & n74838;
  assign n72359 = ~n72268;
  assign n76015 = ~n76039;
  assign n75832 = n75799 & n131;
  assign n75831 = ~n75799;
  assign n75837 = n75871 ^ n75872;
  assign n75796 = n75873 & n75874;
  assign n75848 = n75884 ^ n72900;
  assign n75869 = ~n75871;
  assign n75866 = ~n75890;
  assign n75881 = ~n75884;
  assign n75812 = n75909 ^ n75910;
  assign n75896 = ~n75910;
  assign n75935 = ~n75960;
  assign n75961 = n75808 & n14072;
  assign n75962 = ~n75808;
  assign n75980 = n72359 & n73552;
  assign n75953 = ~n75992;
  assign n75927 = ~n75920;
  assign n75988 = n76015 & n76016;
  assign n75825 = n75831 & n6372;
  assign n75771 = ~n75832;
  assign n75803 = n132 ^ n75837;
  assign n71750 = n75847 ^ n75848;
  assign n75828 = n75796 & n75836;
  assign n75833 = ~n75796;
  assign n75835 = n75866 & n75867;
  assign n75858 = n75868 & n75869;
  assign n75876 = n75812 & n72880;
  assign n75878 = n75881 & n75882;
  assign n75864 = ~n75812;
  assign n75838 = n75896 & n75897;
  assign n75898 = n75935 & n75936;
  assign n75814 = ~n75961;
  assign n75944 = n75962 & n116;
  assign n75952 = ~n75980;
  assign n75959 = n75988 ^ n73483;
  assign n75996 = ~n75988;
  assign n74074 = n75802 ^ n75803;
  assign n75726 = n75803 & n75802;
  assign n75800 = ~n75825;
  assign n75815 = n71750 & n74158;
  assign n75810 = ~n75828;
  assign n75827 = n75833 & n75834;
  assign n71769 = ~n71750;
  assign n75797 = n75835 ^ n75836;
  assign n75809 = ~n75835;
  assign n75829 = ~n75858;
  assign n75856 = n75864 & n72844;
  assign n75778 = ~n75876;
  assign n75842 = ~n75878;
  assign n75841 = ~n75838;
  assign n75870 = n75898 ^ n75880;
  assign n75904 = n75898 & n14111;
  assign n75905 = ~n75898;
  assign n75776 = ~n75944;
  assign n75921 = n75952 & n75953;
  assign n72217 = n75958 ^ n75959;
  assign n75984 = n75996 & n75997;
  assign n75524 = ~n74074;
  assign n75736 = n75796 ^ n75797;
  assign n75732 = ~n75726;
  assign n75805 = n75809 & n75810;
  assign n75795 = n71769 & n72900;
  assign n75784 = ~n75815;
  assign n75780 = ~n75827;
  assign n75798 = n75829 & n75830;
  assign n75811 = n75842 & n75843;
  assign n75817 = ~n75856;
  assign n75839 = n117 ^ n75870;
  assign n75879 = ~n75904;
  assign n75895 = n75905 & n117;
  assign n75753 = n75920 ^ n75921;
  assign n75929 = n72217 & n74833;
  assign n72320 = ~n72217;
  assign n75926 = ~n75921;
  assign n75963 = ~n75984;
  assign n75769 = n75736 & n6286;
  assign n75768 = ~n75736;
  assign n75783 = ~n75795;
  assign n75767 = n75798 ^ n75799;
  assign n75779 = ~n75805;
  assign n75772 = n75811 ^ n75812;
  assign n75801 = ~n75798;
  assign n75816 = ~n75811;
  assign n75710 = n75838 ^ n75839;
  assign n75745 = n75839 & n75841;
  assign n75877 = n75879 & n75880;
  assign n75846 = ~n75895;
  assign n75893 = n75753 & n115;
  assign n75887 = ~n75753;
  assign n75914 = n72320 & n73581;
  assign n75850 = n75926 & n75927;
  assign n75886 = ~n75929;
  assign n75930 = n75963 & n75964;
  assign n75727 = n131 ^ n75767;
  assign n75760 = n75768 & n130;
  assign n75733 = ~n75769;
  assign n71663 = n75772 ^ n72844;
  assign n75741 = n75779 & n75780;
  assign n75742 = n75783 & n75784;
  assign n75773 = n75772 & n72880;
  assign n75790 = n75800 & n75801;
  assign n75804 = n75816 & n75817;
  assign n75845 = ~n75877;
  assign n75883 = n75887 & n14061;
  assign n75709 = ~n75893;
  assign n75885 = ~n75914;
  assign n75891 = n75930 ^ n73466;
  assign n75924 = ~n75930;
  assign n74036 = n75726 ^ n75727;
  assign n75702 = n75741 ^ n75742;
  assign n75747 = n75742 & n75757;
  assign n75731 = ~n75727;
  assign n75699 = ~n75760;
  assign n75750 = ~n75742;
  assign n71700 = ~n71663;
  assign n75725 = ~n75741;
  assign n75713 = ~n75773;
  assign n75770 = ~n75790;
  assign n75777 = ~n75804;
  assign n75807 = n75845 & n75846;
  assign n75744 = ~n75883;
  assign n75851 = n75885 & n75886;
  assign n72146 = n75891 ^ n75892;
  assign n75913 = n75924 & n75925;
  assign n75669 = n75702 ^ n75703;
  assign n75433 = ~n74036;
  assign n75660 = n75731 & n75732;
  assign n75724 = ~n75747;
  assign n75737 = n71700 & n74103;
  assign n75730 = n75750 & n75703;
  assign n75735 = n75770 & n75771;
  assign n75749 = n75777 & n75778;
  assign n75782 = n75807 ^ n75808;
  assign n75813 = ~n75807;
  assign n75637 = n75850 ^ n75851;
  assign n75857 = n72146 & n74729;
  assign n75859 = n72146 & n75865;
  assign n72259 = ~n72146;
  assign n75852 = ~n75851;
  assign n75888 = ~n75913;
  assign n75675 = n75669 & n129;
  assign n75680 = ~n75669;
  assign n75666 = ~n75660;
  assign n75706 = n75724 & n75725;
  assign n75685 = ~n75730;
  assign n75696 = n75735 ^ n75736;
  assign n75712 = ~n75737;
  assign n75711 = n75749 ^ n72799;
  assign n75734 = ~n75735;
  assign n75740 = n75749 & n72808;
  assign n75738 = ~n75749;
  assign n75746 = n116 ^ n75782;
  assign n75794 = n75813 & n75814;
  assign n75826 = n75637 & n14006;
  assign n75824 = ~n75637;
  assign n75786 = n75852 & n75850;
  assign n75840 = n72259 & n74872;
  assign n75821 = ~n75857;
  assign n75849 = n72259 & n73466;
  assign n74869 = ~n75859;
  assign n75853 = n75888 & n75889;
  assign n75606 = ~n75675;
  assign n75662 = n75680 & n6214;
  assign n75661 = n130 ^ n75696;
  assign n75684 = ~n75706;
  assign n71608 = n75710 ^ n75711;
  assign n75653 = n75712 & n75713;
  assign n75718 = n75733 & n75734;
  assign n75728 = n75738 & n72799;
  assign n75723 = ~n75740;
  assign n75614 = n75745 ^ n75746;
  assign n75751 = ~n75746;
  assign n75775 = ~n75794;
  assign n75806 = n75824 & n114;
  assign n75672 = ~n75826;
  assign n74848 = ~n75840;
  assign n75820 = ~n75849;
  assign n75793 = ~n75786;
  assign n75818 = n75853 ^ n73408;
  assign n75854 = ~n75853;
  assign n73999 = n75660 ^ n75661;
  assign n75634 = ~n75662;
  assign n75670 = n71608 & n75682;
  assign n75678 = n75653 & n75683;
  assign n75652 = n75684 & n75685;
  assign n75665 = ~n75661;
  assign n75679 = n71608 & n74067;
  assign n71610 = ~n71608;
  assign n75681 = ~n75653;
  assign n75698 = ~n75718;
  assign n75704 = n75614 & n72747;
  assign n75701 = n75723 & n75710;
  assign n75692 = ~n75728;
  assign n75707 = ~n75614;
  assign n75673 = n75751 & n75745;
  assign n75752 = n75775 & n75776;
  assign n75631 = ~n75806;
  assign n72075 = n75818 ^ n75819;
  assign n75785 = n75820 & n75821;
  assign n75844 = n75854 & n75855;
  assign n75348 = ~n73999;
  assign n75626 = n75652 ^ n75653;
  assign n75600 = n75665 & n75666;
  assign n74161 = ~n75670;
  assign n75659 = n71610 & n72799;
  assign n75650 = ~n75678;
  assign n75641 = ~n75679;
  assign n75651 = ~n75652;
  assign n75664 = n75681 & n75627;
  assign n75663 = n71610 & n74143;
  assign n75668 = n75698 & n75699;
  assign n75691 = ~n75701;
  assign n75622 = ~n75704;
  assign n75697 = n75707 & n72749;
  assign n75705 = n75752 ^ n75753;
  assign n75743 = ~n75752;
  assign n75565 = n75785 ^ n75786;
  assign n75719 = n75785 & n75793;
  assign n75787 = n72075 & n74731;
  assign n72193 = ~n72075;
  assign n75822 = ~n75844;
  assign n75576 = n75626 ^ n75627;
  assign n75633 = n75650 & n75651;
  assign n75598 = ~n75600;
  assign n75640 = ~n75659;
  assign n74138 = ~n75663;
  assign n75617 = ~n75664;
  assign n75628 = n75668 ^ n75669;
  assign n75635 = ~n75668;
  assign n75657 = n75691 & n75692;
  assign n75648 = ~n75697;
  assign n75674 = n115 ^ n75705;
  assign n75729 = n75743 & n75744;
  assign n75762 = n75565 & n113;
  assign n75761 = ~n75565;
  assign n75764 = ~n75787;
  assign n75781 = n72193 & n73408;
  assign n75792 = n75822 & n75823;
  assign n75579 = n75576 & n128;
  assign n75578 = ~n75576;
  assign n75601 = n129 ^ n75628;
  assign n75616 = ~n75633;
  assign n75629 = n75634 & n75635;
  assign n75588 = n75640 & n75641;
  assign n75615 = n75657 ^ n72749;
  assign n75647 = ~n75657;
  assign n75542 = n75673 ^ n75674;
  assign n75603 = n75674 & n75673;
  assign n75708 = ~n75729;
  assign n75739 = n75761 & n13964;
  assign n75570 = ~n75762;
  assign n75763 = ~n75781;
  assign n71958 = n75791 ^ n75792;
  assign n75788 = ~n75792;
  assign n75566 = n75578 & n6136;
  assign n75505 = ~n75579;
  assign n73951 = n75600 ^ n75601;
  assign n75607 = n75588 & n75545;
  assign n71524 = n75614 ^ n75615;
  assign n75597 = ~n75601;
  assign n75587 = n75616 & n75617;
  assign n75612 = ~n75588;
  assign n75605 = ~n75629;
  assign n75639 = n75647 & n75648;
  assign n75561 = ~n75542;
  assign n75677 = n75708 & n75709;
  assign n75611 = ~n75739;
  assign n75720 = n75763 & n75764;
  assign n75755 = n71958 & n75766;
  assign n75765 = n71958 & n74712;
  assign n72131 = ~n71958;
  assign n75774 = n75788 & n75789;
  assign n75555 = ~n75566;
  assign n75289 = ~n73951;
  assign n75544 = n75587 ^ n75588;
  assign n75491 = n75597 & n75598;
  assign n75593 = n71524 & n74108;
  assign n75580 = n71524 & n72747;
  assign n75575 = n75605 & n75606;
  assign n75583 = ~n75587;
  assign n75584 = ~n75607;
  assign n75596 = n75612 & n75613;
  assign n71557 = ~n71524;
  assign n75621 = ~n75639;
  assign n75636 = n114 ^ n75677;
  assign n75671 = ~n75677;
  assign n75530 = n75719 ^ n75720;
  assign n75689 = n75720 & n75719;
  assign n74774 = ~n75755;
  assign n75754 = n72131 & n75756;
  assign n75748 = n72131 & n73331;
  assign n75721 = ~n75765;
  assign n75758 = ~n75774;
  assign n75470 = n75544 ^ n75545;
  assign n75539 = n75575 ^ n75576;
  assign n75541 = ~n75580;
  assign n75567 = n71557 & n74051;
  assign n75562 = n75583 & n75584;
  assign n74107 = ~n75593;
  assign n75517 = ~n75491;
  assign n75573 = n71557 & n75595;
  assign n75551 = ~n75596;
  assign n75556 = ~n75575;
  assign n75581 = n75621 & n75622;
  assign n75604 = n75636 ^ n75637;
  assign n75658 = n75671 & n75672;
  assign n75686 = n75530 & n13918;
  assign n75693 = ~n75530;
  assign n75722 = ~n75748;
  assign n74757 = ~n75754;
  assign n75716 = n75758 & n75759;
  assign n75510 = n75470 & n6045;
  assign n75506 = ~n75470;
  assign n75492 = n128 ^ n75539;
  assign n75536 = n75555 & n75556;
  assign n75550 = ~n75562;
  assign n75540 = ~n75567;
  assign n74124 = ~n75573;
  assign n75543 = n75581 ^ n72710;
  assign n75592 = n75581 & n72715;
  assign n75449 = n75603 ^ n75604;
  assign n75582 = ~n75581;
  assign n75609 = ~n75604;
  assign n75630 = ~n75658;
  assign n75535 = ~n75686;
  assign n75676 = n75693 & n112;
  assign n74775 = n74774 & n74757;
  assign n75694 = n75716 ^ n75717;
  assign n75690 = n75721 & n75722;
  assign n75714 = ~n75716;
  assign n73915 = n75491 ^ n75492;
  assign n75497 = n75506 & n143;
  assign n75478 = ~n75510;
  assign n75406 = n75492 & n75517;
  assign n75504 = ~n75536;
  assign n75521 = n75540 & n75541;
  assign n71469 = n75542 ^ n75543;
  assign n75520 = n75550 & n75551;
  assign n75571 = n75582 & n72710;
  assign n75560 = ~n75592;
  assign n75572 = n75449 & n72665;
  assign n75563 = ~n75449;
  assign n75532 = n75609 & n75603;
  assign n75608 = n75630 & n75631;
  assign n75501 = ~n75676;
  assign n75459 = n75689 ^ n75690;
  assign n71926 = n75694 ^ n73257;
  assign n75695 = n75694 & n73426;
  assign n75585 = n75690 & n75689;
  assign n75700 = n75714 & n75715;
  assign n75228 = ~n73915;
  assign n75442 = ~n75497;
  assign n75469 = n75504 & n75505;
  assign n75465 = n75520 ^ n75521;
  assign n75511 = n71469 & n72710;
  assign n75516 = n71469 & n75524;
  assign n75507 = n75521 & n75525;
  assign n71485 = ~n71469;
  assign n75485 = ~n75520;
  assign n75512 = ~n75521;
  assign n75548 = n75560 & n75561;
  assign n75557 = n75563 & n72714;
  assign n75528 = ~n75571;
  assign n75453 = ~n75572;
  assign n75538 = ~n75532;
  assign n75564 = n113 ^ n75608;
  assign n75610 = ~n75608;
  assign n75649 = n71926 & n75667;
  assign n75646 = n75459 & n13893;
  assign n72076 = ~n71926;
  assign n75654 = ~n75459;
  assign n75619 = ~n75695;
  assign n75687 = ~n75700;
  assign n75412 = n75465 ^ n75466;
  assign n75445 = n75469 ^ n75470;
  assign n75479 = ~n75469;
  assign n75484 = ~n75507;
  assign n75503 = n71485 & n73990;
  assign n75475 = ~n75511;
  assign n75490 = n75512 & n75466;
  assign n74071 = ~n75516;
  assign n75502 = n71485 & n74074;
  assign n75527 = ~n75548;
  assign n75483 = ~n75557;
  assign n75533 = n75564 ^ n75565;
  assign n75599 = n75610 & n75611;
  assign n75461 = ~n75646;
  assign n74714 = ~n75649;
  assign n75638 = n72076 & n74657;
  assign n75632 = n75654 & n127;
  assign n75642 = n72076 & n74739;
  assign n75655 = n75687 & n75688;
  assign n75409 = n143 ^ n75445;
  assign n75443 = n75412 & n142;
  assign n75444 = ~n75412;
  assign n75464 = n75478 & n75479;
  assign n75472 = n75484 & n75485;
  assign n75455 = ~n75490;
  assign n74090 = ~n75502;
  assign n75474 = ~n75503;
  assign n75489 = n75527 & n75528;
  assign n75375 = n75532 ^ n75533;
  assign n75537 = ~n75533;
  assign n75569 = ~n75599;
  assign n75430 = ~n75632;
  assign n75618 = ~n75638;
  assign n74733 = ~n75642;
  assign n75623 = n75655 ^ n75656;
  assign n75644 = ~n75655;
  assign n73878 = n75406 ^ n75409;
  assign n75405 = ~n75409;
  assign n75367 = ~n75443;
  assign n75424 = n75444 & n5959;
  assign n75441 = ~n75464;
  assign n75454 = ~n75472;
  assign n75414 = n75474 & n75475;
  assign n75450 = n75489 ^ n72665;
  assign n75482 = ~n75489;
  assign n75494 = n75375 & n72634;
  assign n75498 = ~n75375;
  assign n75456 = n75537 & n75538;
  assign n75529 = n75569 & n75570;
  assign n75586 = n75618 & n75619;
  assign n71849 = n75623 ^ n73228;
  assign n75620 = n75623 & n73228;
  assign n75643 = n75644 & n75645;
  assign n75143 = ~n73878;
  assign n75342 = n75405 & n75406;
  assign n75404 = ~n75424;
  assign n75411 = n75441 & n75442;
  assign n71407 = n75449 ^ n75450;
  assign n75447 = n75414 & n75451;
  assign n75413 = n75454 & n75455;
  assign n75434 = ~n75414;
  assign n75468 = n75482 & n75483;
  assign n75378 = ~n75494;
  assign n75488 = n75498 & n72638;
  assign n75463 = ~n75456;
  assign n75499 = n75529 ^ n75530;
  assign n75534 = ~n75529;
  assign n75389 = n75585 ^ n75586;
  assign n75522 = n75586 & n75585;
  assign n75577 = n71849 & n75602;
  assign n75594 = n71849 & n74618;
  assign n71986 = ~n71849;
  assign n75559 = ~n75620;
  assign n75624 = ~n75643;
  assign n75374 = n75411 ^ n75412;
  assign n75386 = n75413 ^ n75414;
  assign n75422 = n71407 & n73936;
  assign n75403 = ~n75411;
  assign n75419 = n71407 & n75433;
  assign n75426 = n75434 & n75387;
  assign n75421 = ~n75413;
  assign n71434 = ~n71407;
  assign n75420 = ~n75447;
  assign n75452 = ~n75468;
  assign n75417 = ~n75488;
  assign n75457 = n112 ^ n75499;
  assign n75526 = n75534 & n75535;
  assign n75549 = n75389 & n13832;
  assign n75552 = ~n75389;
  assign n74696 = ~n75577;
  assign n75568 = n71986 & n74679;
  assign n75558 = ~n75594;
  assign n75591 = n75624 & n75625;
  assign n75343 = n142 ^ n75374;
  assign n75329 = n75386 ^ n75387;
  assign n75392 = n75403 & n75404;
  assign n75400 = n71434 & n74036;
  assign n74054 = ~n75419;
  assign n75408 = n71434 & n72665;
  assign n75410 = n75420 & n75421;
  assign n75382 = ~n75422;
  assign n75385 = ~n75426;
  assign n75415 = n75452 & n75453;
  assign n75306 = n75456 ^ n75457;
  assign n75462 = ~n75457;
  assign n75500 = ~n75526;
  assign n75391 = ~n75549;
  assign n75531 = n75552 & n126;
  assign n75523 = n75558 & n75559;
  assign n74675 = ~n75568;
  assign n75553 = n75591 ^ n73171;
  assign n75589 = ~n75591;
  assign n75104 = n75342 ^ n75343;
  assign n75269 = n75343 & n75342;
  assign n75347 = n75329 & n141;
  assign n75358 = ~n75329;
  assign n75366 = ~n75392;
  assign n74035 = ~n75400;
  assign n75381 = ~n75408;
  assign n75384 = ~n75410;
  assign n75376 = n75415 ^ n72634;
  assign n75431 = n75306 & n72581;
  assign n75416 = ~n75415;
  assign n75423 = ~n75306;
  assign n75394 = n75462 & n75463;
  assign n75458 = n75500 & n75501;
  assign n75327 = n75522 ^ n75523;
  assign n75438 = n75523 & n75522;
  assign n75363 = ~n75531;
  assign n71773 = n75553 ^ n75554;
  assign n75574 = n75589 & n75590;
  assign n75092 = ~n75104;
  assign n75272 = ~n75347;
  assign n75340 = n75358 & n5852;
  assign n75328 = n75366 & n75367;
  assign n71368 = n75375 ^ n75376;
  assign n75354 = n75381 & n75382;
  assign n75355 = n75384 & n75385;
  assign n75407 = n75416 & n75417;
  assign n75418 = n75423 & n72609;
  assign n75345 = ~n75431;
  assign n75428 = n75458 ^ n75459;
  assign n75460 = ~n75458;
  assign n75487 = n75327 & n13776;
  assign n75486 = ~n75327;
  assign n75508 = n71773 & n74636;
  assign n75509 = n71773 & n74577;
  assign n71912 = ~n71773;
  assign n75546 = ~n75574;
  assign n75297 = n75328 ^ n75329;
  assign n75309 = ~n75340;
  assign n75304 = n75354 ^ n75355;
  assign n75346 = n75355 & n75303;
  assign n75352 = n71368 & n73938;
  assign n75310 = ~n75328;
  assign n75353 = n71368 & n73999;
  assign n71372 = ~n71368;
  assign n75320 = ~n75354;
  assign n75356 = ~n75355;
  assign n75377 = ~n75407;
  assign n75313 = ~n75418;
  assign n75395 = n127 ^ n75428;
  assign n75448 = n75460 & n75461;
  assign n75473 = n75486 & n125;
  assign n75324 = ~n75487;
  assign n74655 = ~n75508;
  assign n75493 = n71912 & n73171;
  assign n75480 = ~n75509;
  assign n75496 = n71912 & n75513;
  assign n75514 = n75546 & n75547;
  assign n75270 = n141 ^ n75297;
  assign n75243 = n75303 ^ n75304;
  assign n75298 = n75309 & n75310;
  assign n75319 = ~n75346;
  assign n75336 = n71372 & n72634;
  assign n75331 = n71372 & n75348;
  assign n75316 = ~n75352;
  assign n74018 = ~n75353;
  assign n75330 = n75356 & n75357;
  assign n75349 = n75377 & n75378;
  assign n75236 = n75394 ^ n75395;
  assign n75393 = ~n75395;
  assign n75429 = ~n75448;
  assign n75295 = ~n75473;
  assign n75481 = ~n75493;
  assign n74639 = ~n75496;
  assign n75467 = n75514 ^ n75515;
  assign n75518 = ~n75514;
  assign n73807 = n75269 ^ n75270;
  assign n75182 = n75270 & n75269;
  assign n75284 = n75243 & n5747;
  assign n75285 = ~n75243;
  assign n75271 = ~n75298;
  assign n75311 = n75319 & n75320;
  assign n75292 = ~n75330;
  assign n74002 = ~n75331;
  assign n75317 = ~n75336;
  assign n75307 = n75349 ^ n72581;
  assign n75344 = ~n75349;
  assign n75321 = n75393 & n75394;
  assign n75388 = n75429 & n75430;
  assign n71696 = n73117 ^ n75467;
  assign n75437 = n75480 & n75481;
  assign n75471 = n75467 & n73111;
  assign n75495 = n75518 & n75519;
  assign n75040 = ~n73807;
  assign n75242 = n75271 & n75272;
  assign n75245 = ~n75284;
  assign n75261 = n75285 & n140;
  assign n71316 = n75306 ^ n75307;
  assign n75291 = ~n75311;
  assign n75249 = n75316 & n75317;
  assign n75335 = n75344 & n75345;
  assign n75332 = ~n75321;
  assign n75360 = n75388 ^ n75389;
  assign n75390 = ~n75388;
  assign n75253 = n75437 ^ n75438;
  assign n75372 = n75437 & n75438;
  assign n75446 = n71696 & n74596;
  assign n71846 = ~n71696;
  assign n75397 = ~n75471;
  assign n75476 = ~n75495;
  assign n75210 = n75242 ^ n75243;
  assign n75217 = ~n75261;
  assign n75246 = ~n75242;
  assign n75283 = n75249 & n75225;
  assign n75278 = n71316 & n75289;
  assign n75248 = n75291 & n75292;
  assign n75279 = n71316 & n73895;
  assign n71343 = ~n71316;
  assign n75274 = ~n75249;
  assign n75312 = ~n75335;
  assign n75322 = n126 ^ n75360;
  assign n75383 = n75390 & n75391;
  assign n75231 = ~n75253;
  assign n75427 = n71846 & n74474;
  assign n75370 = ~n75372;
  assign n75432 = n71846 & n75439;
  assign n74593 = ~n75446;
  assign n75440 = n75476 & n75477;
  assign n75183 = n140 ^ n75210;
  assign n75229 = n75245 & n75246;
  assign n75224 = n75248 ^ n75249;
  assign n75256 = ~n75248;
  assign n75259 = n71343 & n72609;
  assign n75265 = n75274 & n75275;
  assign n73980 = ~n75278;
  assign n75238 = ~n75279;
  assign n75264 = n71343 & n73951;
  assign n75255 = ~n75283;
  assign n75280 = n75312 & n75313;
  assign n75160 = n75321 ^ n75322;
  assign n75257 = n75322 & n75332;
  assign n75362 = ~n75383;
  assign n75396 = ~n75427;
  assign n74621 = ~n75432;
  assign n75399 = n75440 ^ n73033;
  assign n75435 = ~n75440;
  assign n73752 = n75182 ^ n75183;
  assign n75185 = ~n75183;
  assign n75187 = n75224 ^ n75225;
  assign n75216 = ~n75229;
  assign n75240 = n75255 & n75256;
  assign n75239 = ~n75259;
  assign n73954 = ~n75264;
  assign n75220 = ~n75265;
  assign n75237 = n75280 ^ n72544;
  assign n75286 = n75280 & n72553;
  assign n75288 = n75160 & n72557;
  assign n75273 = ~n75280;
  assign n75287 = ~n75160;
  assign n75326 = n75362 & n75363;
  assign n75373 = n75396 & n75397;
  assign n71606 = n75398 ^ n75399;
  assign n75425 = n75435 & n75436;
  assign n74996 = ~n73752;
  assign n75132 = n75185 & n75182;
  assign n75190 = n75187 & n5694;
  assign n75198 = ~n75187;
  assign n75186 = n75216 & n75217;
  assign n71269 = n75236 ^ n75237;
  assign n75197 = n75238 & n75239;
  assign n75219 = ~n75240;
  assign n75260 = n75273 & n72544;
  assign n75250 = ~n75286;
  assign n75277 = n75287 & n72496;
  assign n75189 = ~n75288;
  assign n75296 = n75326 ^ n75327;
  assign n75323 = ~n75326;
  assign n75175 = n75372 ^ n75373;
  assign n75368 = n71606 & n73210;
  assign n75371 = n71606 & n75380;
  assign n75369 = ~n75373;
  assign n71774 = ~n71606;
  assign n75401 = ~n75425;
  assign n75151 = ~n75132;
  assign n75159 = n75186 ^ n75187;
  assign n75172 = ~n75190;
  assign n75180 = n75198 & n139;
  assign n75173 = ~n75186;
  assign n75196 = n75219 & n75220;
  assign n75212 = n71269 & n73810;
  assign n75211 = n75197 & n75163;
  assign n75207 = n71269 & n75228;
  assign n75214 = ~n75197;
  assign n71271 = ~n71269;
  assign n75244 = n75250 & n75236;
  assign n75222 = ~n75260;
  assign n75171 = ~n75277;
  assign n75258 = n125 ^ n75296;
  assign n75308 = n75323 & n75324;
  assign n75337 = n75175 & n123;
  assign n75341 = ~n75175;
  assign n75333 = ~n75368;
  assign n75361 = n71774 & n74488;
  assign n75300 = n75369 & n75370;
  assign n74554 = ~n75371;
  assign n75359 = n71774 & n74551;
  assign n75365 = n75401 & n75402;
  assign n75133 = n139 ^ n75159;
  assign n75169 = n75172 & n75173;
  assign n75157 = ~n75180;
  assign n75162 = n75196 ^ n75197;
  assign n73941 = ~n75207;
  assign n75204 = n71271 & n73915;
  assign n75202 = n71271 & n72544;
  assign n75193 = ~n75211;
  assign n75192 = ~n75196;
  assign n75179 = ~n75212;
  assign n75203 = n75214 & n75215;
  assign n75221 = ~n75244;
  assign n75109 = n75257 ^ n75258;
  assign n75194 = n75258 & n75257;
  assign n75294 = ~n75308;
  assign n75153 = ~n75337;
  assign n75325 = n75341 & n13696;
  assign n74579 = ~n75359;
  assign n75334 = ~n75361;
  assign n75305 = ~n75300;
  assign n75338 = n75365 ^ n72974;
  assign n75364 = n75365 & n75379;
  assign n73706 = n75132 ^ n75133;
  assign n75080 = n75133 & n75151;
  assign n75131 = n75162 ^ n75163;
  assign n75156 = ~n75169;
  assign n75181 = n75192 & n75193;
  assign n75178 = ~n75202;
  assign n75168 = ~n75203;
  assign n73914 = ~n75204;
  assign n75199 = n75221 & n75222;
  assign n75223 = n75109 & n72459;
  assign n75227 = ~n75109;
  assign n75252 = n75294 & n75295;
  assign n75177 = ~n75325;
  assign n75299 = n75333 & n75334;
  assign n71553 = n75338 ^ n75339;
  assign n75350 = ~n75364;
  assign n74949 = ~n73706;
  assign n75141 = n75131 & n5626;
  assign n75130 = n75156 & n75157;
  assign n75147 = ~n75131;
  assign n75111 = n75178 & n75179;
  assign n75167 = ~n75181;
  assign n75161 = n75199 ^ n72496;
  assign n75188 = ~n75199;
  assign n75118 = ~n75223;
  assign n75213 = n75227 & n72467;
  assign n75226 = n75252 ^ n75253;
  assign n75251 = n75252 & n13745;
  assign n75247 = ~n75252;
  assign n75127 = n75299 ^ n75300;
  assign n75232 = n75299 & n75305;
  assign n75301 = n71553 & n72974;
  assign n75302 = n71553 & n75318;
  assign n71692 = ~n71553;
  assign n75314 = n75350 & n75351;
  assign n75103 = n75130 ^ n75131;
  assign n75123 = ~n75141;
  assign n75124 = ~n75130;
  assign n75134 = n75147 & n138;
  assign n71200 = n75160 ^ n75161;
  assign n75142 = n75167 & n75168;
  assign n75129 = ~n75111;
  assign n75184 = n75188 & n75189;
  assign n75146 = ~n75213;
  assign n75195 = n124 ^ n75226;
  assign n75241 = n75247 & n124;
  assign n75230 = ~n75251;
  assign n75263 = n75127 & n122;
  assign n75262 = ~n75127;
  assign n75293 = n71692 & n74511;
  assign n75290 = n71692 & n74448;
  assign n75268 = ~n75301;
  assign n74516 = ~n75302;
  assign n71657 = n75314 ^ n75315;
  assign n75081 = n138 ^ n75103;
  assign n75115 = n75123 & n75124;
  assign n75100 = ~n75134;
  assign n75112 = n75142 ^ n75140;
  assign n75150 = n71200 & n72496;
  assign n75148 = n71200 & n73878;
  assign n75149 = n75142 & n75154;
  assign n75139 = ~n75142;
  assign n71259 = ~n71200;
  assign n75170 = ~n75184;
  assign n75090 = n75194 ^ n75195;
  assign n75122 = n75195 & n75194;
  assign n75218 = n75230 & n75231;
  assign n75206 = ~n75241;
  assign n75254 = n75262 & n13622;
  assign n75106 = ~n75263;
  assign n74492 = n75281 ^ n71657;
  assign n75282 = n71657 & n74423;
  assign n75267 = ~n75290;
  assign n74532 = ~n75293;
  assign n75276 = ~n71657;
  assign n73679 = n75080 ^ n75081;
  assign n75021 = n75081 & n75080;
  assign n75057 = n75111 ^ n75112;
  assign n75099 = ~n75115;
  assign n75137 = n75139 & n75140;
  assign n75136 = n71259 & n73761;
  assign n75138 = n71259 & n75143;
  assign n73881 = ~n75148;
  assign n75128 = ~n75149;
  assign n75114 = ~n75150;
  assign n75144 = n75170 & n75171;
  assign n75164 = n75090 & n72387;
  assign n75166 = ~n75090;
  assign n75205 = ~n75218;
  assign n75120 = ~n75254;
  assign n75233 = n75267 & n75268;
  assign n75266 = n75276 & n73123;
  assign n75235 = ~n75282;
  assign n74917 = ~n73679;
  assign n75085 = n75099 & n75100;
  assign n75116 = n75128 & n75129;
  assign n75113 = ~n75136;
  assign n75102 = ~n75137;
  assign n73905 = ~n75138;
  assign n75110 = n75144 ^ n72459;
  assign n75145 = ~n75144;
  assign n75062 = ~n75164;
  assign n75158 = n75166 & n72487;
  assign n75174 = n75205 & n75206;
  assign n75084 = n75232 ^ n75233;
  assign n75209 = n75233 & n75232;
  assign n75234 = ~n75266;
  assign n75048 = n75085 ^ n75057;
  assign n75071 = n75085 & n5602;
  assign n75082 = ~n75085;
  assign n71127 = n75109 ^ n75110;
  assign n75075 = n75113 & n75114;
  assign n75101 = ~n75116;
  assign n75135 = n75145 & n75146;
  assign n75094 = ~n75158;
  assign n75155 = n75174 ^ n75175;
  assign n75176 = ~n75174;
  assign n75201 = n75084 & n13583;
  assign n75200 = ~n75084;
  assign n75208 = n75234 & n75235;
  assign n75026 = n137 ^ n75048;
  assign n75056 = ~n75071;
  assign n75064 = n75082 & n137;
  assign n75076 = n75101 & n75102;
  assign n75096 = n71127 & n73701;
  assign n75095 = n71127 & n75104;
  assign n71204 = ~n71127;
  assign n75059 = ~n75075;
  assign n75117 = ~n75135;
  assign n75125 = n123 ^ n75155;
  assign n75165 = n75176 & n75177;
  assign n75191 = n75200 & n121;
  assign n75073 = ~n75201;
  assign n75019 = n75208 ^ n75209;
  assign n73633 = n75021 ^ n75026;
  assign n75020 = ~n75026;
  assign n75049 = n75056 & n75057;
  assign n75033 = ~n75064;
  assign n75045 = n75075 ^ n75076;
  assign n75079 = n75076 & n75046;
  assign n75077 = ~n75076;
  assign n75088 = n71204 & n75092;
  assign n75087 = n71204 & n72459;
  assign n73857 = ~n75095;
  assign n75065 = ~n75096;
  assign n75089 = n75117 & n75118;
  assign n75016 = n75122 ^ n75125;
  assign n75121 = ~n75125;
  assign n75152 = ~n75165;
  assign n75053 = ~n75191;
  assign n74874 = ~n73633;
  assign n74964 = n75020 & n75021;
  assign n75006 = n75045 ^ n75046;
  assign n75032 = ~n75049;
  assign n75068 = n75077 & n75078;
  assign n75058 = ~n75079;
  assign n75066 = ~n75087;
  assign n73841 = ~n75088;
  assign n75067 = n75089 ^ n75090;
  assign n75107 = n75016 & n72450;
  assign n75093 = ~n75089;
  assign n75098 = ~n75016;
  assign n75070 = n75121 & n75122;
  assign n75126 = n75152 & n75153;
  assign n75005 = n75032 & n75033;
  assign n74989 = ~n75006;
  assign n75055 = n75058 & n75059;
  assign n73866 = n73857 & n73841;
  assign n75013 = n75065 & n75066;
  assign n71100 = n72387 ^ n75067;
  assign n75030 = ~n75068;
  assign n75063 = n75067 & n72387;
  assign n75086 = n75093 & n75094;
  assign n75091 = n75098 & n72364;
  assign n75044 = ~n75107;
  assign n75097 = n75126 ^ n75127;
  assign n75119 = ~n75126;
  assign n74980 = n75005 ^ n75006;
  assign n75011 = n75005 & n5544;
  assign n75010 = ~n75005;
  assign n75041 = n71100 & n73807;
  assign n75039 = n75013 & n75050;
  assign n75037 = n71100 & n73744;
  assign n75029 = ~n75055;
  assign n71098 = ~n71100;
  assign n75042 = ~n75013;
  assign n75025 = ~n75063;
  assign n75061 = ~n75086;
  assign n75015 = ~n75091;
  assign n75074 = n122 ^ n75097;
  assign n75108 = n75119 & n75120;
  assign n74965 = n136 ^ n74980;
  assign n75002 = n75010 & n136;
  assign n74988 = ~n75011;
  assign n75012 = n75029 & n75030;
  assign n75024 = ~n75037;
  assign n75008 = ~n75039;
  assign n75031 = n71098 & n75040;
  assign n73822 = ~n75041;
  assign n75035 = n75042 & n74986;
  assign n75036 = n75061 & n75062;
  assign n74969 = n75070 ^ n75074;
  assign n75069 = ~n75074;
  assign n75105 = ~n75108;
  assign n73598 = n74964 ^ n74965;
  assign n74909 = n74965 & n74964;
  assign n74987 = n74988 & n74989;
  assign n74976 = ~n75002;
  assign n74985 = n75012 ^ n75013;
  assign n74943 = n75024 & n75025;
  assign n75007 = ~n75012;
  assign n73786 = ~n75031;
  assign n74982 = ~n75035;
  assign n75017 = n75036 ^ n72364;
  assign n75047 = n74969 & n72316;
  assign n75043 = ~n75036;
  assign n75051 = ~n74969;
  assign n75027 = n75069 & n75070;
  assign n75083 = n75105 & n75106;
  assign n74824 = ~n73598;
  assign n74951 = n74985 ^ n74986;
  assign n74975 = ~n74987;
  assign n75004 = n75007 & n75008;
  assign n75001 = n74943 & n75009;
  assign n74999 = ~n74943;
  assign n70999 = n75016 ^ n75017;
  assign n75034 = n75043 & n75044;
  assign n74993 = ~n75047;
  assign n75038 = n75051 & n72403;
  assign n75023 = ~n75027;
  assign n75054 = n75083 ^ n75084;
  assign n75072 = ~n75083;
  assign n74968 = n74951 & n151;
  assign n74950 = n74975 & n74976;
  assign n74961 = ~n74951;
  assign n74990 = n74999 & n74963;
  assign n74991 = n70999 & n73752;
  assign n74997 = n70999 & n72364;
  assign n74967 = ~n75001;
  assign n74981 = ~n75004;
  assign n71018 = ~n70999;
  assign n75014 = ~n75034;
  assign n74974 = ~n75038;
  assign n75028 = n121 ^ n75054;
  assign n75060 = n75072 & n75073;
  assign n74933 = n74950 ^ n74951;
  assign n74958 = n74961 & n5509;
  assign n74938 = ~n74950;
  assign n74920 = ~n74968;
  assign n74962 = n74981 & n74982;
  assign n74983 = n71018 & n73626;
  assign n74936 = ~n74990;
  assign n73755 = ~n74991;
  assign n74984 = n71018 & n74996;
  assign n74972 = ~n74997;
  assign n74994 = n75014 & n75015;
  assign n74929 = n75027 ^ n75028;
  assign n75022 = ~n75028;
  assign n75052 = ~n75060;
  assign n74914 = n151 ^ n74933;
  assign n74939 = ~n74958;
  assign n74944 = n74962 ^ n74963;
  assign n74966 = ~n74962;
  assign n74971 = ~n74983;
  assign n73769 = ~n74984;
  assign n74970 = n74994 ^ n72316;
  assign n74998 = n74929 & n72268;
  assign n74992 = ~n74994;
  assign n75000 = ~n74929;
  assign n74977 = n75022 & n75023;
  assign n75018 = n75052 & n75053;
  assign n73574 = n74909 ^ n74914;
  assign n74908 = ~n74914;
  assign n74934 = n74938 & n74939;
  assign n74902 = n74943 ^ n74944;
  assign n74959 = n74966 & n74967;
  assign n70908 = n74969 ^ n74970;
  assign n74922 = n74971 & n74972;
  assign n74979 = n74992 & n74993;
  assign n74948 = ~n74998;
  assign n74995 = n75000 & n72359;
  assign n75003 = n75018 ^ n75019;
  assign n74767 = ~n73574;
  assign n74862 = n74908 & n74909;
  assign n74923 = n74902 & n150;
  assign n74924 = ~n74902;
  assign n74919 = ~n74934;
  assign n74946 = n74922 & n74956;
  assign n74945 = n70908 & n73706;
  assign n74935 = ~n74959;
  assign n74952 = n70908 & n73660;
  assign n74955 = ~n74922;
  assign n71005 = ~n70908;
  assign n74973 = ~n74979;
  assign n74932 = ~n74995;
  assign n74978 = n120 ^ n75003;
  assign n74901 = n74919 & n74920;
  assign n74884 = ~n74923;
  assign n74915 = n74924 & n5464;
  assign n74921 = n74935 & n74936;
  assign n73737 = ~n74945;
  assign n74926 = ~n74946;
  assign n74942 = n71005 & n72403;
  assign n74941 = n71005 & n74949;
  assign n74927 = ~n74952;
  assign n74937 = n74955 & n74899;
  assign n74953 = n74973 & n74974;
  assign n74888 = n74977 ^ n74978;
  assign n74885 = n74901 ^ n74902;
  assign n74904 = ~n74915;
  assign n74903 = ~n74901;
  assign n74898 = n74921 ^ n74922;
  assign n74925 = ~n74921;
  assign n74895 = ~n74937;
  assign n73719 = ~n74941;
  assign n74928 = ~n74942;
  assign n74930 = n74953 ^ n72268;
  assign n74947 = ~n74953;
  assign n74960 = n74888 & n72217;
  assign n74957 = ~n74888;
  assign n74864 = n150 ^ n74885;
  assign n74867 = n74898 ^ n74899;
  assign n74892 = n74903 & n74904;
  assign n74918 = n74925 & n74926;
  assign n74878 = n74927 & n74928;
  assign n70833 = n74929 ^ n74930;
  assign n74940 = n74947 & n74948;
  assign n74954 = n74957 & n72320;
  assign n74913 = ~n74960;
  assign n73538 = n74862 ^ n74864;
  assign n74861 = ~n74864;
  assign n74882 = n74867 & n149;
  assign n74883 = ~n74892;
  assign n74881 = ~n74867;
  assign n74906 = n74878 & n74916;
  assign n74907 = n70833 & n74917;
  assign n74911 = n70833 & n73552;
  assign n74894 = ~n74918;
  assign n70941 = ~n70833;
  assign n74910 = ~n74878;
  assign n74931 = ~n74940;
  assign n74891 = ~n74954;
  assign n74755 = ~n73538;
  assign n74822 = n74861 & n74862;
  assign n74875 = n74881 & n5423;
  assign n74844 = ~n74882;
  assign n74866 = n74883 & n74884;
  assign n74877 = n74894 & n74895;
  assign n74896 = n70941 & n72359;
  assign n74880 = ~n74906;
  assign n73693 = ~n74907;
  assign n74900 = n74910 & n74857;
  assign n74897 = n70941 & n73679;
  assign n74887 = ~n74911;
  assign n74905 = n74931 & n74932;
  assign n74831 = ~n74822;
  assign n74840 = n74866 ^ n74867;
  assign n74854 = ~n74866;
  assign n74855 = ~n74875;
  assign n74856 = n74877 ^ n74878;
  assign n74879 = ~n74877;
  assign n74886 = ~n74896;
  assign n73675 = ~n74897;
  assign n74860 = ~n74900;
  assign n74889 = n74905 ^ n72217;
  assign n74912 = ~n74905;
  assign n74823 = n149 ^ n74840;
  assign n74853 = n74854 & n74855;
  assign n74821 = n74856 ^ n74857;
  assign n74876 = n74879 & n74880;
  assign n74811 = n74886 & n74887;
  assign n70760 = n74888 ^ n74889;
  assign n74893 = n74912 & n74913;
  assign n73478 = n74822 ^ n74823;
  assign n74781 = n74823 & n74831;
  assign n74842 = n74821 & n148;
  assign n74841 = ~n74821;
  assign n74843 = ~n74853;
  assign n74873 = n70760 & n73581;
  assign n74870 = n70760 & n73633;
  assign n74859 = ~n74876;
  assign n70859 = ~n70760;
  assign n74826 = ~n74811;
  assign n74890 = ~n74893;
  assign n74697 = ~n73478;
  assign n74836 = n74841 & n5391;
  assign n74802 = ~n74842;
  assign n74820 = n74843 & n74844;
  assign n74837 = n74859 & n74860;
  assign n74858 = n70859 & n72320;
  assign n73654 = ~n74870;
  assign n74851 = ~n74873;
  assign n74865 = n70859 & n74874;
  assign n74871 = n74890 & n74891;
  assign n74800 = n74820 ^ n74821;
  assign n74815 = ~n74820;
  assign n74816 = ~n74836;
  assign n74812 = n74837 ^ n74838;
  assign n74839 = n74837 & n74846;
  assign n74845 = ~n74837;
  assign n74852 = ~n74858;
  assign n73632 = ~n74865;
  assign n74849 = n74871 ^ n74872;
  assign n74868 = ~n74871;
  assign n74782 = n148 ^ n74800;
  assign n74784 = n74811 ^ n74812;
  assign n74810 = n74815 & n74816;
  assign n74825 = ~n74839;
  assign n74834 = n74845 & n74838;
  assign n70682 = n72146 ^ n74849;
  assign n74788 = n74851 & n74852;
  assign n74850 = n74849 & n72259;
  assign n74863 = n74868 & n74869;
  assign n73439 = n74781 ^ n74782;
  assign n74740 = n74782 & n74781;
  assign n74798 = n74784 & n147;
  assign n74799 = ~n74784;
  assign n74801 = ~n74810;
  assign n74818 = n74825 & n74826;
  assign n74805 = ~n74834;
  assign n74828 = n74788 & n74769;
  assign n74829 = n70682 & n73598;
  assign n70800 = ~n70682;
  assign n74832 = ~n74788;
  assign n74807 = ~n74850;
  assign n74847 = ~n74863;
  assign n74664 = ~n73439;
  assign n74762 = ~n74798;
  assign n74797 = n74799 & n5352;
  assign n74783 = n74801 & n74802;
  assign n74804 = ~n74818;
  assign n74813 = n70800 & n74824;
  assign n74793 = ~n74828;
  assign n73597 = ~n74829;
  assign n74814 = n74832 & n74833;
  assign n74817 = n70800 & n73466;
  assign n74835 = n74847 & n74848;
  assign n74760 = n74783 ^ n74784;
  assign n74779 = ~n74783;
  assign n74780 = ~n74797;
  assign n74787 = n74804 & n74805;
  assign n73619 = ~n74813;
  assign n74766 = ~n74814;
  assign n74806 = ~n74817;
  assign n74827 = n74835 & n72075;
  assign n74830 = ~n74835;
  assign n74741 = n147 ^ n74760;
  assign n74777 = n74779 & n74780;
  assign n74768 = n74787 ^ n74788;
  assign n74792 = ~n74787;
  assign n74754 = n74806 & n74807;
  assign n74808 = ~n74827;
  assign n74819 = n74830 & n72193;
  assign n73393 = n74740 ^ n74741;
  assign n74700 = n74741 & n74740;
  assign n74721 = n74768 ^ n74769;
  assign n74761 = ~n74777;
  assign n74778 = n74792 & n74793;
  assign n74789 = n74754 & n74794;
  assign n74786 = ~n74754;
  assign n74803 = n74808 & n74809;
  assign n74796 = ~n74819;
  assign n74616 = ~n73393;
  assign n74751 = n74721 & n5311;
  assign n74744 = n74761 & n74762;
  assign n74752 = ~n74721;
  assign n74765 = ~n74778;
  assign n74785 = n74786 & n74729;
  assign n74749 = ~n74789;
  assign n74795 = ~n74803;
  assign n74790 = n74796 & n74808;
  assign n74720 = n146 ^ n74744;
  assign n74736 = ~n74751;
  assign n74743 = n74752 & n146;
  assign n74737 = ~n74744;
  assign n74753 = n74765 & n74766;
  assign n74727 = ~n74785;
  assign n70594 = n74790 ^ n74791;
  assign n74776 = n74795 & n74796;
  assign n74701 = n74720 ^ n74721;
  assign n74723 = n74736 & n74737;
  assign n74719 = ~n74743;
  assign n74728 = n74753 ^ n74754;
  assign n74748 = ~n74753;
  assign n70479 = n74775 ^ n74776;
  assign n74772 = n70594 & n73408;
  assign n74771 = n70594 & n73574;
  assign n70696 = ~n70594;
  assign n74773 = ~n74776;
  assign n73348 = n74700 ^ n74701;
  assign n74699 = ~n74701;
  assign n74718 = ~n74723;
  assign n74694 = n74728 ^ n74729;
  assign n74742 = n74748 & n74749;
  assign n74758 = n70479 & n73538;
  assign n74759 = n70479 & n73331;
  assign n70656 = ~n70479;
  assign n74763 = n70696 & n72193;
  assign n74764 = n70696 & n74767;
  assign n73577 = ~n74771;
  assign n74745 = ~n74772;
  assign n74770 = n74773 & n74774;
  assign n74580 = ~n73348;
  assign n74661 = n74699 & n74700;
  assign n74709 = n74694 & n145;
  assign n74693 = n74718 & n74719;
  assign n74706 = ~n74694;
  assign n74726 = ~n74742;
  assign n74750 = n70656 & n74755;
  assign n73533 = ~n74758;
  assign n74735 = ~n74759;
  assign n74747 = n70656 & n72131;
  assign n74746 = ~n74763;
  assign n73557 = ~n74764;
  assign n74756 = ~n74770;
  assign n74678 = n74693 ^ n74694;
  assign n74702 = n74706 & n5261;
  assign n74670 = ~n74709;
  assign n74690 = ~n74693;
  assign n74704 = n74726 & n74727;
  assign n74705 = n74745 & n74746;
  assign n74734 = ~n74747;
  assign n73515 = ~n74750;
  assign n74738 = n74756 & n74757;
  assign n74662 = n145 ^ n74678;
  assign n74689 = ~n74702;
  assign n74687 = n74704 ^ n74705;
  assign n74707 = ~n74704;
  assign n74672 = n74734 & n74735;
  assign n74725 = n74705 & n74688;
  assign n74715 = n74738 ^ n74739;
  assign n74730 = ~n74705;
  assign n74732 = ~n74738;
  assign n73299 = n74661 ^ n74662;
  assign n74609 = n74662 & n74661;
  assign n74646 = n74687 ^ n74688;
  assign n74681 = n74689 & n74690;
  assign n70441 = n71926 ^ n74715;
  assign n74717 = n74672 & n74649;
  assign n74711 = ~n74672;
  assign n74708 = ~n74725;
  assign n74722 = n74730 & n74731;
  assign n74716 = ~n74715;
  assign n74724 = n74732 & n74733;
  assign n74539 = ~n73299;
  assign n74619 = ~n74609;
  assign n74668 = n74646 & n5208;
  assign n74673 = ~n74646;
  assign n74669 = ~n74681;
  assign n74691 = n70441 & n73478;
  assign n70460 = ~n70441;
  assign n74698 = n74707 & n74708;
  assign n74710 = n74711 & n74712;
  assign n74703 = n74716 & n71926;
  assign n74667 = ~n74717;
  assign n74686 = ~n74722;
  assign n74713 = ~n74724;
  assign n74642 = ~n74668;
  assign n74645 = n74669 & n74670;
  assign n74665 = n74673 & n144;
  assign n73477 = ~n74691;
  assign n74683 = n70460 & n73426;
  assign n74684 = n70460 & n74697;
  assign n74685 = ~n74698;
  assign n74677 = ~n74703;
  assign n74652 = ~n74710;
  assign n74692 = n74713 & n74714;
  assign n74631 = n74645 ^ n74646;
  assign n74630 = ~n74665;
  assign n74643 = ~n74645;
  assign n74676 = ~n74683;
  assign n73499 = ~n74684;
  assign n74671 = n74685 & n74686;
  assign n74680 = n74692 ^ n71849;
  assign n74695 = ~n74692;
  assign n74610 = n144 ^ n74631;
  assign n74640 = n74642 & n74643;
  assign n74648 = n74671 ^ n74672;
  assign n74626 = n74676 & n74677;
  assign n70296 = n74679 ^ n74680;
  assign n74666 = ~n74671;
  assign n74682 = n74695 & n74696;
  assign n73235 = n74609 ^ n74610;
  assign n74560 = n74610 & n74619;
  assign n74629 = ~n74640;
  assign n74612 = n74648 ^ n74649;
  assign n74653 = n70296 & n71986;
  assign n74660 = n70296 & n74664;
  assign n74658 = n74626 & n74606;
  assign n74656 = ~n74626;
  assign n70489 = ~n70296;
  assign n74663 = n74666 & n74667;
  assign n74674 = ~n74682;
  assign n74496 = ~n73235;
  assign n74569 = ~n74560;
  assign n74611 = n74629 & n74630;
  assign n74633 = n74612 & n5179;
  assign n74632 = ~n74612;
  assign n74647 = n70489 & n73439;
  assign n74635 = ~n74653;
  assign n74644 = n74656 & n74657;
  assign n74650 = n70489 & n73228;
  assign n74628 = ~n74658;
  assign n73444 = ~n74660;
  assign n74651 = ~n74663;
  assign n74659 = n74674 & n74675;
  assign n74585 = n74611 ^ n74612;
  assign n74599 = ~n74611;
  assign n74623 = n74632 & n159;
  assign n74600 = ~n74633;
  assign n74602 = ~n74644;
  assign n73463 = ~n74647;
  assign n74634 = ~n74650;
  assign n74625 = n74651 & n74652;
  assign n74637 = n74659 ^ n71773;
  assign n74654 = ~n74659;
  assign n74561 = n159 ^ n74585;
  assign n74598 = n74599 & n74600;
  assign n74587 = ~n74623;
  assign n74605 = n74625 ^ n74626;
  assign n74584 = n74634 & n74635;
  assign n70249 = n74636 ^ n74637;
  assign n74627 = ~n74625;
  assign n74641 = n74654 & n74655;
  assign n74468 = n74560 ^ n74561;
  assign n74568 = ~n74561;
  assign n74586 = ~n74598;
  assign n74557 = n74605 ^ n74606;
  assign n74622 = n70249 & n73171;
  assign n74614 = n70249 & n73393;
  assign n74613 = n74584 & n74571;
  assign n74617 = ~n74584;
  assign n74624 = n74627 & n74628;
  assign n70257 = ~n70249;
  assign n74638 = ~n74641;
  assign n74522 = n74568 & n74569;
  assign n74556 = n74586 & n74587;
  assign n74591 = n74557 & n5130;
  assign n74588 = ~n74557;
  assign n74590 = ~n74613;
  assign n73420 = ~n74614;
  assign n74608 = n70257 & n74616;
  assign n74603 = n74617 & n74618;
  assign n74604 = n70257 & n71912;
  assign n74595 = ~n74622;
  assign n74601 = ~n74624;
  assign n74615 = n74638 & n74639;
  assign n74534 = ~n74522;
  assign n74546 = n74556 ^ n74557;
  assign n74558 = ~n74556;
  assign n74581 = n74588 & n158;
  assign n74559 = ~n74591;
  assign n74583 = n74601 & n74602;
  assign n74567 = ~n74603;
  assign n74594 = ~n74604;
  assign n73398 = ~n74608;
  assign n74597 = n74615 ^ n71696;
  assign n74620 = ~n74615;
  assign n74523 = n158 ^ n74546;
  assign n74555 = n74558 & n74559;
  assign n74548 = ~n74581;
  assign n74570 = n74583 ^ n74584;
  assign n74543 = n74594 & n74595;
  assign n70158 = n74596 ^ n74597;
  assign n74589 = ~n74583;
  assign n74607 = n74620 & n74621;
  assign n74502 = n74522 ^ n74523;
  assign n74477 = n74523 & n74534;
  assign n74547 = ~n74555;
  assign n74525 = n74570 ^ n74571;
  assign n74573 = n70158 & n74580;
  assign n74574 = n70158 & n73111;
  assign n74575 = n74543 & n74529;
  assign n74576 = ~n74543;
  assign n74582 = n74589 & n74590;
  assign n70298 = ~n70158;
  assign n74592 = ~n74607;
  assign n71288 = n74502 ^ n72331;
  assign n74500 = n74502 & n72331;
  assign n74501 = ~n74502;
  assign n74484 = ~n74477;
  assign n74524 = n74547 & n74548;
  assign n74544 = n74525 & n5088;
  assign n74545 = ~n74525;
  assign n73369 = ~n74573;
  assign n74550 = ~n74574;
  assign n74541 = ~n74575;
  assign n74562 = n74576 & n74577;
  assign n74564 = n70298 & n71696;
  assign n74563 = n70298 & n73348;
  assign n74566 = ~n74582;
  assign n74572 = n74592 & n74593;
  assign n74471 = n71288 & n73382;
  assign n71284 = ~n71288;
  assign n74463 = ~n74500;
  assign n74415 = n74501 & n72331;
  assign n74505 = n74524 ^ n74525;
  assign n74520 = ~n74524;
  assign n74521 = ~n74544;
  assign n74537 = n74545 & n157;
  assign n74527 = ~n74562;
  assign n73345 = ~n74563;
  assign n74549 = ~n74564;
  assign n74542 = n74566 & n74567;
  assign n74552 = n74572 ^ n71606;
  assign n74578 = ~n74572;
  assign n74462 = ~n74471;
  assign n74478 = n157 ^ n74505;
  assign n74517 = n74520 & n74521;
  assign n74509 = ~n74537;
  assign n74528 = n74542 ^ n74543;
  assign n74503 = n74549 & n74550;
  assign n70084 = n74551 ^ n74552;
  assign n74540 = ~n74542;
  assign n74565 = n74578 & n74579;
  assign n74449 = n74462 & n74463;
  assign n74469 = n74477 ^ n74478;
  assign n74483 = ~n74478;
  assign n74508 = ~n74517;
  assign n74481 = n74528 ^ n74529;
  assign n74536 = n70084 & n71606;
  assign n74535 = n70084 & n74539;
  assign n74538 = n74540 & n74541;
  assign n70239 = ~n70084;
  assign n74490 = ~n74503;
  assign n74553 = ~n74565;
  assign n74416 = n74449 ^ n74445;
  assign n74444 = ~n74449;
  assign n74459 = n74469 & n72201;
  assign n74455 = ~n74469;
  assign n74431 = n74483 & n74484;
  assign n74480 = n74508 & n74509;
  assign n74499 = n74481 & n5043;
  assign n74498 = ~n74481;
  assign n74530 = n70239 & n73210;
  assign n74519 = n70239 & n73299;
  assign n73293 = ~n74535;
  assign n74513 = ~n74536;
  assign n74526 = ~n74538;
  assign n74533 = n74553 & n74554;
  assign n72723 = n167 ^ n74416;
  assign n74417 = ~n74416;
  assign n74323 = n74444 & n74445;
  assign n74451 = n74455 & n72191;
  assign n74434 = ~n74459;
  assign n74443 = ~n74431;
  assign n74454 = n74480 ^ n74481;
  assign n74475 = ~n74480;
  assign n74497 = n74498 & n156;
  assign n74476 = ~n74499;
  assign n73318 = ~n74519;
  assign n74504 = n74526 & n74527;
  assign n74514 = ~n74530;
  assign n74512 = n74533 ^ n71553;
  assign n74531 = ~n74533;
  assign n73976 = ~n72723;
  assign n74265 = n74417 & n167;
  assign n74428 = n74434 & n74415;
  assign n74419 = ~n74451;
  assign n74432 = n156 ^ n74454;
  assign n74470 = n74475 & n74476;
  assign n74453 = ~n74497;
  assign n74473 = n74503 ^ n74504;
  assign n74507 = n74504 & n74510;
  assign n70016 = n74511 ^ n74512;
  assign n74440 = n74513 & n74514;
  assign n74506 = ~n74504;
  assign n74518 = n74531 & n74532;
  assign n74418 = ~n74428;
  assign n74380 = n74431 ^ n74432;
  assign n74414 = n74419 & n74434;
  assign n74396 = n74432 & n74443;
  assign n74452 = ~n74470;
  assign n74436 = n74473 ^ n74474;
  assign n74486 = n70016 & n71553;
  assign n74493 = n70016 & n74496;
  assign n74494 = n74440 & n74421;
  assign n74487 = ~n74440;
  assign n70026 = ~n70016;
  assign n74495 = n74506 & n74474;
  assign n74489 = ~n74507;
  assign n74515 = ~n74518;
  assign n71172 = n74414 ^ n74415;
  assign n74399 = n74418 & n74419;
  assign n74409 = n74380 & n72098;
  assign n74413 = ~n74380;
  assign n74400 = ~n74396;
  assign n74435 = n74452 & n74453;
  assign n74457 = n74436 & n155;
  assign n74456 = ~n74436;
  assign n74461 = ~n74486;
  assign n74472 = n74487 & n74488;
  assign n74482 = n74489 & n74490;
  assign n74485 = n70026 & n72974;
  assign n73246 = ~n74493;
  assign n74479 = n70026 & n73235;
  assign n74438 = ~n74494;
  assign n74465 = ~n74495;
  assign n74491 = n74515 & n74516;
  assign n74381 = n74399 ^ n72098;
  assign n74390 = n71172 & n72191;
  assign n71175 = ~n71172;
  assign n74404 = ~n74409;
  assign n74408 = n74413 & n72117;
  assign n74403 = ~n74399;
  assign n74410 = n74435 ^ n74436;
  assign n74429 = ~n74435;
  assign n74450 = n74456 & n5010;
  assign n74412 = ~n74457;
  assign n74425 = ~n74472;
  assign n73262 = ~n74479;
  assign n74464 = ~n74482;
  assign n74460 = ~n74485;
  assign n70079 = n74491 ^ n74492;
  assign n71089 = n74380 ^ n74381;
  assign n74374 = ~n74390;
  assign n74389 = n71175 & n73273;
  assign n74392 = n74403 & n74404;
  assign n74386 = ~n74408;
  assign n74397 = n155 ^ n74410;
  assign n74430 = ~n74450;
  assign n74402 = n74460 & n74461;
  assign n74439 = n74464 & n74465;
  assign n73213 = n74468 ^ n70079;
  assign n74467 = n70079 & n73123;
  assign n74466 = ~n70079;
  assign n74368 = n71089 & n73187;
  assign n71118 = ~n71089;
  assign n74373 = ~n74389;
  assign n74385 = ~n74392;
  assign n74345 = n74396 ^ n74397;
  assign n74355 = n74397 & n74400;
  assign n74426 = n74429 & n74430;
  assign n74420 = n74439 ^ n74440;
  assign n74446 = n74402 & n74379;
  assign n74447 = ~n74402;
  assign n74437 = ~n74439;
  assign n74458 = n74466 & n71657;
  assign n74442 = ~n74467;
  assign n74342 = ~n74368;
  assign n74353 = n71118 & n72117;
  assign n74365 = n74373 & n74374;
  assign n74377 = n74345 & n72025;
  assign n74363 = n74385 & n74386;
  assign n74376 = ~n74345;
  assign n74395 = n74420 ^ n74421;
  assign n74411 = ~n74426;
  assign n74427 = n74437 & n74438;
  assign n74406 = ~n74446;
  assign n74433 = n74447 & n74448;
  assign n74441 = ~n74458;
  assign n74343 = ~n74353;
  assign n74346 = n74363 ^ n72029;
  assign n74361 = n74365 & n74366;
  assign n74358 = ~n74365;
  assign n74370 = n74376 & n72029;
  assign n74338 = ~n74377;
  assign n74356 = ~n74363;
  assign n74407 = n74395 & n4987;
  assign n74394 = n74411 & n74412;
  assign n74398 = ~n74395;
  assign n74424 = ~n74427;
  assign n74383 = ~n74433;
  assign n74422 = n74441 & n74442;
  assign n74284 = n74342 & n74343;
  assign n71030 = n74345 ^ n74346;
  assign n74347 = n74358 & n74359;
  assign n74336 = ~n74361;
  assign n74357 = ~n74370;
  assign n74375 = n74394 ^ n74395;
  assign n74391 = n74398 & n154;
  assign n74387 = ~n74407;
  assign n74388 = ~n74394;
  assign n74341 = n74422 ^ n74423;
  assign n74401 = n74424 & n74425;
  assign n74329 = n71030 & n72025;
  assign n74326 = n74284 & n74305;
  assign n74324 = ~n74284;
  assign n71049 = ~n71030;
  assign n74334 = n74336 & n74323;
  assign n74328 = ~n74347;
  assign n74350 = n74356 & n74357;
  assign n74362 = n154 ^ n74375;
  assign n74384 = n74387 & n74388;
  assign n74372 = ~n74391;
  assign n74378 = n74401 ^ n74402;
  assign n74405 = ~n74401;
  assign n74317 = n74324 & n74325;
  assign n74308 = ~n74326;
  assign n74320 = n71049 & n73104;
  assign n74307 = ~n74329;
  assign n74327 = ~n74334;
  assign n74322 = n74328 & n74336;
  assign n74337 = ~n74350;
  assign n74302 = n74355 ^ n74362;
  assign n74354 = ~n74362;
  assign n74349 = n74378 ^ n74379;
  assign n74371 = ~n74384;
  assign n74393 = n74405 & n74406;
  assign n74290 = ~n74317;
  assign n74306 = ~n74320;
  assign n74310 = n74322 ^ n74323;
  assign n74304 = n74327 & n74328;
  assign n74321 = n74337 & n74338;
  assign n74339 = n74302 & n71934;
  assign n74335 = ~n74302;
  assign n74312 = n74354 & n74355;
  assign n74369 = n74349 & n4946;
  assign n74348 = n74371 & n74372;
  assign n74367 = ~n74349;
  assign n74382 = ~n74393;
  assign n74285 = n74304 ^ n74305;
  assign n74255 = n74306 & n74307;
  assign n74300 = n74310 & n166;
  assign n74299 = ~n74310;
  assign n74309 = ~n74304;
  assign n74303 = n74321 ^ n71928;
  assign n74319 = ~n74321;
  assign n74330 = n74335 & n71928;
  assign n74298 = ~n74339;
  assign n74331 = n74348 ^ n74349;
  assign n74360 = n74367 & n153;
  assign n74352 = ~n74348;
  assign n74351 = ~n74369;
  assign n74364 = n74382 & n74383;
  assign n74249 = n74284 ^ n74285;
  assign n74291 = n74255 & n74270;
  assign n74293 = n74299 & n17578;
  assign n74267 = ~n74300;
  assign n74287 = ~n74255;
  assign n70934 = n74302 ^ n74303;
  assign n74301 = n74308 & n74309;
  assign n74318 = ~n74330;
  assign n74314 = n153 ^ n74331;
  assign n74344 = n74351 & n74352;
  assign n74333 = ~n74360;
  assign n74340 = n152 ^ n74364;
  assign n74275 = n74249 & n17487;
  assign n74272 = ~n74249;
  assign n74282 = n70934 & n71934;
  assign n74280 = n74287 & n74288;
  assign n74274 = ~n74291;
  assign n70953 = ~n70934;
  assign n74283 = ~n74293;
  assign n74289 = ~n74301;
  assign n74260 = n74312 ^ n74314;
  assign n74313 = n74318 & n74319;
  assign n74311 = ~n74314;
  assign n74316 = n74340 ^ n74341;
  assign n74332 = ~n74344;
  assign n74259 = n74272 & n165;
  assign n74250 = ~n74275;
  assign n74254 = ~n74280;
  assign n74279 = n70953 & n73035;
  assign n74263 = ~n74282;
  assign n74264 = n74283 & n74267;
  assign n74276 = n74283 & n74265;
  assign n74269 = n74289 & n74290;
  assign n74292 = n74260 & n71828;
  assign n74294 = ~n74260;
  assign n74295 = n74311 & n74312;
  assign n74297 = ~n74313;
  assign n74315 = n74332 & n74333;
  assign n74233 = ~n74259;
  assign n72666 = n74264 ^ n74265;
  assign n74256 = n74269 ^ n74270;
  assign n74266 = ~n74276;
  assign n74262 = ~n74279;
  assign n74273 = ~n74269;
  assign n74258 = ~n74292;
  assign n74286 = n74294 & n71872;
  assign n74281 = n74297 & n74298;
  assign n74296 = n74315 ^ n74316;
  assign n74217 = n74255 ^ n74256;
  assign n72685 = ~n72666;
  assign n74218 = n74262 & n74263;
  assign n74248 = n74266 & n74267;
  assign n74268 = n74273 & n74274;
  assign n74261 = n74281 ^ n71828;
  assign n74277 = ~n74286;
  assign n74278 = ~n74281;
  assign n74221 = n74295 ^ n74296;
  assign n74241 = n74217 & n17421;
  assign n74234 = n74248 ^ n74249;
  assign n74237 = ~n74217;
  assign n74225 = ~n74218;
  assign n74251 = ~n74248;
  assign n70845 = n74260 ^ n74261;
  assign n74253 = ~n74268;
  assign n74271 = n74277 & n74278;
  assign n74231 = ~n74221;
  assign n74213 = n165 ^ n74234;
  assign n74229 = n74237 & n164;
  assign n74211 = ~n74241;
  assign n74246 = n74250 & n74251;
  assign n74252 = n70845 & n72955;
  assign n74235 = n74253 & n74254;
  assign n70851 = ~n70845;
  assign n74257 = ~n74271;
  assign n72642 = n74213 ^ n72666;
  assign n74181 = n74213 & n72666;
  assign n74200 = ~n74229;
  assign n74219 = n74235 ^ n74236;
  assign n74232 = ~n74246;
  assign n74240 = n74235 & n74247;
  assign n74244 = n70851 & n71828;
  assign n74228 = ~n74252;
  assign n74238 = ~n74235;
  assign n74243 = n74257 & n74258;
  assign n73893 = ~n72642;
  assign n74184 = ~n74181;
  assign n74173 = n74218 ^ n74219;
  assign n74216 = n74232 & n74233;
  assign n74226 = n74238 & n74236;
  assign n74224 = ~n74240;
  assign n74222 = n74243 ^ n71750;
  assign n74227 = ~n74244;
  assign n74242 = n74243 & n71750;
  assign n74245 = ~n74243;
  assign n74203 = n74216 ^ n74217;
  assign n74212 = ~n74216;
  assign n70745 = n74221 ^ n74222;
  assign n74220 = n74224 & n74225;
  assign n74209 = ~n74226;
  assign n74174 = n74227 & n74228;
  assign n74230 = ~n74242;
  assign n74239 = n74245 & n71769;
  assign n74182 = n164 ^ n74203;
  assign n74210 = n74211 & n74212;
  assign n74207 = n70745 & n72900;
  assign n70743 = ~n70745;
  assign n74208 = ~n74220;
  assign n74180 = ~n74174;
  assign n74223 = n74230 & n74231;
  assign n74215 = ~n74239;
  assign n72603 = n74181 ^ n74182;
  assign n74183 = ~n74182;
  assign n74197 = ~n74207;
  assign n74198 = n74208 & n74209;
  assign n74206 = n70743 & n71769;
  assign n74199 = ~n74210;
  assign n74214 = ~n74223;
  assign n73861 = ~n72603;
  assign n74152 = n74183 & n74184;
  assign n74175 = n74198 ^ n74193;
  assign n74185 = n74199 & n74200;
  assign n74194 = n74198 & n74202;
  assign n74196 = ~n74206;
  assign n74192 = ~n74198;
  assign n74205 = n74214 & n74215;
  assign n74132 = n74174 ^ n74175;
  assign n74156 = ~n74152;
  assign n74169 = n74185 ^ n74173;
  assign n74189 = n74185 & n17333;
  assign n74190 = n74192 & n74193;
  assign n74179 = ~n74194;
  assign n74188 = ~n74185;
  assign n74134 = n74196 & n74197;
  assign n74201 = n74205 & n71700;
  assign n74204 = ~n74205;
  assign n74153 = n163 ^ n74169;
  assign n74178 = n74179 & n74180;
  assign n74177 = n74188 & n163;
  assign n74172 = ~n74189;
  assign n74141 = ~n74134;
  assign n74167 = ~n74190;
  assign n74187 = ~n74201;
  assign n74195 = n74204 & n71663;
  assign n73833 = n74152 ^ n74153;
  assign n74155 = ~n74153;
  assign n74168 = n74172 & n74173;
  assign n74163 = ~n74177;
  assign n74166 = ~n74178;
  assign n74186 = n74187 & n74191;
  assign n74171 = ~n74195;
  assign n73843 = ~n73833;
  assign n74111 = n74155 & n74156;
  assign n74150 = n74166 & n74167;
  assign n74162 = ~n74168;
  assign n74170 = ~n74186;
  assign n74176 = n74171 & n74187;
  assign n74117 = ~n74111;
  assign n74135 = n74150 ^ n74151;
  assign n74154 = n74150 & n74151;
  assign n74145 = n74162 & n74163;
  assign n74157 = ~n74150;
  assign n74159 = n74170 & n74171;
  assign n74164 = ~n74176;
  assign n74098 = n74134 ^ n74135;
  assign n74125 = n74145 ^ n74132;
  assign n74139 = n74145 & n17249;
  assign n74142 = ~n74145;
  assign n74140 = ~n74154;
  assign n74148 = n74157 & n74158;
  assign n74144 = n74159 ^ n71608;
  assign n70634 = n74164 ^ n74165;
  assign n74160 = ~n74159;
  assign n74112 = n162 ^ n74125;
  assign n74079 = ~n74098;
  assign n74131 = ~n74139;
  assign n74136 = n74140 & n74141;
  assign n74133 = n74142 & n162;
  assign n70554 = n74143 ^ n74144;
  assign n74127 = ~n74148;
  assign n74147 = n70634 & n71663;
  assign n70684 = ~n70634;
  assign n74149 = n74160 & n74161;
  assign n72526 = n74111 ^ n74112;
  assign n74057 = n74112 & n74117;
  assign n74121 = n70554 & n71610;
  assign n74128 = n74131 & n74132;
  assign n70603 = ~n70554;
  assign n74115 = ~n74133;
  assign n74126 = ~n74136;
  assign n74146 = n70684 & n72880;
  assign n74130 = ~n74147;
  assign n74137 = ~n74149;
  assign n73779 = ~n72526;
  assign n74065 = ~n74057;
  assign n74119 = n70603 & n72799;
  assign n74105 = ~n74121;
  assign n74102 = n74126 & n74127;
  assign n74114 = ~n74128;
  assign n74122 = n74137 & n74138;
  assign n74129 = ~n74146;
  assign n74093 = n74102 ^ n74103;
  assign n74097 = n74114 & n74115;
  assign n74100 = ~n74102;
  assign n74104 = ~n74119;
  assign n74109 = n74122 ^ n71524;
  assign n74092 = n74129 & n74130;
  assign n74123 = ~n74122;
  assign n74045 = n74092 ^ n74093;
  assign n74077 = n74097 ^ n74098;
  assign n74094 = n74097 & n17182;
  assign n74041 = n74104 & n74105;
  assign n74095 = ~n74097;
  assign n70491 = n74108 ^ n74109;
  assign n74113 = n74092 & n74118;
  assign n74116 = ~n74092;
  assign n74120 = n74123 & n74124;
  assign n74073 = n74045 & n160;
  assign n74058 = n161 ^ n74077;
  assign n74072 = ~n74045;
  assign n74078 = ~n74094;
  assign n74086 = n74095 & n161;
  assign n74091 = n74041 & n74096;
  assign n74085 = n70491 & n72747;
  assign n74087 = ~n74041;
  assign n70514 = ~n70491;
  assign n74101 = ~n74113;
  assign n74110 = n74116 & n74103;
  assign n74106 = ~n74120;
  assign n72513 = n74057 ^ n74058;
  assign n74013 = n74058 & n74065;
  assign n74062 = n74072 & n17111;
  assign n74026 = ~n74073;
  assign n74076 = n74078 & n74079;
  assign n74068 = ~n74085;
  assign n74064 = ~n74086;
  assign n74082 = n74087 & n74067;
  assign n74081 = n70514 & n71524;
  assign n74061 = ~n74091;
  assign n74099 = n74100 & n74101;
  assign n74088 = n74106 & n74107;
  assign n74084 = ~n74110;
  assign n73735 = ~n72513;
  assign n74046 = ~n74062;
  assign n74063 = ~n74076;
  assign n74069 = ~n74081;
  assign n74049 = ~n74082;
  assign n74075 = n74088 ^ n71469;
  assign n74083 = ~n74099;
  assign n74089 = ~n74088;
  assign n74044 = n74063 & n74064;
  assign n74005 = n74068 & n74069;
  assign n70407 = n74074 ^ n74075;
  assign n74066 = n74083 & n74084;
  assign n74080 = n74089 & n74090;
  assign n74029 = n74044 ^ n74045;
  assign n74055 = n70407 & n71469;
  assign n74052 = n74005 & n74024;
  assign n74047 = ~n74044;
  assign n70430 = ~n70407;
  assign n74042 = n74066 ^ n74067;
  assign n74050 = ~n74005;
  assign n74060 = ~n74066;
  assign n74070 = ~n74080;
  assign n74014 = n160 ^ n74029;
  assign n74008 = n74041 ^ n74042;
  assign n74038 = n74046 & n74047;
  assign n74043 = n70430 & n72710;
  assign n74040 = n74050 & n74051;
  assign n74031 = ~n74052;
  assign n74032 = ~n74055;
  assign n74059 = n74060 & n74061;
  assign n74056 = n74070 & n74071;
  assign n72462 = n74013 ^ n74014;
  assign n74012 = ~n74014;
  assign n74028 = n74008 & n175;
  assign n74027 = ~n74008;
  assign n74025 = ~n74038;
  assign n74016 = ~n74040;
  assign n74033 = ~n74043;
  assign n74037 = n74056 ^ n71407;
  assign n74048 = ~n74059;
  assign n74053 = ~n74056;
  assign n73695 = ~n72462;
  assign n73963 = n74012 & n74013;
  assign n74007 = n74025 & n74026;
  assign n74021 = n74027 & n17044;
  assign n73996 = ~n74028;
  assign n73966 = n74032 & n74033;
  assign n70313 = n74036 ^ n74037;
  assign n74023 = n74048 & n74049;
  assign n74039 = n74053 & n74054;
  assign n73991 = n74007 ^ n74008;
  assign n74009 = ~n74007;
  assign n74010 = ~n74021;
  assign n74020 = n70313 & n71434;
  assign n73983 = ~n73966;
  assign n74006 = n74023 ^ n74024;
  assign n70340 = ~n70313;
  assign n74030 = ~n74023;
  assign n74034 = ~n74039;
  assign n73972 = n175 ^ n73991;
  assign n73961 = n74005 ^ n74006;
  assign n74003 = n74009 & n74010;
  assign n74004 = n70340 & n72665;
  assign n73997 = ~n74020;
  assign n74022 = n74030 & n74031;
  assign n74019 = n74034 & n74035;
  assign n72425 = n73963 ^ n73972;
  assign n73962 = ~n73972;
  assign n73992 = n73961 & n17004;
  assign n73995 = ~n74003;
  assign n73993 = ~n73961;
  assign n73998 = ~n74004;
  assign n74000 = n74019 ^ n71368;
  assign n74015 = ~n74022;
  assign n74017 = ~n74019;
  assign n73668 = ~n72425;
  assign n73922 = n73962 & n73963;
  assign n73965 = ~n73992;
  assign n73986 = n73993 & n174;
  assign n73960 = n73995 & n73996;
  assign n73911 = n73997 & n73998;
  assign n70216 = n73999 ^ n74000;
  assign n73987 = n74015 & n74016;
  assign n74011 = n74017 & n74018;
  assign n73925 = ~n73922;
  assign n73946 = n73960 ^ n73961;
  assign n73981 = n73911 & n73985;
  assign n73964 = ~n73960;
  assign n73950 = ~n73986;
  assign n73975 = n70216 & n72634;
  assign n73977 = n70216 & n72723;
  assign n73967 = n73987 ^ n73988;
  assign n73974 = ~n73911;
  assign n70252 = ~n70216;
  assign n73994 = n73987 & n73988;
  assign n73989 = ~n73987;
  assign n74001 = ~n74011;
  assign n73923 = n174 ^ n73946;
  assign n73959 = n73964 & n73965;
  assign n73928 = n73966 ^ n73967;
  assign n73968 = n73974 & n73936;
  assign n73956 = ~n73975;
  assign n73973 = n70252 & n73976;
  assign n72733 = ~n73977;
  assign n73970 = n70252 & n71372;
  assign n73944 = ~n73981;
  assign n73984 = n73989 & n73990;
  assign n73982 = ~n73994;
  assign n73978 = n74001 & n74002;
  assign n72401 = n73922 ^ n73923;
  assign n73924 = ~n73923;
  assign n73947 = n73928 & n16960;
  assign n73949 = ~n73959;
  assign n73948 = ~n73928;
  assign n73918 = ~n73968;
  assign n73955 = ~n73970;
  assign n72719 = ~n73973;
  assign n73952 = n73978 ^ n71316;
  assign n73969 = n73982 & n73983;
  assign n73958 = ~n73984;
  assign n73979 = ~n73978;
  assign n73614 = ~n72401;
  assign n73882 = n73924 & n73925;
  assign n73932 = ~n73947;
  assign n73945 = n73948 & n173;
  assign n73927 = n73949 & n73950;
  assign n70144 = n73951 ^ n73952;
  assign n73876 = n73955 & n73956;
  assign n73957 = ~n73969;
  assign n73971 = n73979 & n73980;
  assign n73908 = n73927 ^ n73928;
  assign n73933 = ~n73927;
  assign n73942 = n73876 & n73898;
  assign n73910 = ~n73945;
  assign n73939 = n70144 & n71343;
  assign n73937 = ~n73876;
  assign n70166 = ~n70144;
  assign n73935 = n73957 & n73958;
  assign n73953 = ~n73971;
  assign n73883 = n173 ^ n73908;
  assign n73921 = n73932 & n73933;
  assign n73931 = n70166 & n72609;
  assign n73912 = n73935 ^ n73936;
  assign n73929 = n73937 & n73938;
  assign n73919 = ~n73939;
  assign n73901 = ~n73942;
  assign n73943 = ~n73935;
  assign n73934 = n73953 & n73954;
  assign n72335 = n73882 ^ n73883;
  assign n73889 = ~n73883;
  assign n73892 = n73911 ^ n73912;
  assign n73909 = ~n73921;
  assign n73873 = ~n73929;
  assign n73920 = ~n73931;
  assign n73916 = n73934 ^ n71269;
  assign n73926 = n73943 & n73944;
  assign n73940 = ~n73934;
  assign n73591 = ~n72335;
  assign n73846 = n73889 & n73882;
  assign n73903 = n73892 & n172;
  assign n73896 = ~n73892;
  assign n73891 = n73909 & n73910;
  assign n70058 = n73915 ^ n73916;
  assign n73829 = n73919 & n73920;
  assign n73917 = ~n73926;
  assign n73930 = n73940 & n73941;
  assign n73845 = ~n73846;
  assign n73869 = n73891 ^ n73892;
  assign n73888 = n73896 & n16911;
  assign n73863 = ~n73903;
  assign n73902 = n70058 & n72642;
  assign n73899 = n70058 & n71271;
  assign n73906 = n73829 & n73855;
  assign n73871 = ~n73891;
  assign n70093 = ~n70058;
  assign n73894 = ~n73829;
  assign n73897 = n73917 & n73918;
  assign n73913 = ~n73930;
  assign n73847 = n172 ^ n73869;
  assign n73870 = ~n73888;
  assign n73884 = n70093 & n73893;
  assign n73887 = n73894 & n73895;
  assign n73877 = n73897 ^ n73898;
  assign n73875 = ~n73899;
  assign n73890 = n70093 & n72544;
  assign n72644 = ~n73902;
  assign n73865 = ~n73906;
  assign n73900 = ~n73897;
  assign n73907 = n73913 & n73914;
  assign n72286 = n73846 ^ n73847;
  assign n73844 = ~n73847;
  assign n73868 = n73870 & n73871;
  assign n73813 = n73876 ^ n73877;
  assign n72660 = ~n73884;
  assign n73832 = ~n73887;
  assign n73874 = ~n73890;
  assign n73886 = n73900 & n73901;
  assign n73879 = n73907 ^ n71200;
  assign n73904 = ~n73907;
  assign n73547 = ~n72286;
  assign n73796 = n73844 & n73845;
  assign n73853 = n73813 & n16887;
  assign n73860 = ~n73813;
  assign n73862 = ~n73868;
  assign n73794 = n73874 & n73875;
  assign n69994 = n73878 ^ n73879;
  assign n73872 = ~n73886;
  assign n73885 = n73904 & n73905;
  assign n73837 = ~n73853;
  assign n73852 = n73860 & n171;
  assign n73839 = n73862 & n73863;
  assign n73858 = n69994 & n72496;
  assign n73859 = n69994 & n72603;
  assign n70020 = ~n69994;
  assign n73800 = ~n73794;
  assign n73854 = n73872 & n73873;
  assign n73880 = ~n73885;
  assign n73812 = n171 ^ n73839;
  assign n73819 = ~n73852;
  assign n73836 = ~n73839;
  assign n73850 = n70020 & n71200;
  assign n73830 = n73854 ^ n73855;
  assign n73834 = ~n73858;
  assign n72625 = ~n73859;
  assign n73849 = n70020 & n73861;
  assign n73864 = ~n73854;
  assign n73867 = n73880 & n73881;
  assign n73797 = n73812 ^ n73813;
  assign n73792 = n73829 ^ n73830;
  assign n73828 = n73836 & n73837;
  assign n72602 = ~n73849;
  assign n73835 = ~n73850;
  assign n73848 = n73864 & n73865;
  assign n69904 = n73866 ^ n73867;
  assign n73856 = ~n73867;
  assign n72233 = n73796 ^ n73797;
  assign n73749 = n73797 & n73796;
  assign n73820 = n73792 & n16859;
  assign n73824 = ~n73792;
  assign n73818 = ~n73828;
  assign n73739 = n73834 & n73835;
  assign n73838 = n69904 & n73843;
  assign n73842 = n69904 & n72459;
  assign n73831 = ~n73848;
  assign n69950 = ~n69904;
  assign n73851 = n73856 & n73857;
  assign n73507 = ~n72233;
  assign n73791 = n73818 & n73819;
  assign n73787 = ~n73820;
  assign n73803 = n73824 & n170;
  assign n73808 = n73739 & n73825;
  assign n73811 = ~n73739;
  assign n73814 = n73831 & n73832;
  assign n73826 = n69950 & n73833;
  assign n72591 = ~n73838;
  assign n73816 = ~n73842;
  assign n73827 = n69950 & n71204;
  assign n73840 = ~n73851;
  assign n73767 = n73791 ^ n73792;
  assign n73788 = ~n73791;
  assign n73771 = ~n73803;
  assign n73759 = ~n73808;
  assign n73805 = n73811 & n73761;
  assign n73795 = n73814 ^ n73815;
  assign n73823 = n73814 & n73815;
  assign n72571 = ~n73826;
  assign n73817 = ~n73827;
  assign n73809 = ~n73814;
  assign n73806 = n73840 & n73841;
  assign n73750 = n170 ^ n73767;
  assign n73782 = n73787 & n73788;
  assign n73757 = n73794 ^ n73795;
  assign n73742 = ~n73805;
  assign n73790 = n73806 ^ n73807;
  assign n73804 = n73809 & n73810;
  assign n73725 = n73816 & n73817;
  assign n73799 = ~n73823;
  assign n73802 = n72591 & n72571;
  assign n73821 = ~n73806;
  assign n72206 = n73749 ^ n73750;
  assign n73712 = n73750 & n73749;
  assign n73774 = n73757 & n16793;
  assign n73776 = ~n73757;
  assign n73770 = ~n73782;
  assign n69888 = n73790 ^ n71100;
  assign n73784 = n73725 & n73798;
  assign n73789 = n73799 & n73800;
  assign n73783 = ~n73725;
  assign n73793 = ~n73790;
  assign n72589 = ~n73802;
  assign n73778 = ~n73804;
  assign n73801 = n73821 & n73822;
  assign n73472 = ~n72206;
  assign n73715 = ~n73712;
  assign n73756 = n73770 & n73771;
  assign n73748 = ~n73774;
  assign n73764 = n73776 & n169;
  assign n73772 = n69888 & n72387;
  assign n73773 = n69888 & n73779;
  assign n69893 = ~n69888;
  assign n73781 = n73783 & n73701;
  assign n73722 = ~n73784;
  assign n73777 = ~n73789;
  assign n73780 = n73793 & n71098;
  assign n73785 = ~n73801;
  assign n73738 = n73756 ^ n73757;
  assign n73747 = ~n73756;
  assign n73733 = ~n73764;
  assign n73765 = n69893 & n72526;
  assign n73762 = ~n73772;
  assign n72552 = ~n73773;
  assign n73760 = n73777 & n73778;
  assign n73763 = ~n73780;
  assign n73705 = ~n73781;
  assign n73775 = n73785 & n73786;
  assign n73713 = n169 ^ n73738;
  assign n73746 = n73747 & n73748;
  assign n73740 = n73760 ^ n73761;
  assign n73687 = n73762 & n73763;
  assign n72531 = ~n73765;
  assign n73758 = ~n73760;
  assign n73753 = n73775 ^ n70999;
  assign n73768 = ~n73775;
  assign n72109 = n73712 ^ n73713;
  assign n73714 = ~n73713;
  assign n73709 = n73739 ^ n73740;
  assign n73732 = ~n73746;
  assign n73745 = n73687 & n73663;
  assign n73743 = ~n73687;
  assign n69831 = n73752 ^ n73753;
  assign n73751 = n73758 & n73759;
  assign n73766 = n73768 & n73769;
  assign n73429 = ~n72109;
  assign n73676 = n73714 & n73715;
  assign n73720 = n73709 & n168;
  assign n73723 = ~n73709;
  assign n73708 = n73732 & n73733;
  assign n73729 = n69831 & n72364;
  assign n73734 = n69831 & n72513;
  assign n73731 = n73743 & n73744;
  assign n73682 = ~n73745;
  assign n69839 = ~n69831;
  assign n73741 = ~n73751;
  assign n73754 = ~n73766;
  assign n73698 = n73708 ^ n73709;
  assign n73684 = ~n73720;
  assign n73717 = n73723 & n16739;
  assign n73703 = ~n73708;
  assign n73711 = ~n73729;
  assign n73670 = ~n73731;
  assign n72517 = ~n73734;
  assign n73727 = n69839 & n70999;
  assign n73726 = n69839 & n73735;
  assign n73724 = n73741 & n73742;
  assign n73730 = n73754 & n73755;
  assign n73677 = n168 ^ n73698;
  assign n73702 = ~n73717;
  assign n73700 = n73724 ^ n73725;
  assign n72504 = ~n73726;
  assign n73710 = ~n73727;
  assign n73707 = n73730 ^ n70908;
  assign n73721 = ~n73724;
  assign n73736 = ~n73730;
  assign n72037 = n73676 ^ n73677;
  assign n73623 = n73677 & n73676;
  assign n73667 = n73700 ^ n73701;
  assign n73694 = n73702 & n73703;
  assign n69781 = n73706 ^ n73707;
  assign n73642 = n73710 & n73711;
  assign n73716 = n73721 & n73722;
  assign n73728 = n73736 & n73737;
  assign n73374 = ~n72037;
  assign n73688 = n73667 & n183;
  assign n73683 = ~n73694;
  assign n73685 = ~n73667;
  assign n73696 = n69781 & n72462;
  assign n73699 = n69781 & n72403;
  assign n73630 = ~n73642;
  assign n69793 = ~n69781;
  assign n73704 = ~n73716;
  assign n73718 = ~n73728;
  assign n73666 = n73683 & n73684;
  assign n73678 = n73685 & n16715;
  assign n73647 = ~n73688;
  assign n73690 = n69793 & n73695;
  assign n73689 = n69793 & n71005;
  assign n72483 = ~n73696;
  assign n73671 = ~n73699;
  assign n73686 = n73704 & n73705;
  assign n73697 = n73718 & n73719;
  assign n73644 = n73666 ^ n73667;
  assign n73664 = ~n73666;
  assign n73665 = ~n73678;
  assign n73662 = n73686 ^ n73687;
  assign n73672 = ~n73689;
  assign n72461 = ~n73690;
  assign n73680 = n73697 ^ n70833;
  assign n73681 = ~n73686;
  assign n73692 = ~n73697;
  assign n73624 = n183 ^ n73644;
  assign n73607 = n73662 ^ n73663;
  assign n73658 = n73664 & n73665;
  assign n73570 = n73671 & n73672;
  assign n69745 = n73679 ^ n73680;
  assign n73673 = n73681 & n73682;
  assign n73691 = n73692 & n73693;
  assign n71953 = n73623 ^ n73624;
  assign n73583 = n73624 & n73623;
  assign n73641 = n73607 & n16633;
  assign n73646 = ~n73658;
  assign n73640 = ~n73607;
  assign n73656 = n73570 & n73593;
  assign n73655 = n69745 & n70941;
  assign n73657 = n69745 & n73668;
  assign n73659 = ~n73570;
  assign n69750 = ~n69745;
  assign n73669 = ~n73673;
  assign n73674 = ~n73691;
  assign n73329 = ~n71953;
  assign n73635 = n73640 & n182;
  assign n73622 = ~n73641;
  assign n73628 = n73646 & n73647;
  assign n73638 = ~n73655;
  assign n73595 = ~n73656;
  assign n73651 = n69750 & n72425;
  assign n72424 = ~n73657;
  assign n73649 = n73659 & n73660;
  assign n73652 = n69750 & n72359;
  assign n73643 = n73669 & n73670;
  assign n73661 = n73674 & n73675;
  assign n73606 = n182 ^ n73628;
  assign n73604 = ~n73635;
  assign n73621 = ~n73628;
  assign n73625 = n73642 ^ n73643;
  assign n73639 = n73643 & n73648;
  assign n73566 = ~n73649;
  assign n72444 = ~n73651;
  assign n73637 = ~n73652;
  assign n73645 = ~n73643;
  assign n73634 = n73661 ^ n70760;
  assign n73653 = ~n73661;
  assign n73584 = n73606 ^ n73607;
  assign n73615 = n73621 & n73622;
  assign n73586 = n73625 ^ n73626;
  assign n69690 = n73633 ^ n73634;
  assign n73527 = n73637 & n73638;
  assign n73629 = ~n73639;
  assign n73636 = n73645 & n73626;
  assign n73650 = n73653 & n73654;
  assign n71864 = n73583 ^ n73584;
  assign n73587 = ~n73584;
  assign n73608 = n73586 & n181;
  assign n73605 = ~n73586;
  assign n73603 = ~n73615;
  assign n73616 = n69690 & n72401;
  assign n73617 = n69690 & n72320;
  assign n73540 = ~n73527;
  assign n69707 = ~n69690;
  assign n73627 = n73629 & n73630;
  assign n73611 = ~n73636;
  assign n73631 = ~n73650;
  assign n73263 = ~n71864;
  assign n73544 = n73587 & n73583;
  assign n73585 = n73603 & n73604;
  assign n73602 = n73605 & n16558;
  assign n73563 = ~n73608;
  assign n73609 = n69707 & n73614;
  assign n72406 = ~n73616;
  assign n73601 = ~n73617;
  assign n73613 = n69707 & n70859;
  assign n73610 = ~n73627;
  assign n73620 = n73631 & n73632;
  assign n73564 = n73585 ^ n73586;
  assign n73588 = ~n73585;
  assign n73589 = ~n73602;
  assign n72380 = ~n73609;
  assign n73592 = n73610 & n73611;
  assign n73600 = ~n73613;
  assign n73599 = n73620 ^ n70682;
  assign n73618 = ~n73620;
  assign n73545 = n181 ^ n73564;
  assign n73582 = n73588 & n73589;
  assign n73571 = n73592 ^ n73593;
  assign n69656 = n73598 ^ n73599;
  assign n73504 = n73600 & n73601;
  assign n73594 = ~n73592;
  assign n73612 = n73618 & n73619;
  assign n71787 = n73544 ^ n73545;
  assign n73178 = n73545 & n73544;
  assign n73542 = n73570 ^ n73571;
  assign n73562 = ~n73582;
  assign n73578 = n73504 & n73483;
  assign n73579 = n69656 & n73591;
  assign n73575 = n69656 & n72259;
  assign n73580 = ~n73504;
  assign n69653 = ~n69656;
  assign n73590 = n73594 & n73595;
  assign n73596 = ~n73612;
  assign n73223 = ~n71787;
  assign n73511 = ~n73178;
  assign n73553 = n73542 & n16510;
  assign n73541 = n73562 & n73563;
  assign n73548 = ~n73542;
  assign n73559 = ~n73575;
  assign n73502 = ~n73578;
  assign n73569 = n69653 & n70682;
  assign n72351 = ~n73579;
  assign n73572 = n73580 & n73581;
  assign n73567 = n69653 & n72335;
  assign n73565 = ~n73590;
  assign n73573 = n73596 & n73597;
  assign n73524 = n73541 ^ n73542;
  assign n73546 = n73548 & n180;
  assign n73535 = ~n73553;
  assign n73536 = ~n73541;
  assign n73549 = n73565 & n73566;
  assign n72329 = ~n73567;
  assign n73560 = ~n73569;
  assign n73475 = ~n73572;
  assign n73561 = n73573 ^ n73574;
  assign n73576 = ~n73573;
  assign n73147 = n180 ^ n73524;
  assign n73525 = n73535 & n73536;
  assign n73520 = ~n73546;
  assign n73528 = n73549 ^ n73550;
  assign n73435 = n73559 & n73560;
  assign n69600 = n70594 ^ n73561;
  assign n73555 = n73549 & n73550;
  assign n73551 = ~n73549;
  assign n73558 = ~n73561;
  assign n73568 = n73576 & n73577;
  assign n73457 = n73147 & n73511;
  assign n73519 = ~n73525;
  assign n73494 = n73527 ^ n73528;
  assign n73531 = n69600 & n72193;
  assign n73534 = n69600 & n73547;
  assign n69614 = ~n69600;
  assign n73543 = n73551 & n73552;
  assign n73449 = ~n73435;
  assign n73539 = ~n73555;
  assign n73554 = n73558 & n70696;
  assign n73556 = ~n73568;
  assign n73509 = n73494 & n16437;
  assign n73493 = n73519 & n73520;
  assign n73513 = ~n73494;
  assign n73522 = ~n73531;
  assign n72310 = ~n73534;
  assign n73529 = n69614 & n72286;
  assign n73530 = n73539 & n73540;
  assign n73518 = ~n73543;
  assign n73523 = ~n73554;
  assign n73537 = n73556 & n73557;
  assign n73484 = n73493 ^ n73494;
  assign n73492 = ~n73509;
  assign n73491 = ~n73493;
  assign n73508 = n73513 & n179;
  assign n73387 = n73522 & n73523;
  assign n72289 = ~n73529;
  assign n73517 = ~n73530;
  assign n73516 = n73537 ^ n73538;
  assign n73532 = ~n73537;
  assign n73458 = n179 ^ n73484;
  assign n73487 = n73491 & n73492;
  assign n73481 = ~n73508;
  assign n73505 = n73387 & n73510;
  assign n73506 = ~n73387;
  assign n69544 = n70479 ^ n73516;
  assign n73503 = n73517 & n73518;
  assign n73521 = ~n73516;
  assign n73526 = n73532 & n73533;
  assign n73437 = n73457 ^ n73458;
  assign n73417 = n73458 & n73457;
  assign n73480 = ~n73487;
  assign n73482 = n73503 ^ n73504;
  assign n73405 = ~n73505;
  assign n73497 = n73506 & n73408;
  assign n73496 = n69544 & n72131;
  assign n73495 = n69544 & n73507;
  assign n69581 = ~n69544;
  assign n73501 = ~n73503;
  assign n73512 = n73521 & n70656;
  assign n73514 = ~n73526;
  assign n69342 = n73437 ^ n71288;
  assign n73343 = n73437 & n71284;
  assign n73445 = ~n73437;
  assign n73459 = n73480 & n73481;
  assign n73460 = n73482 ^ n73483;
  assign n73490 = n69581 & n72233;
  assign n72252 = ~n73495;
  assign n73485 = ~n73496;
  assign n73386 = ~n73497;
  assign n73489 = n73501 & n73502;
  assign n73486 = ~n73512;
  assign n73500 = n73514 & n73515;
  assign n73416 = n69342 & n72331;
  assign n69344 = ~n69342;
  assign n73434 = n73445 & n71284;
  assign n73446 = n73459 ^ n73460;
  assign n73471 = n73460 & n16378;
  assign n73451 = ~n73459;
  assign n73470 = ~n73460;
  assign n73355 = n73485 & n73486;
  assign n73474 = ~n73489;
  assign n72228 = ~n73490;
  assign n73479 = n73500 ^ n70441;
  assign n73498 = ~n73500;
  assign n73402 = ~n73416;
  assign n73403 = ~n73434;
  assign n73418 = n178 ^ n73446;
  assign n73452 = n73470 & n178;
  assign n73450 = ~n73471;
  assign n73337 = ~n73355;
  assign n73468 = n73474 & n73475;
  assign n69532 = n73478 ^ n73479;
  assign n73488 = n73498 & n73499;
  assign n73379 = n73402 & n73403;
  assign n73406 = n73417 ^ n73418;
  assign n73358 = n73418 & n73417;
  assign n73438 = n73450 & n73451;
  assign n73431 = ~n73452;
  assign n73436 = n73468 ^ n73466;
  assign n73467 = n69532 & n71926;
  assign n73469 = n69532 & n73472;
  assign n73461 = n73468 & n73473;
  assign n73465 = ~n73468;
  assign n69517 = ~n69532;
  assign n73476 = ~n73488;
  assign n73352 = n73379 ^ n73380;
  assign n73381 = ~n73379;
  assign n73399 = n73406 & n71172;
  assign n73391 = ~n73406;
  assign n73410 = n73435 ^ n73436;
  assign n73430 = ~n73438;
  assign n73448 = ~n73461;
  assign n73453 = n69517 & n72206;
  assign n73455 = n73465 & n73466;
  assign n73442 = ~n73467;
  assign n72208 = ~n73469;
  assign n73454 = n69517 & n70441;
  assign n73464 = n73476 & n73477;
  assign n71196 = n199 ^ n73352;
  assign n73099 = n73352 & n199;
  assign n73203 = n73381 & n73382;
  assign n73390 = n73391 & n71175;
  assign n73339 = ~n73399;
  assign n73409 = n73430 & n73431;
  assign n73423 = n73410 & n177;
  assign n73422 = ~n73410;
  assign n73447 = n73448 & n73449;
  assign n72174 = ~n73453;
  assign n73441 = ~n73454;
  assign n73433 = ~n73455;
  assign n73440 = n73464 ^ n70296;
  assign n73462 = ~n73464;
  assign n71237 = ~n71196;
  assign n73373 = ~n73390;
  assign n73384 = n73409 ^ n73410;
  assign n73411 = n73422 & n16277;
  assign n73371 = ~n73423;
  assign n73401 = ~n73409;
  assign n69467 = n73439 ^ n73440;
  assign n73286 = n73441 & n73442;
  assign n73432 = ~n73447;
  assign n73456 = n73462 & n73463;
  assign n73362 = n73373 & n73343;
  assign n73342 = n73373 & n73339;
  assign n73359 = n177 ^ n73384;
  assign n73400 = ~n73411;
  assign n73427 = n69467 & n73429;
  assign n73424 = n69467 & n70296;
  assign n73428 = n73286 & n73257;
  assign n73407 = n73432 & n73433;
  assign n73425 = ~n73286;
  assign n69510 = ~n69467;
  assign n73443 = ~n73456;
  assign n69260 = n73342 ^ n73343;
  assign n73297 = n73358 ^ n73359;
  assign n73338 = ~n73362;
  assign n73360 = ~n73359;
  assign n73389 = n73400 & n73401;
  assign n73388 = n73407 ^ n73408;
  assign n73404 = ~n73407;
  assign n73415 = n69510 & n72109;
  assign n73414 = n69510 & n71986;
  assign n73396 = ~n73424;
  assign n73413 = n73425 & n73426;
  assign n72096 = ~n73427;
  assign n73284 = ~n73428;
  assign n73421 = n73443 & n73444;
  assign n73320 = n69260 & n71172;
  assign n69266 = ~n69260;
  assign n73324 = n73338 & n73339;
  assign n73302 = ~n73297;
  assign n73287 = n73360 & n73358;
  assign n73347 = n73387 ^ n73388;
  assign n73370 = ~n73389;
  assign n73392 = n73404 & n73405;
  assign n73252 = ~n73413;
  assign n73395 = ~n73414;
  assign n72144 = ~n73415;
  assign n73394 = n73421 ^ n70249;
  assign n73419 = ~n73421;
  assign n73290 = ~n73320;
  assign n73315 = n69266 & n72191;
  assign n73298 = n73324 ^ n71089;
  assign n73328 = n73324 & n71089;
  assign n73323 = ~n73324;
  assign n73307 = ~n73287;
  assign n73354 = n73347 & n176;
  assign n73346 = n73370 & n73371;
  assign n73357 = ~n73347;
  assign n73385 = ~n73392;
  assign n69427 = n73393 ^ n73394;
  assign n73196 = n73395 & n73396;
  assign n73412 = n73419 & n73420;
  assign n69191 = n73297 ^ n73298;
  assign n73289 = ~n73315;
  assign n73308 = n73323 & n71118;
  assign n73301 = ~n73328;
  assign n73319 = n73346 ^ n73347;
  assign n73304 = ~n73354;
  assign n73341 = n73357 & n16229;
  assign n73333 = ~n73346;
  assign n73375 = n73196 & n73383;
  assign n73376 = n69427 & n72037;
  assign n73378 = n69427 & n71912;
  assign n73356 = n73385 & n73386;
  assign n73372 = ~n73196;
  assign n69472 = ~n69427;
  assign n73397 = ~n73412;
  assign n73271 = n69191 & n72117;
  assign n69218 = ~n69191;
  assign n73279 = n73289 & n73290;
  assign n73291 = n73301 & n73302;
  assign n73275 = ~n73308;
  assign n73288 = n176 ^ n73319;
  assign n73332 = ~n73341;
  assign n73330 = n73355 ^ n73356;
  assign n73353 = n73356 & n73366;
  assign n73363 = n73372 & n73228;
  assign n73361 = ~n73356;
  assign n73367 = n69472 & n73374;
  assign n73230 = ~n73375;
  assign n73365 = n69472 & n70257;
  assign n72071 = ~n73376;
  assign n73351 = ~n73378;
  assign n73377 = n73397 & n73398;
  assign n73259 = n69218 & n71118;
  assign n73239 = ~n73271;
  assign n73270 = n73279 & n73280;
  assign n73272 = ~n73279;
  assign n73216 = n73287 ^ n73288;
  assign n73274 = ~n73291;
  assign n73219 = n73288 & n73307;
  assign n73277 = n73330 ^ n73331;
  assign n73316 = n73332 & n73333;
  assign n73336 = ~n73353;
  assign n73340 = n73361 & n73331;
  assign n73201 = ~n73363;
  assign n73350 = ~n73365;
  assign n72020 = ~n73367;
  assign n73349 = n73377 ^ n70158;
  assign n73368 = ~n73377;
  assign n73240 = ~n73259;
  assign n73242 = ~n73270;
  assign n73253 = n73272 & n73273;
  assign n73250 = n73274 & n73275;
  assign n73266 = n73216 & n71030;
  assign n73269 = ~n73216;
  assign n73305 = n73277 & n191;
  assign n73303 = ~n73316;
  assign n73306 = ~n73277;
  assign n73334 = n73336 & n73337;
  assign n73313 = ~n73340;
  assign n69381 = n73348 ^ n73349;
  assign n73139 = n73350 & n73351;
  assign n73364 = n73368 & n73369;
  assign n73157 = n73239 & n73240;
  assign n73217 = n73250 ^ n71030;
  assign n73241 = n73242 & n73203;
  assign n73222 = ~n73253;
  assign n73244 = ~n73250;
  assign n73215 = ~n73266;
  assign n73260 = n73269 & n71049;
  assign n73276 = n73303 & n73304;
  assign n73248 = ~n73305;
  assign n73296 = n73306 & n16084;
  assign n73325 = n69381 & n73329;
  assign n73326 = n69381 & n70298;
  assign n73312 = ~n73334;
  assign n73321 = n73139 & n73335;
  assign n73322 = ~n73139;
  assign n69430 = ~n69381;
  assign n73344 = ~n73364;
  assign n69172 = n73216 ^ n73217;
  assign n73162 = ~n73157;
  assign n73221 = ~n73241;
  assign n73231 = n73222 & n73242;
  assign n73243 = ~n73260;
  assign n73249 = n73276 ^ n73277;
  assign n73281 = ~n73276;
  assign n73282 = ~n73296;
  assign n73285 = n73312 & n73313;
  assign n73309 = n69430 & n71953;
  assign n73168 = ~n73321;
  assign n73314 = n73322 & n73171;
  assign n71956 = ~n73325;
  assign n73311 = n69430 & n71696;
  assign n73294 = ~n73326;
  assign n73327 = n73344 & n73345;
  assign n73189 = n69172 & n72025;
  assign n69170 = ~n69172;
  assign n73186 = n73221 & n73222;
  assign n73204 = ~n73231;
  assign n73234 = n73243 & n73244;
  assign n73220 = n191 ^ n73249;
  assign n73267 = n73281 & n73282;
  assign n73256 = n73285 ^ n73286;
  assign n73283 = ~n73285;
  assign n71996 = ~n73309;
  assign n73295 = ~n73311;
  assign n73135 = ~n73314;
  assign n73300 = n73327 ^ n70084;
  assign n73317 = ~n73327;
  assign n73158 = n73186 ^ n73187;
  assign n73180 = n69170 & n71030;
  assign n73154 = ~n73189;
  assign n73191 = n73186 & n73198;
  assign n73179 = n73203 ^ n73204;
  assign n73193 = ~n73186;
  assign n73141 = n73219 ^ n73220;
  assign n73214 = ~n73234;
  assign n73151 = n73220 & n73219;
  assign n73225 = n73256 ^ n73257;
  assign n73247 = ~n73267;
  assign n73278 = n73283 & n73284;
  assign n73078 = n73294 & n73295;
  assign n69336 = n73299 ^ n73300;
  assign n73310 = n73317 & n73318;
  assign n73070 = n73157 ^ n73158;
  assign n73164 = n73179 & n8617;
  assign n73153 = ~n73180;
  assign n73161 = ~n73191;
  assign n73163 = ~n73179;
  assign n73177 = n73193 & n73187;
  assign n73192 = n73141 & n70953;
  assign n73188 = ~n73141;
  assign n73174 = n73214 & n73215;
  assign n73232 = n73225 & n16051;
  assign n73224 = n73247 & n73248;
  assign n73233 = ~n73225;
  assign n73268 = n69336 & n70084;
  assign n73251 = ~n73278;
  assign n73264 = n69336 & n71864;
  assign n69394 = ~n69336;
  assign n73092 = ~n73078;
  assign n73292 = ~n73310;
  assign n73071 = n73153 & n73154;
  assign n73152 = n73161 & n73162;
  assign n73149 = n73163 & n198;
  assign n73138 = ~n73164;
  assign n73142 = n73174 ^ n70934;
  assign n73130 = ~n73177;
  assign n73184 = n73188 & n70934;
  assign n73165 = ~n73192;
  assign n73166 = ~n73174;
  assign n73190 = n73224 ^ n73225;
  assign n73206 = ~n73232;
  assign n73226 = n73233 & n190;
  assign n73207 = ~n73224;
  assign n73227 = n73251 & n73252;
  assign n73254 = n69394 & n73263;
  assign n71863 = ~n73264;
  assign n73258 = n69394 & n71606;
  assign n73238 = ~n73268;
  assign n73265 = n73292 & n73293;
  assign n69115 = n73141 ^ n73142;
  assign n73094 = ~n73071;
  assign n73131 = n73138 & n73099;
  assign n73121 = ~n73149;
  assign n73129 = ~n73152;
  assign n73155 = n73165 & n73166;
  assign n73137 = ~n73184;
  assign n73156 = n190 ^ n73190;
  assign n73194 = n73206 & n73207;
  assign n73176 = ~n73226;
  assign n73197 = n73227 ^ n73228;
  assign n73229 = ~n73227;
  assign n71903 = ~n73254;
  assign n73237 = ~n73258;
  assign n73236 = n73265 ^ n70016;
  assign n73261 = ~n73265;
  assign n73124 = n69115 & n70934;
  assign n73108 = n73129 & n73130;
  assign n73120 = ~n73131;
  assign n69131 = ~n69115;
  assign n73128 = n73138 & n73121;
  assign n73136 = ~n73155;
  assign n73080 = n73151 ^ n73156;
  assign n73150 = ~n73156;
  assign n73175 = ~n73194;
  assign n73146 = n73196 ^ n73197;
  assign n73218 = n73229 & n73230;
  assign n69297 = n73235 ^ n73236;
  assign n73003 = n73237 & n73238;
  assign n73255 = n73261 & n73262;
  assign n73072 = n73108 ^ n73109;
  assign n73083 = n73120 & n73121;
  assign n73088 = ~n73124;
  assign n73114 = n69131 & n71934;
  assign n73115 = n73108 & n73109;
  assign n73103 = ~n73108;
  assign n73100 = ~n73128;
  assign n73127 = n73080 & n70851;
  assign n73113 = n73136 & n73137;
  assign n73125 = ~n73080;
  assign n73089 = n73150 & n73151;
  assign n73145 = n73175 & n73176;
  assign n73172 = n73146 & n189;
  assign n73173 = ~n73146;
  assign n73208 = n69297 & n70016;
  assign n73200 = ~n73218;
  assign n73211 = n69297 & n73223;
  assign n73205 = n73003 & n73033;
  assign n73209 = ~n73003;
  assign n69306 = ~n69297;
  assign n73245 = ~n73255;
  assign n73010 = n73071 ^ n73072;
  assign n73056 = n73083 ^ n73070;
  assign n73065 = n73099 ^ n73100;
  assign n73085 = n73083 & n8554;
  assign n73101 = n73103 & n73104;
  assign n73084 = ~n73083;
  assign n73081 = n73113 ^ n70845;
  assign n73087 = ~n73114;
  assign n73093 = ~n73115;
  assign n73119 = n73125 & n70845;
  assign n73067 = ~n73127;
  assign n73097 = ~n73113;
  assign n73118 = n73145 ^ n73146;
  assign n73132 = ~n73145;
  assign n73107 = ~n73172;
  assign n73160 = n73173 & n15951;
  assign n73170 = n73200 & n73201;
  assign n73041 = ~n73205;
  assign n73199 = n69306 & n71787;
  assign n73183 = ~n73208;
  assign n73202 = n69306 & n71553;
  assign n73195 = n73209 & n73210;
  assign n71847 = ~n73211;
  assign n73212 = n73245 & n73246;
  assign n73030 = n197 ^ n73056;
  assign n72988 = ~n73010;
  assign n72486 = n73065 ^ n71237;
  assign n73029 = n73065 & n71237;
  assign n69077 = n73080 ^ n73081;
  assign n73076 = n73084 & n197;
  assign n73069 = ~n73085;
  assign n72996 = n73087 & n73088;
  assign n73082 = n73093 & n73094;
  assign n73058 = ~n73101;
  assign n73090 = n189 ^ n73118;
  assign n73096 = ~n73119;
  assign n73133 = ~n73160;
  assign n73140 = n73170 ^ n73171;
  assign n73167 = ~n73170;
  assign n73002 = ~n73195;
  assign n71807 = ~n73199;
  assign n73182 = ~n73202;
  assign n69315 = n73212 ^ n73213;
  assign n71104 = n73029 ^ n73030;
  assign n73036 = ~n73030;
  assign n71160 = ~n72486;
  assign n73052 = n69077 & n70851;
  assign n73037 = ~n73029;
  assign n69094 = ~n69077;
  assign n73059 = n73069 & n73070;
  assign n73047 = ~n73076;
  assign n73057 = ~n73082;
  assign n73012 = ~n72996;
  assign n73000 = n73089 ^ n73090;
  assign n73086 = n73096 & n73097;
  assign n73024 = n73090 & n73089;
  assign n73126 = n73132 & n73133;
  assign n73055 = n73139 ^ n73140;
  assign n73159 = n73167 & n73168;
  assign n73148 = n73178 ^ n69315;
  assign n72945 = n73182 & n73183;
  assign n73185 = n69315 & n71657;
  assign n73181 = ~n69315;
  assign n72445 = ~n71104;
  assign n72948 = n73036 & n73037;
  assign n73044 = n69094 & n71828;
  assign n73027 = ~n73052;
  assign n73034 = n73057 & n73058;
  assign n73046 = ~n73059;
  assign n73061 = n73000 & n70745;
  assign n73062 = ~n73000;
  assign n73066 = ~n73086;
  assign n73020 = ~n73024;
  assign n73102 = n73055 & n188;
  assign n73106 = ~n73126;
  assign n73105 = ~n73055;
  assign n71771 = n73147 ^ n73148;
  assign n73134 = ~n73159;
  assign n72951 = ~n72945;
  assign n73169 = n73181 & n70079;
  assign n73144 = ~n73185;
  assign n72997 = n73034 ^ n73035;
  assign n73026 = ~n73044;
  assign n73031 = n73034 & n73045;
  assign n73009 = n73046 & n73047;
  assign n73038 = ~n73034;
  assign n73042 = ~n73061;
  assign n73051 = n73062 & n70743;
  assign n73060 = n73066 & n73067;
  assign n73050 = ~n73102;
  assign n73098 = n73105 & n15860;
  assign n73077 = n73106 & n73107;
  assign n73116 = n73134 & n73135;
  assign n73143 = ~n73169;
  assign n72922 = n72996 ^ n72997;
  assign n72986 = n73009 ^ n73010;
  assign n73008 = n73009 & n8495;
  assign n72927 = n73026 & n73027;
  assign n73007 = ~n73009;
  assign n73011 = ~n73031;
  assign n73016 = n73038 & n73035;
  assign n73015 = ~n73051;
  assign n73039 = ~n73060;
  assign n73054 = n188 ^ n73077;
  assign n73073 = ~n73098;
  assign n73074 = ~n73077;
  assign n73079 = n73116 ^ n73117;
  assign n73112 = n73116 & n73117;
  assign n73110 = ~n73116;
  assign n73122 = n73143 & n73144;
  assign n72949 = n196 ^ n72986;
  assign n72991 = n72927 & n73005;
  assign n72998 = n73007 & n196;
  assign n72995 = ~n72927;
  assign n72987 = ~n73008;
  assign n73006 = n73011 & n73012;
  assign n72982 = ~n73016;
  assign n72999 = n73039 ^ n70743;
  assign n73028 = n73042 & n73039;
  assign n73025 = n73054 ^ n73055;
  assign n73068 = n73073 & n73074;
  assign n73018 = n73078 ^ n73079;
  assign n73095 = n73110 & n73111;
  assign n73091 = ~n73112;
  assign n72874 = n73122 ^ n73123;
  assign n71077 = n72948 ^ n72949;
  assign n72884 = n72949 & n72948;
  assign n72979 = n72987 & n72988;
  assign n72957 = ~n72991;
  assign n72985 = n72995 & n72955;
  assign n72971 = ~n72998;
  assign n69039 = n72999 ^ n73000;
  assign n72981 = ~n73006;
  assign n72959 = n73024 ^ n73025;
  assign n73014 = ~n73028;
  assign n73019 = ~n73025;
  assign n73053 = n73018 & n15777;
  assign n73048 = ~n73018;
  assign n73049 = ~n73068;
  assign n73075 = n73091 & n73092;
  assign n73064 = ~n73095;
  assign n72407 = ~n71077;
  assign n72898 = ~n72884;
  assign n72970 = ~n72979;
  assign n72976 = n69039 & n71769;
  assign n72954 = n72981 & n72982;
  assign n72926 = ~n72985;
  assign n69048 = ~n69039;
  assign n72989 = n72959 & n70634;
  assign n72990 = ~n72959;
  assign n72980 = n73014 & n73015;
  assign n72968 = n73019 & n73020;
  assign n73043 = n73048 & n187;
  assign n73017 = n73049 & n73050;
  assign n73023 = ~n73053;
  assign n73063 = ~n73075;
  assign n72928 = n72954 ^ n72955;
  assign n72940 = n72970 & n72971;
  assign n72958 = ~n72954;
  assign n72964 = n69048 & n70743;
  assign n72941 = ~n72976;
  assign n72960 = n72980 ^ n70634;
  assign n72938 = ~n72989;
  assign n72984 = n72990 & n70684;
  assign n72961 = ~n72980;
  assign n72994 = n73017 ^ n73018;
  assign n72993 = ~n73043;
  assign n73022 = ~n73017;
  assign n73032 = n73063 & n73064;
  assign n72863 = n72927 ^ n72928;
  assign n72911 = n72940 ^ n72922;
  assign n72935 = n72940 & n8474;
  assign n72939 = ~n72940;
  assign n72944 = n72957 & n72958;
  assign n68999 = n72959 ^ n72960;
  assign n72942 = ~n72964;
  assign n72962 = ~n72984;
  assign n72969 = n187 ^ n72994;
  assign n73013 = n73022 & n73023;
  assign n73004 = n73032 ^ n73033;
  assign n73040 = ~n73032;
  assign n72885 = n195 ^ n72911;
  assign n72905 = n72863 & n194;
  assign n72904 = ~n72863;
  assign n72929 = n68999 & n71663;
  assign n72921 = ~n72935;
  assign n72932 = n72939 & n195;
  assign n72871 = n72941 & n72942;
  assign n69008 = ~n68999;
  assign n72925 = ~n72944;
  assign n72956 = n72961 & n72962;
  assign n72889 = n72968 ^ n72969;
  assign n72917 = n72969 & n72968;
  assign n72966 = n73003 ^ n73004;
  assign n72992 = ~n73013;
  assign n73021 = n73040 & n73041;
  assign n70958 = n72884 ^ n72885;
  assign n72826 = n72885 & n72898;
  assign n72895 = n72904 & n8425;
  assign n72849 = ~n72905;
  assign n72912 = n72921 & n72922;
  assign n72899 = n72925 & n72926;
  assign n72908 = ~n72929;
  assign n72894 = ~n72932;
  assign n72924 = n69008 & n70634;
  assign n72883 = ~n72871;
  assign n72937 = ~n72956;
  assign n72977 = n72966 & n15671;
  assign n72972 = ~n72966;
  assign n72965 = n72992 & n72993;
  assign n73001 = ~n73021;
  assign n72369 = ~n70958;
  assign n72832 = ~n72826;
  assign n72869 = ~n72895;
  assign n72872 = n72899 ^ n72900;
  assign n72893 = ~n72912;
  assign n72909 = n72899 & n72916;
  assign n72910 = ~n72899;
  assign n72907 = ~n72924;
  assign n72913 = n72937 & n72938;
  assign n72936 = n72965 ^ n72966;
  assign n72967 = n72972 & n186;
  assign n72952 = ~n72977;
  assign n72953 = ~n72965;
  assign n72973 = n73001 & n73002;
  assign n72825 = n72871 ^ n72872;
  assign n72862 = n72893 & n72894;
  assign n72817 = n72907 & n72908;
  assign n72882 = ~n72909;
  assign n72892 = n72910 & n72900;
  assign n72890 = n72913 ^ n70554;
  assign n72915 = n72913 & n70603;
  assign n72919 = ~n72913;
  assign n72918 = n186 ^ n72936;
  assign n72947 = n72952 & n72953;
  assign n72934 = ~n72967;
  assign n72946 = n72973 ^ n72974;
  assign n72978 = n72973 & n72983;
  assign n72975 = ~n72973;
  assign n72853 = n72825 & n193;
  assign n72847 = n72862 ^ n72863;
  assign n72854 = ~n72825;
  assign n72877 = n72882 & n72883;
  assign n72870 = ~n72862;
  assign n72876 = n72817 & n72844;
  assign n68963 = n72889 ^ n72890;
  assign n72861 = ~n72892;
  assign n72879 = ~n72817;
  assign n72891 = ~n72915;
  assign n72822 = n72917 ^ n72918;
  assign n72906 = n72919 & n70554;
  assign n72855 = n72918 & n72917;
  assign n72902 = n72945 ^ n72946;
  assign n72933 = ~n72947;
  assign n72963 = n72975 & n72974;
  assign n72950 = ~n72978;
  assign n72827 = n194 ^ n72847;
  assign n72807 = ~n72853;
  assign n72846 = n72854 & n8392;
  assign n72857 = n68963 & n71610;
  assign n72859 = n72869 & n72870;
  assign n68972 = ~n68963;
  assign n72836 = ~n72876;
  assign n72860 = ~n72877;
  assign n72866 = n72879 & n72880;
  assign n72886 = n72891 & n72889;
  assign n72888 = n72822 & n70514;
  assign n72868 = ~n72906;
  assign n72881 = ~n72822;
  assign n72858 = ~n72855;
  assign n72923 = n72902 & n185;
  assign n72901 = n72933 & n72934;
  assign n72920 = ~n72902;
  assign n72943 = n72950 & n72951;
  assign n72931 = ~n72963;
  assign n70893 = n72826 ^ n72827;
  assign n72831 = ~n72827;
  assign n72828 = ~n72846;
  assign n72841 = ~n72857;
  assign n72848 = ~n72859;
  assign n72843 = n72860 & n72861;
  assign n72852 = n68972 & n70554;
  assign n72816 = ~n72866;
  assign n72875 = n72881 & n70491;
  assign n72867 = ~n72886;
  assign n72821 = ~n72888;
  assign n72878 = n72901 ^ n72902;
  assign n72914 = n72920 & n15638;
  assign n72896 = ~n72901;
  assign n72865 = ~n72923;
  assign n72930 = ~n72943;
  assign n72311 = ~n70893;
  assign n72777 = n72831 & n72832;
  assign n72818 = n72843 ^ n72844;
  assign n72824 = n72848 & n72849;
  assign n72842 = ~n72852;
  assign n72837 = ~n72843;
  assign n72845 = n72867 & n72868;
  assign n72851 = ~n72875;
  assign n72856 = n185 ^ n72878;
  assign n72897 = ~n72914;
  assign n72903 = n72930 & n72931;
  assign n72787 = n72817 ^ n72818;
  assign n72805 = n72824 ^ n72825;
  assign n72829 = ~n72824;
  assign n72834 = n72836 & n72837;
  assign n72773 = n72841 & n72842;
  assign n72823 = n72845 ^ n70491;
  assign n72790 = n72855 ^ n72856;
  assign n72850 = ~n72845;
  assign n72839 = n72856 & n72858;
  assign n72887 = n72896 & n72897;
  assign n72873 = n184 ^ n72903;
  assign n72778 = n193 ^ n72805;
  assign n72797 = n72787 & n8358;
  assign n72801 = ~n72787;
  assign n68920 = n72822 ^ n72823;
  assign n72819 = n72828 & n72829;
  assign n72783 = ~n72773;
  assign n72815 = ~n72834;
  assign n72835 = n72790 & n70407;
  assign n72833 = ~n72790;
  assign n72840 = n72850 & n72851;
  assign n72814 = n72873 ^ n72874;
  assign n72864 = ~n72887;
  assign n70828 = n72777 ^ n72778;
  assign n72784 = ~n72797;
  assign n72779 = ~n72778;
  assign n72792 = n72801 & n192;
  assign n72810 = n68920 & n70514;
  assign n72798 = n72815 & n72816;
  assign n68947 = ~n68920;
  assign n72806 = ~n72819;
  assign n72830 = n72833 & n70430;
  assign n72789 = ~n72835;
  assign n72820 = ~n72840;
  assign n72838 = n72864 & n72865;
  assign n72269 = ~n70828;
  assign n72750 = n72779 & n72777;
  assign n72768 = ~n72792;
  assign n72774 = n72798 ^ n72799;
  assign n72802 = n68947 & n71524;
  assign n72786 = n72806 & n72807;
  assign n72796 = n72798 & n72808;
  assign n72781 = ~n72810;
  assign n72803 = ~n72798;
  assign n72809 = n72820 & n72821;
  assign n72812 = ~n72830;
  assign n72813 = n72838 ^ n72839;
  assign n72741 = n72773 ^ n72774;
  assign n72769 = n72786 ^ n72787;
  assign n72782 = ~n72796;
  assign n72780 = ~n72802;
  assign n72785 = ~n72786;
  assign n72793 = n72803 & n72799;
  assign n72791 = n72809 ^ n70407;
  assign n72811 = ~n72809;
  assign n72757 = n72813 ^ n72814;
  assign n72751 = n192 ^ n72769;
  assign n72734 = n72780 & n72781;
  assign n72776 = n72782 & n72783;
  assign n72775 = n72784 & n72785;
  assign n68880 = n72790 ^ n72791;
  assign n72766 = ~n72793;
  assign n72795 = n72757 & n70313;
  assign n72800 = n72811 & n72812;
  assign n72804 = ~n72757;
  assign n72212 = n72750 ^ n72751;
  assign n72720 = n72751 & n72750;
  assign n72772 = n68880 & n71469;
  assign n68878 = ~n68880;
  assign n72767 = ~n72775;
  assign n72743 = ~n72734;
  assign n72765 = ~n72776;
  assign n72755 = ~n72795;
  assign n72788 = ~n72800;
  assign n72794 = n72804 & n70340;
  assign n72199 = ~n72212;
  assign n72748 = n72765 & n72766;
  assign n72756 = n72767 & n72768;
  assign n72752 = ~n72772;
  assign n72763 = n68878 & n70407;
  assign n72764 = n72788 & n72789;
  assign n72771 = ~n72794;
  assign n72735 = n72748 ^ n72749;
  assign n72738 = n72756 ^ n72741;
  assign n72759 = n72756 & n8317;
  assign n72760 = n72748 & n72749;
  assign n72746 = ~n72748;
  assign n72761 = ~n72756;
  assign n72753 = ~n72763;
  assign n72758 = n72764 ^ n70313;
  assign n72770 = ~n72764;
  assign n72708 = n72734 ^ n72735;
  assign n72721 = n207 ^ n72738;
  assign n72745 = n72746 & n72747;
  assign n72688 = n72752 & n72753;
  assign n68823 = n72757 ^ n72758;
  assign n72740 = ~n72759;
  assign n72742 = ~n72760;
  assign n72744 = n72761 & n207;
  assign n72762 = n72770 & n72771;
  assign n70709 = n72720 ^ n72721;
  assign n72695 = ~n72708;
  assign n72722 = ~n72721;
  assign n72739 = n68823 & n71434;
  assign n72737 = n72740 & n72741;
  assign n72736 = n72742 & n72743;
  assign n68845 = ~n68823;
  assign n72728 = ~n72744;
  assign n72692 = ~n72688;
  assign n72726 = ~n72745;
  assign n72754 = ~n72762;
  assign n72152 = ~n70709;
  assign n72672 = n72722 & n72720;
  assign n72729 = n68845 & n70313;
  assign n72725 = ~n72736;
  assign n72727 = ~n72737;
  assign n72717 = ~n72739;
  assign n72731 = n72754 & n72755;
  assign n72671 = ~n72672;
  assign n72709 = n72725 & n72726;
  assign n72707 = n72727 & n72728;
  assign n72716 = ~n72729;
  assign n72724 = n72731 ^ n70216;
  assign n72732 = ~n72731;
  assign n72686 = n72707 ^ n72708;
  assign n72689 = n72709 ^ n72710;
  assign n72711 = n72709 & n72715;
  assign n72713 = n72707 & n8278;
  assign n72712 = ~n72709;
  assign n72650 = n72716 & n72717;
  assign n72706 = ~n72707;
  assign n68786 = n72723 ^ n72724;
  assign n72730 = n72732 & n72733;
  assign n72673 = n206 ^ n72686;
  assign n72654 = n72688 ^ n72689;
  assign n72703 = n72706 & n206;
  assign n72691 = ~n72711;
  assign n72699 = n68786 & n71372;
  assign n72702 = n72712 & n72710;
  assign n72694 = ~n72713;
  assign n72704 = n72650 & n72714;
  assign n72700 = ~n72650;
  assign n68814 = ~n68786;
  assign n72718 = ~n72730;
  assign n70627 = n72672 ^ n72673;
  assign n72670 = ~n72673;
  assign n72687 = n72691 & n72692;
  assign n72690 = n72694 & n72695;
  assign n72684 = ~n72699;
  assign n72697 = n72700 & n72665;
  assign n72680 = ~n72702;
  assign n72678 = ~n72703;
  assign n72669 = ~n72704;
  assign n72693 = n68814 & n70252;
  assign n72705 = n72718 & n72719;
  assign n72079 = ~n70627;
  assign n72629 = n72670 & n72671;
  assign n72679 = ~n72687;
  assign n72677 = ~n72690;
  assign n72683 = ~n72693;
  assign n72647 = ~n72697;
  assign n72701 = n72705 & n70166;
  assign n72698 = ~n72705;
  assign n72661 = n72677 & n72678;
  assign n72664 = n72679 & n72680;
  assign n72613 = n72683 & n72684;
  assign n72696 = n72698 & n70144;
  assign n72681 = ~n72701;
  assign n72652 = n72661 ^ n72654;
  assign n72651 = n72664 ^ n72665;
  assign n72662 = n72661 & n8239;
  assign n72668 = ~n72664;
  assign n72663 = ~n72661;
  assign n72617 = ~n72613;
  assign n72682 = n72681 & n72685;
  assign n72675 = ~n72696;
  assign n72621 = n72650 ^ n72651;
  assign n72630 = n205 ^ n72652;
  assign n72653 = ~n72662;
  assign n72657 = n72663 & n205;
  assign n72656 = n72668 & n72669;
  assign n72676 = n72675 & n72681;
  assign n72674 = ~n72682;
  assign n70506 = n72629 ^ n72630;
  assign n72632 = n72621 & n204;
  assign n72585 = n72630 & n72629;
  assign n72628 = ~n72621;
  assign n72648 = n72653 & n72654;
  assign n72646 = ~n72656;
  assign n72640 = ~n72657;
  assign n72658 = n72674 & n72675;
  assign n72667 = ~n72676;
  assign n71988 = ~n70506;
  assign n72627 = n72628 & n8227;
  assign n72595 = ~n72632;
  assign n72579 = ~n72585;
  assign n72635 = n72646 & n72647;
  assign n72639 = ~n72648;
  assign n72641 = n72658 ^ n70058;
  assign n68748 = n72666 ^ n72667;
  assign n72659 = ~n72658;
  assign n72611 = ~n72627;
  assign n72614 = n72635 ^ n72634;
  assign n72631 = n72635 & n72638;
  assign n72620 = n72639 & n72640;
  assign n68706 = n72641 ^ n72642;
  assign n72633 = ~n72635;
  assign n72649 = n68748 & n70144;
  assign n68780 = ~n68748;
  assign n72655 = n72659 & n72660;
  assign n72574 = n72613 ^ n72614;
  assign n72597 = n72620 ^ n72621;
  assign n72616 = ~n72631;
  assign n72612 = ~n72620;
  assign n72623 = n72633 & n72634;
  assign n72626 = n68706 & n71271;
  assign n68740 = ~n68706;
  assign n72645 = n68780 & n71343;
  assign n72636 = ~n72649;
  assign n72643 = ~n72655;
  assign n72596 = n72574 & n203;
  assign n72586 = n204 ^ n72597;
  assign n72593 = ~n72574;
  assign n72607 = n72611 & n72612;
  assign n72610 = n72616 & n72617;
  assign n72599 = ~n72623;
  assign n72605 = ~n72626;
  assign n72618 = n68740 & n70058;
  assign n72622 = n72643 & n72644;
  assign n72637 = ~n72645;
  assign n70428 = n72585 ^ n72586;
  assign n72592 = n72593 & n8167;
  assign n72578 = ~n72586;
  assign n72559 = ~n72596;
  assign n72594 = ~n72607;
  assign n72598 = ~n72610;
  assign n72606 = ~n72618;
  assign n72604 = n72622 ^ n69994;
  assign n72564 = n72636 & n72637;
  assign n72624 = ~n72622;
  assign n71917 = ~n70428;
  assign n72535 = n72578 & n72579;
  assign n72576 = ~n72592;
  assign n72573 = n72594 & n72595;
  assign n72580 = n72598 & n72599;
  assign n68661 = n72603 ^ n72604;
  assign n72524 = n72605 & n72606;
  assign n72615 = n72564 & n72581;
  assign n72608 = ~n72564;
  assign n72619 = n72624 & n72625;
  assign n72560 = n72573 ^ n72574;
  assign n72565 = n72580 ^ n72581;
  assign n72575 = ~n72573;
  assign n72587 = n68661 & n71200;
  assign n72582 = ~n72580;
  assign n68695 = ~n68661;
  assign n72533 = ~n72524;
  assign n72600 = n72608 & n72609;
  assign n72583 = ~n72615;
  assign n72601 = ~n72619;
  assign n72537 = n203 ^ n72560;
  assign n72540 = n72564 ^ n72565;
  assign n72566 = n72575 & n72576;
  assign n72572 = n72582 & n72583;
  assign n72569 = ~n72587;
  assign n72584 = n68695 & n70020;
  assign n72563 = ~n72600;
  assign n72588 = n72601 & n72602;
  assign n70347 = n72535 ^ n72537;
  assign n72541 = n72540 & n8128;
  assign n72534 = ~n72537;
  assign n72542 = ~n72540;
  assign n72558 = ~n72566;
  assign n72562 = ~n72572;
  assign n72568 = ~n72584;
  assign n68621 = n72588 ^ n72589;
  assign n72590 = ~n72588;
  assign n71834 = ~n70347;
  assign n72506 = n72534 & n72535;
  assign n72528 = ~n72541;
  assign n72536 = n72542 & n202;
  assign n72539 = n72558 & n72559;
  assign n72543 = n72562 & n72563;
  assign n72484 = n72568 & n72569;
  assign n72567 = n68621 & n69904;
  assign n68658 = ~n68621;
  assign n72577 = n72590 & n72591;
  assign n72519 = ~n72536;
  assign n72521 = n72539 ^ n72540;
  assign n72525 = n72543 ^ n72544;
  assign n72529 = ~n72539;
  assign n72546 = n72543 & n72553;
  assign n72549 = n72484 & n72557;
  assign n72548 = ~n72543;
  assign n72556 = ~n72484;
  assign n72555 = ~n72567;
  assign n72561 = n68658 & n71127;
  assign n72570 = ~n72577;
  assign n72507 = n202 ^ n72521;
  assign n72501 = n72524 ^ n72525;
  assign n72522 = n72528 & n72529;
  assign n72532 = ~n72546;
  assign n72538 = n72548 & n72544;
  assign n72499 = ~n72549;
  assign n72547 = n72556 & n72496;
  assign n72554 = ~n72561;
  assign n72550 = n72570 & n72571;
  assign n70270 = n72506 ^ n72507;
  assign n72455 = n72507 & n72506;
  assign n72509 = n72501 & n201;
  assign n72511 = ~n72501;
  assign n72518 = ~n72522;
  assign n72523 = n72532 & n72533;
  assign n72515 = ~n72538;
  assign n72476 = ~n72547;
  assign n72527 = n72550 ^ n69888;
  assign n72413 = n72554 & n72555;
  assign n72551 = ~n72550;
  assign n71758 = ~n70270;
  assign n72468 = ~n72455;
  assign n72470 = ~n72509;
  assign n72505 = n72511 & n8107;
  assign n72500 = n72518 & n72519;
  assign n72514 = ~n72523;
  assign n68565 = n72526 ^ n72527;
  assign n72545 = n72551 & n72552;
  assign n72477 = n72500 ^ n72501;
  assign n72492 = ~n72505;
  assign n72491 = ~n72500;
  assign n72495 = n72514 & n72515;
  assign n72520 = n68565 & n69893;
  assign n68622 = ~n68565;
  assign n72530 = ~n72545;
  assign n72456 = n201 ^ n72477;
  assign n72488 = n72491 & n72492;
  assign n72485 = n72495 ^ n72496;
  assign n72498 = ~n72495;
  assign n72494 = ~n72520;
  assign n72510 = n68622 & n71098;
  assign n72512 = n72530 & n72531;
  assign n70178 = n72455 ^ n72456;
  assign n72415 = n72456 & n72468;
  assign n72452 = n72484 ^ n72485;
  assign n72469 = ~n72488;
  assign n72490 = n72498 & n72499;
  assign n72493 = ~n72510;
  assign n72497 = n72512 ^ n72513;
  assign n72516 = ~n72512;
  assign n72418 = ~n72415;
  assign n72457 = n72452 & n200;
  assign n72451 = n72469 & n72470;
  assign n72453 = ~n72452;
  assign n72475 = ~n72490;
  assign n72410 = n72493 & n72494;
  assign n68543 = n69831 ^ n72497;
  assign n72502 = ~n72497;
  assign n72508 = n72516 & n72517;
  assign n72434 = n72451 ^ n72452;
  assign n72448 = n72453 & n8067;
  assign n72420 = ~n72457;
  assign n72438 = ~n72451;
  assign n72466 = n72475 & n72476;
  assign n72480 = n68543 & n72486;
  assign n72479 = n68543 & n70999;
  assign n72478 = n72410 & n72487;
  assign n72474 = ~n72410;
  assign n68574 = ~n68543;
  assign n72489 = n72502 & n69839;
  assign n72503 = ~n72508;
  assign n72416 = n200 ^ n72434;
  assign n72437 = ~n72448;
  assign n72454 = n72466 & n72467;
  assign n72458 = ~n72466;
  assign n72471 = n72474 & n72387;
  assign n72473 = n68574 & n71160;
  assign n72412 = ~n72478;
  assign n72464 = ~n72479;
  assign n71186 = ~n72480;
  assign n72465 = ~n72489;
  assign n72481 = n72503 & n72504;
  assign n72394 = n72415 ^ n72416;
  assign n72417 = ~n72416;
  assign n72429 = n72437 & n72438;
  assign n72436 = ~n72454;
  assign n72449 = n72458 & n72459;
  assign n72342 = n72464 & n72465;
  assign n72384 = ~n72471;
  assign n71165 = ~n72473;
  assign n72463 = n72481 ^ n69781;
  assign n72482 = ~n72481;
  assign n68287 = n72394 ^ n69342;
  assign n72273 = n72394 & n69344;
  assign n72388 = ~n72394;
  assign n72345 = n72417 & n72418;
  assign n72419 = ~n72429;
  assign n72435 = n72436 & n72413;
  assign n72428 = ~n72449;
  assign n72447 = n72342 & n72450;
  assign n68496 = n72462 ^ n72463;
  assign n72446 = ~n72342;
  assign n72472 = n72482 & n72483;
  assign n72373 = n68287 & n71284;
  assign n68277 = ~n68287;
  assign n72385 = n72388 & n69344;
  assign n72389 = n72419 & n72420;
  assign n72427 = ~n72435;
  assign n72432 = n72428 & n72436;
  assign n72439 = n68496 & n72445;
  assign n72441 = n72446 & n72364;
  assign n72440 = n68496 & n71005;
  assign n72368 = ~n72447;
  assign n68504 = ~n68496;
  assign n72460 = ~n72472;
  assign n72361 = ~n72373;
  assign n72362 = ~n72385;
  assign n72375 = ~n72389;
  assign n72409 = n72427 & n72428;
  assign n72414 = ~n72432;
  assign n71136 = ~n72439;
  assign n72422 = ~n72440;
  assign n72339 = ~n72441;
  assign n72433 = n68504 & n71104;
  assign n72430 = n68504 & n69793;
  assign n72442 = n72460 & n72461;
  assign n72330 = n72361 & n72362;
  assign n72386 = n72409 ^ n72410;
  assign n72390 = n72413 ^ n72414;
  assign n72411 = ~n72409;
  assign n72421 = ~n72430;
  assign n71109 = ~n72433;
  assign n72426 = n72442 ^ n69745;
  assign n72443 = ~n72442;
  assign n72299 = n72330 ^ n72331;
  assign n72332 = ~n72330;
  assign n72334 = n72386 ^ n72387;
  assign n72370 = n72389 ^ n72390;
  assign n72396 = n72390 & n8015;
  assign n72392 = ~n72390;
  assign n72398 = n72411 & n72412;
  assign n72290 = n72421 & n72422;
  assign n68450 = n72425 ^ n72426;
  assign n72431 = n72443 & n72444;
  assign n69708 = n231 ^ n72299;
  assign n72302 = ~n72299;
  assign n72124 = n72332 & n72331;
  assign n72346 = n215 ^ n72370;
  assign n72365 = n72334 & n214;
  assign n72366 = ~n72334;
  assign n72382 = n72392 & n215;
  assign n72374 = ~n72396;
  assign n72383 = ~n72398;
  assign n72404 = n68450 & n71077;
  assign n72408 = n68450 & n69745;
  assign n72399 = n72290 & n72316;
  assign n68494 = ~n68450;
  assign n72402 = ~n72290;
  assign n72423 = ~n72431;
  assign n71984 = ~n69708;
  assign n72018 = n72302 & n231;
  assign n72337 = n72345 ^ n72346;
  assign n72279 = n72346 & n72345;
  assign n72304 = ~n72365;
  assign n72355 = n72366 & n7981;
  assign n72372 = n72374 & n72375;
  assign n72354 = ~n72382;
  assign n72363 = n72383 & n72384;
  assign n72322 = ~n72399;
  assign n72397 = n72402 & n72403;
  assign n71043 = ~n72404;
  assign n72395 = n68494 & n72407;
  assign n72393 = n68494 & n70941;
  assign n72377 = ~n72408;
  assign n72400 = n72423 & n72424;
  assign n72324 = n72337 & n69260;
  assign n72325 = ~n72337;
  assign n72326 = ~n72355;
  assign n72343 = n72363 ^ n72364;
  assign n72353 = ~n72372;
  assign n72367 = ~n72363;
  assign n72378 = ~n72393;
  assign n71068 = ~n72395;
  assign n72293 = ~n72397;
  assign n72381 = n72400 ^ n72401;
  assign n72405 = ~n72400;
  assign n72275 = ~n72324;
  assign n72317 = n72325 & n69266;
  assign n72282 = n72342 ^ n72343;
  assign n72333 = n72353 & n72354;
  assign n72357 = n72367 & n72368;
  assign n72236 = n72377 & n72378;
  assign n68405 = n69690 ^ n72381;
  assign n72376 = ~n72381;
  assign n72391 = n72405 & n72406;
  assign n72296 = ~n72317;
  assign n72314 = n72282 & n213;
  assign n72318 = ~n72282;
  assign n72312 = n72333 ^ n72334;
  assign n72327 = ~n72333;
  assign n72338 = ~n72357;
  assign n72352 = n68405 & n70859;
  assign n72360 = n68405 & n72369;
  assign n72349 = n72236 & n72268;
  assign n72358 = ~n72236;
  assign n68411 = ~n68405;
  assign n72371 = n72376 & n69707;
  assign n72379 = ~n72391;
  assign n72294 = n72296 & n72273;
  assign n72272 = n72296 & n72275;
  assign n72280 = n214 ^ n72312;
  assign n72262 = ~n72314;
  assign n72300 = n72318 & n7930;
  assign n72323 = n72326 & n72327;
  assign n72315 = n72338 & n72339;
  assign n72266 = ~n72349;
  assign n72340 = ~n72352;
  assign n72347 = n68411 & n70958;
  assign n72344 = n72358 & n72359;
  assign n71007 = ~n72360;
  assign n72341 = ~n72371;
  assign n72356 = n72379 & n72380;
  assign n68251 = n72272 ^ n72273;
  assign n72218 = n72279 ^ n72280;
  assign n72274 = ~n72294;
  assign n72283 = ~n72280;
  assign n72284 = ~n72300;
  assign n72291 = n72315 ^ n72316;
  assign n72303 = ~n72323;
  assign n72321 = ~n72315;
  assign n72180 = n72340 & n72341;
  assign n72241 = ~n72344;
  assign n70963 = ~n72347;
  assign n72336 = n72356 ^ n69656;
  assign n72350 = ~n72356;
  assign n72249 = n68251 & n69260;
  assign n68262 = ~n68251;
  assign n72250 = n72218 & n69191;
  assign n72244 = n72274 & n72275;
  assign n72263 = ~n72218;
  assign n72231 = n72283 & n72279;
  assign n72224 = n72290 ^ n72291;
  assign n72281 = n72303 & n72304;
  assign n72308 = n72321 & n72322;
  assign n72313 = n72180 & n72217;
  assign n72319 = ~n72180;
  assign n68354 = n72335 ^ n72336;
  assign n72348 = n72350 & n72351;
  assign n72219 = n72244 ^ n69191;
  assign n72242 = n68262 & n71172;
  assign n72221 = ~n72249;
  assign n72238 = ~n72250;
  assign n72246 = n72263 & n69218;
  assign n72239 = ~n72244;
  assign n72271 = n72224 & n7900;
  assign n72270 = ~n72224;
  assign n72264 = n72281 ^ n72282;
  assign n72285 = ~n72281;
  assign n72292 = ~n72308;
  assign n72215 = ~n72313;
  assign n72307 = n68354 & n70893;
  assign n72306 = n72319 & n72320;
  assign n72301 = n68354 & n69653;
  assign n68415 = ~n68354;
  assign n72328 = ~n72348;
  assign n68068 = n72218 ^ n72219;
  assign n72235 = n72238 & n72239;
  assign n72222 = ~n72242;
  assign n72210 = ~n72246;
  assign n72232 = n72264 ^ n7930;
  assign n72253 = n72270 & n212;
  assign n72229 = ~n72271;
  assign n72276 = n72284 & n72285;
  assign n72267 = n72292 & n72293;
  assign n72277 = ~n72301;
  assign n72178 = ~n72306;
  assign n70898 = ~n72307;
  assign n72298 = n68415 & n72311;
  assign n72295 = n68415 & n70682;
  assign n72305 = n72328 & n72329;
  assign n72189 = n68068 & n71118;
  assign n68083 = ~n68068;
  assign n72200 = n72221 & n72222;
  assign n72156 = n72231 ^ n72232;
  assign n72209 = ~n72235;
  assign n72168 = n72232 & n72231;
  assign n72195 = ~n72253;
  assign n72237 = n72267 ^ n72268;
  assign n72261 = ~n72276;
  assign n72265 = ~n72267;
  assign n72278 = ~n72295;
  assign n70926 = ~n72298;
  assign n72287 = n72305 ^ n69600;
  assign n72309 = ~n72305;
  assign n72176 = n68083 & n69218;
  assign n72161 = ~n72189;
  assign n72185 = n72200 & n72201;
  assign n72190 = ~n72200;
  assign n72182 = n72209 & n72210;
  assign n72165 = n72236 ^ n72237;
  assign n72223 = n72261 & n72262;
  assign n72255 = n72265 & n72266;
  assign n72114 = n72277 & n72278;
  assign n68315 = n72286 ^ n72287;
  assign n72297 = n72309 & n72310;
  assign n72160 = ~n72176;
  assign n72158 = n72182 ^ n72156;
  assign n72179 = n72182 & n69172;
  assign n72159 = ~n72185;
  assign n72175 = n72190 & n72191;
  assign n72183 = ~n72182;
  assign n72213 = n72165 & n7845;
  assign n72202 = n72223 ^ n72224;
  assign n72211 = ~n72165;
  assign n72230 = ~n72223;
  assign n72240 = ~n72255;
  assign n72254 = n68315 & n69614;
  assign n72257 = n68315 & n72269;
  assign n72260 = n72114 & n72146;
  assign n68320 = ~n68315;
  assign n72258 = ~n72114;
  assign n72288 = ~n72297;
  assign n72147 = n72158 & n69170;
  assign n72065 = n72160 & n72161;
  assign n72157 = n72159 & n72124;
  assign n72135 = ~n72158;
  assign n72134 = ~n72175;
  assign n72155 = ~n72179;
  assign n72170 = n72183 & n69170;
  assign n72169 = n212 ^ n72202;
  assign n72196 = n72211 & n211;
  assign n72172 = ~n72213;
  assign n72220 = n72229 & n72230;
  assign n72216 = n72240 & n72241;
  assign n72243 = n68320 & n70828;
  assign n72226 = ~n72254;
  assign n70826 = ~n72257;
  assign n72245 = n72258 & n72259;
  assign n72150 = ~n72260;
  assign n72247 = n68320 & n70696;
  assign n72256 = n72288 & n72289;
  assign n68013 = n72135 ^ n69170;
  assign n72126 = n72065 & n72098;
  assign n72059 = ~n72147;
  assign n72116 = ~n72065;
  assign n72151 = n72155 & n72156;
  assign n72133 = ~n72157;
  assign n72123 = n72134 & n72159;
  assign n72047 = n72168 ^ n72169;
  assign n72122 = ~n72170;
  assign n72101 = n72169 & n72168;
  assign n72140 = ~n72196;
  assign n72181 = n72216 ^ n72217;
  assign n72194 = ~n72220;
  assign n72214 = ~n72216;
  assign n70854 = ~n72243;
  assign n72113 = ~n72245;
  assign n72225 = ~n72247;
  assign n72234 = n72256 ^ n69544;
  assign n72251 = ~n72256;
  assign n72111 = n72116 & n72117;
  assign n67991 = ~n68013;
  assign n72094 = n72123 ^ n72124;
  assign n72099 = ~n72126;
  assign n72097 = n72133 & n72134;
  assign n72137 = n72047 & n69115;
  assign n72121 = ~n72151;
  assign n72128 = ~n72047;
  assign n72104 = ~n72101;
  assign n72093 = n72180 ^ n72181;
  assign n72164 = n72194 & n72195;
  assign n72197 = n72214 & n72215;
  assign n72039 = n72225 & n72226;
  assign n68212 = n72233 ^ n72234;
  assign n72248 = n72251 & n72252;
  assign n72088 = n72094 & n230;
  assign n72086 = n67991 & n71030;
  assign n72066 = n72097 ^ n72098;
  assign n72055 = ~n72111;
  assign n72091 = ~n72094;
  assign n72100 = ~n72097;
  assign n72090 = n72121 & n72122;
  assign n72127 = n72128 & n69131;
  assign n72052 = ~n72137;
  assign n72153 = n72093 & n7794;
  assign n72148 = ~n72093;
  assign n72136 = n72164 ^ n72165;
  assign n72171 = ~n72164;
  assign n72177 = ~n72197;
  assign n72203 = n68212 & n69581;
  assign n72198 = n68212 & n72212;
  assign n72204 = n72039 & n72075;
  assign n68336 = ~n68212;
  assign n72192 = ~n72039;
  assign n72227 = ~n72248;
  assign n71979 = n72065 ^ n72066;
  assign n72058 = ~n72086;
  assign n72015 = ~n72088;
  assign n72048 = n72090 ^ n69115;
  assign n72080 = n72091 & n19809;
  assign n72087 = n72099 & n72100;
  assign n72084 = ~n72090;
  assign n72085 = ~n72127;
  assign n72102 = n211 ^ n72136;
  assign n72132 = n72148 & n210;
  assign n72108 = ~n72153;
  assign n72154 = n72171 & n72172;
  assign n72145 = n72177 & n72178;
  assign n72184 = n72192 & n72193;
  assign n70736 = ~n72198;
  assign n72186 = n68336 & n72199;
  assign n72167 = ~n72203;
  assign n72083 = ~n72204;
  assign n72187 = n68336 & n70656;
  assign n72205 = n72227 & n72228;
  assign n72036 = n71979 & n19742;
  assign n67937 = n72047 ^ n72048;
  assign n72023 = ~n71979;
  assign n71980 = n72058 & n72059;
  assign n72046 = ~n72080;
  assign n72078 = n72084 & n72085;
  assign n72054 = ~n72087;
  assign n71973 = n72101 ^ n72102;
  assign n72103 = ~n72102;
  assign n72063 = ~n72132;
  assign n72115 = n72145 ^ n72146;
  assign n72139 = ~n72154;
  assign n72149 = ~n72145;
  assign n72043 = ~n72184;
  assign n70779 = ~n72186;
  assign n72166 = ~n72187;
  assign n72163 = n72205 ^ n72206;
  assign n72207 = ~n72205;
  assign n72012 = n67937 & n70934;
  assign n72016 = n72023 & n229;
  assign n71976 = ~n72036;
  assign n67930 = ~n67937;
  assign n72004 = ~n71980;
  assign n72041 = n72046 & n72018;
  assign n72017 = n72046 & n72015;
  assign n72028 = n72054 & n72055;
  assign n72064 = n71973 & n69094;
  assign n72051 = ~n72078;
  assign n72072 = ~n71973;
  assign n72021 = n72103 & n72104;
  assign n72031 = n72114 ^ n72115;
  assign n72092 = n72139 & n72140;
  assign n72141 = n72149 & n72150;
  assign n68191 = n69532 ^ n72163;
  assign n71999 = n72166 & n72167;
  assign n70790 = n70736 & n70779;
  assign n72162 = n72163 & n69517;
  assign n72188 = n72207 & n72208;
  assign n72000 = n67930 & n69115;
  assign n71966 = ~n72012;
  assign n71942 = ~n72016;
  assign n71975 = n72017 ^ n72018;
  assign n71981 = n72028 ^ n72029;
  assign n72033 = n72028 & n72029;
  assign n72014 = ~n72041;
  assign n72024 = ~n72028;
  assign n72013 = n72051 & n72052;
  assign n72009 = ~n72064;
  assign n72049 = n72072 & n69077;
  assign n72081 = n72031 & n7739;
  assign n72056 = n72092 ^ n72093;
  assign n72077 = ~n72031;
  assign n72107 = ~n72092;
  assign n72112 = ~n72141;
  assign n72142 = n68191 & n72152;
  assign n72138 = n71999 & n71958;
  assign n68196 = ~n68191;
  assign n72130 = ~n71999;
  assign n72106 = ~n72162;
  assign n72173 = ~n72188;
  assign n69676 = n71975 ^ n69708;
  assign n71859 = n71980 ^ n71981;
  assign n71888 = n71975 & n71984;
  assign n71967 = ~n72000;
  assign n71974 = n72013 ^ n69077;
  assign n71978 = n72014 & n72015;
  assign n72011 = n72024 & n72025;
  assign n72003 = ~n72033;
  assign n72010 = ~n72013;
  assign n71970 = ~n72049;
  assign n72022 = n210 ^ n72056;
  assign n72057 = n72077 & n209;
  assign n72027 = ~n72081;
  assign n72089 = n72107 & n72108;
  assign n72074 = n72112 & n72113;
  assign n72118 = n68196 & n70441;
  assign n72125 = n68196 & n70709;
  assign n72120 = n72130 & n72131;
  assign n72007 = ~n72138;
  assign n70674 = ~n72142;
  assign n72129 = n72173 & n72174;
  assign n71946 = n71859 & n19716;
  assign n70805 = ~n69676;
  assign n71880 = n71966 & n71967;
  assign n71943 = ~n71859;
  assign n67852 = n71973 ^ n71974;
  assign n71932 = n71978 ^ n71979;
  assign n71977 = ~n71978;
  assign n71990 = n72003 & n72004;
  assign n72001 = n72009 & n72010;
  assign n71962 = ~n72011;
  assign n71916 = n72021 ^ n72022;
  assign n72032 = ~n72022;
  assign n71992 = ~n72057;
  assign n72040 = n72074 ^ n72075;
  assign n72062 = ~n72089;
  assign n72082 = ~n72074;
  assign n72105 = ~n72118;
  assign n71960 = ~n72120;
  assign n70715 = ~n72125;
  assign n72110 = n72129 ^ n69467;
  assign n72143 = ~n72129;
  assign n71889 = n229 ^ n71932;
  assign n71935 = n71943 & n228;
  assign n71890 = ~n71946;
  assign n71939 = n71880 & n71928;
  assign n71936 = n67852 & n69077;
  assign n67876 = ~n67852;
  assign n71933 = ~n71880;
  assign n71964 = n71976 & n71977;
  assign n71961 = ~n71990;
  assign n71969 = ~n72001;
  assign n71944 = n72032 & n72021;
  assign n71950 = n72039 ^ n72040;
  assign n72030 = n72062 & n72063;
  assign n72068 = n72082 & n72083;
  assign n71877 = n72105 & n72106;
  assign n68111 = n72109 ^ n72110;
  assign n72119 = n72143 & n72144;
  assign n69631 = n71888 ^ n71889;
  assign n71819 = n71889 & n71888;
  assign n71920 = n71933 & n71934;
  assign n71855 = ~n71935;
  assign n71897 = ~n71936;
  assign n71922 = n67876 & n70851;
  assign n71918 = ~n71939;
  assign n71927 = n71961 & n71962;
  assign n71941 = ~n71964;
  assign n71938 = n71969 & n71970;
  assign n71963 = ~n71944;
  assign n72005 = n71950 & n7684;
  assign n72002 = ~n71950;
  assign n71989 = n72030 ^ n72031;
  assign n72026 = ~n72030;
  assign n72042 = ~n72068;
  assign n72061 = n71877 & n72076;
  assign n72060 = n68111 & n69467;
  assign n72067 = n68111 & n72079;
  assign n68233 = ~n68111;
  assign n72073 = ~n71877;
  assign n72095 = ~n72119;
  assign n70766 = ~n69631;
  assign n71861 = ~n71920;
  assign n71896 = ~n71922;
  assign n71881 = n71927 ^ n71928;
  assign n71899 = n71938 ^ n71916;
  assign n71885 = n71941 & n71942;
  assign n71940 = n71938 & n69039;
  assign n71919 = ~n71927;
  assign n71937 = ~n71938;
  assign n71945 = n209 ^ n71989;
  assign n71982 = n72002 & n208;
  assign n71948 = ~n72005;
  assign n72008 = n72026 & n72027;
  assign n71998 = n72042 & n72043;
  assign n72035 = ~n72060;
  assign n71924 = ~n72061;
  assign n70577 = ~n72067;
  assign n72050 = n68233 & n70296;
  assign n72044 = n68233 & n70627;
  assign n72045 = n72073 & n71926;
  assign n72069 = n72095 & n72096;
  assign n71816 = n71880 ^ n71881;
  assign n71858 = n228 ^ n71885;
  assign n71799 = n71896 & n71897;
  assign n67782 = n69039 ^ n71899;
  assign n71895 = n71899 & n69048;
  assign n71898 = n71918 & n71919;
  assign n71891 = ~n71885;
  assign n71930 = n71937 & n69048;
  assign n71915 = ~n71940;
  assign n71795 = n71944 ^ n71945;
  assign n71866 = n71945 & n71963;
  assign n71907 = ~n71982;
  assign n71957 = n71998 ^ n71999;
  assign n71991 = ~n72008;
  assign n72006 = ~n71998;
  assign n70625 = ~n72044;
  assign n71883 = ~n72045;
  assign n72034 = ~n72050;
  assign n72038 = n72069 ^ n69427;
  assign n72070 = ~n72069;
  assign n71852 = n71816 & n19695;
  assign n71820 = n71858 ^ n71859;
  assign n71851 = ~n71816;
  assign n71853 = n71799 & n71872;
  assign n67796 = ~n67782;
  assign n71857 = ~n71799;
  assign n71879 = n71890 & n71891;
  assign n71809 = ~n71895;
  assign n71860 = ~n71898;
  assign n71887 = n71915 & n71916;
  assign n71910 = n71795 & n68999;
  assign n71874 = ~n71930;
  assign n71900 = ~n71795;
  assign n71876 = n71957 ^ n71958;
  assign n71949 = n71991 & n71992;
  assign n71994 = n72006 & n72007;
  assign n71801 = n72034 & n72035;
  assign n68036 = n72037 ^ n72038;
  assign n72053 = n72070 & n72071;
  assign n69620 = n71819 ^ n71820;
  assign n71745 = n71820 & n71819;
  assign n71826 = n71851 & n227;
  assign n71811 = ~n71852;
  assign n71829 = ~n71853;
  assign n71845 = n71857 & n71828;
  assign n71850 = n67796 & n70743;
  assign n71827 = n71860 & n71861;
  assign n71854 = ~n71879;
  assign n71873 = ~n71887;
  assign n71886 = n71900 & n69008;
  assign n71825 = ~n71910;
  assign n71921 = n71876 & n7559;
  assign n71929 = ~n71876;
  assign n71908 = n71949 ^ n71950;
  assign n71947 = ~n71949;
  assign n71959 = ~n71994;
  assign n71997 = n68036 & n70506;
  assign n71987 = n68036 & n70257;
  assign n71983 = n71801 & n71849;
  assign n68038 = ~n68036;
  assign n71985 = ~n71801;
  assign n72019 = ~n72053;
  assign n70620 = ~n69620;
  assign n71780 = ~n71826;
  assign n71800 = n71827 ^ n71828;
  assign n71784 = ~n71845;
  assign n71808 = ~n71850;
  assign n71815 = n71854 & n71855;
  assign n71830 = ~n71827;
  assign n71840 = n71873 & n71874;
  assign n71798 = ~n71886;
  assign n71867 = n208 ^ n71908;
  assign n71869 = ~n71921;
  assign n71905 = n71929 & n223;
  assign n71931 = n71947 & n71948;
  assign n71925 = n71959 & n71960;
  assign n71965 = n68038 & n69472;
  assign n71842 = ~n71983;
  assign n71972 = n71985 & n71986;
  assign n71952 = ~n71987;
  assign n71971 = n68038 & n71988;
  assign n70543 = ~n71997;
  assign n71993 = n72019 & n72020;
  assign n71742 = n71799 ^ n71800;
  assign n71723 = n71808 & n71809;
  assign n71782 = n71815 ^ n71816;
  assign n71814 = n71829 & n71830;
  assign n71796 = n71840 ^ n68999;
  assign n71812 = ~n71815;
  assign n71824 = ~n71840;
  assign n71718 = n71866 ^ n71867;
  assign n71793 = n71867 & n71866;
  assign n71839 = ~n71905;
  assign n71878 = n71925 ^ n71926;
  assign n71906 = ~n71931;
  assign n71923 = ~n71925;
  assign n71951 = ~n71965;
  assign n70509 = ~n71971;
  assign n71805 = ~n71972;
  assign n71954 = n71993 ^ n69381;
  assign n71995 = ~n71993;
  assign n71766 = n71742 & n226;
  assign n71767 = ~n71742;
  assign n71746 = n227 ^ n71782;
  assign n67720 = n71795 ^ n71796;
  assign n71732 = ~n71723;
  assign n71803 = n71811 & n71812;
  assign n71783 = ~n71814;
  assign n71813 = n71824 & n71825;
  assign n71786 = n71877 ^ n71878;
  assign n71875 = n71906 & n71907;
  assign n71904 = n71923 & n71924;
  assign n71730 = n71951 & n71952;
  assign n67963 = n71953 ^ n71954;
  assign n71968 = n71995 & n71996;
  assign n69559 = n71745 ^ n71746;
  assign n71672 = n71746 & n71745;
  assign n71680 = ~n71766;
  assign n71740 = n71767 & n19641;
  assign n71752 = n67720 & n70634;
  assign n67747 = ~n67720;
  assign n71749 = n71783 & n71784;
  assign n71779 = ~n71803;
  assign n71797 = ~n71813;
  assign n71844 = n71786 & n222;
  assign n71843 = ~n71786;
  assign n71831 = n71875 ^ n71876;
  assign n71868 = ~n71875;
  assign n71882 = ~n71904;
  assign n71913 = n71730 & n71773;
  assign n71914 = n67963 & n70428;
  assign n71909 = n67963 & n69381;
  assign n71911 = ~n71730;
  assign n68127 = ~n67963;
  assign n71955 = ~n71968;
  assign n70550 = ~n69559;
  assign n71713 = ~n71740;
  assign n71724 = n71749 ^ n71750;
  assign n71725 = ~n71752;
  assign n71744 = n67747 & n69008;
  assign n71751 = n71749 & n71750;
  assign n71741 = n71779 & n71780;
  assign n71768 = ~n71749;
  assign n71747 = n71797 & n71798;
  assign n71794 = n223 ^ n71831;
  assign n71833 = n71843 & n7536;
  assign n71757 = ~n71844;
  assign n71856 = n71868 & n71869;
  assign n71848 = n71882 & n71883;
  assign n71871 = ~n71909;
  assign n71893 = n71911 & n71912;
  assign n71778 = ~n71913;
  assign n70427 = ~n71914;
  assign n71894 = n68127 & n71917;
  assign n71884 = n68127 & n70298;
  assign n71901 = n71955 & n71956;
  assign n71653 = n71723 ^ n71724;
  assign n71705 = n71741 ^ n71742;
  assign n71726 = ~n71744;
  assign n71719 = n71747 ^ n68963;
  assign n71733 = ~n71751;
  assign n71737 = n71768 & n71769;
  assign n71714 = ~n71741;
  assign n71755 = n71747 & n68963;
  assign n71763 = ~n71747;
  assign n71636 = n71793 ^ n71794;
  assign n71715 = n71794 & n71793;
  assign n71792 = ~n71833;
  assign n71802 = n71848 ^ n71849;
  assign n71838 = ~n71856;
  assign n71841 = ~n71848;
  assign n71870 = ~n71884;
  assign n71729 = ~n71893;
  assign n70471 = ~n71894;
  assign n71865 = n71901 ^ n69336;
  assign n71902 = ~n71901;
  assign n71673 = n226 ^ n71705;
  assign n71625 = ~n71653;
  assign n71706 = n71713 & n71714;
  assign n67678 = n71718 ^ n71719;
  assign n71632 = n71725 & n71726;
  assign n71720 = n71732 & n71733;
  assign n71702 = ~n71737;
  assign n71734 = ~n71755;
  assign n71735 = n71763 & n68972;
  assign n71765 = n71636 & n68920;
  assign n71748 = ~n71636;
  assign n71710 = n71801 ^ n71802;
  assign n71785 = n71838 & n71839;
  assign n71832 = n71841 & n71842;
  assign n67905 = n71864 ^ n71865;
  assign n71660 = n71870 & n71871;
  assign n71892 = n71902 & n71903;
  assign n69549 = n71672 ^ n71673;
  assign n71689 = n67678 & n68972;
  assign n71686 = n71632 & n71700;
  assign n71671 = ~n71673;
  assign n71688 = ~n71632;
  assign n67688 = ~n67678;
  assign n71679 = ~n71706;
  assign n71701 = ~n71720;
  assign n71717 = n71734 & n71718;
  assign n71699 = ~n71735;
  assign n71743 = n71748 & n68947;
  assign n71635 = ~n71765;
  assign n71775 = n71710 & n7384;
  assign n71754 = n71785 ^ n71786;
  assign n71776 = ~n71710;
  assign n71791 = ~n71785;
  assign n71804 = ~n71832;
  assign n71836 = n67905 & n70084;
  assign n71823 = n67905 & n70347;
  assign n71822 = n71660 & n71846;
  assign n67899 = ~n67905;
  assign n71835 = ~n71660;
  assign n71862 = ~n71892;
  assign n70464 = ~n69549;
  assign n71600 = n71671 & n71672;
  assign n71652 = n71679 & n71680;
  assign n71670 = n67688 & n70554;
  assign n71667 = ~n71686;
  assign n71669 = n71688 & n71663;
  assign n71645 = ~n71689;
  assign n71662 = n71701 & n71702;
  assign n71698 = ~n71717;
  assign n71659 = ~n71743;
  assign n71716 = n222 ^ n71754;
  assign n71712 = ~n71775;
  assign n71762 = n71776 & n221;
  assign n71781 = n71791 & n71792;
  assign n71772 = n71804 & n71805;
  assign n71810 = n67899 & n69336;
  assign n71691 = ~n71822;
  assign n70391 = ~n71823;
  assign n71817 = n67899 & n71834;
  assign n71818 = n71835 & n71696;
  assign n71789 = ~n71836;
  assign n71837 = n71862 & n71863;
  assign n71623 = n71652 ^ n71653;
  assign n71650 = n71652 & n19596;
  assign n71633 = n71662 ^ n71663;
  assign n71631 = ~n71669;
  assign n71646 = ~n71670;
  assign n71649 = ~n71652;
  assign n71668 = ~n71662;
  assign n71666 = n71698 & n71699;
  assign n71580 = n71715 ^ n71716;
  assign n71721 = ~n71716;
  assign n71678 = ~n71762;
  assign n71731 = n71772 ^ n71773;
  assign n71756 = ~n71781;
  assign n71777 = ~n71772;
  assign n71790 = ~n71810;
  assign n70351 = ~n71817;
  assign n71665 = ~n71818;
  assign n71788 = n71837 ^ n69297;
  assign n71821 = n71837 & n71847;
  assign n71601 = n225 ^ n71623;
  assign n71556 = n71632 ^ n71633;
  assign n71582 = n71645 & n71646;
  assign n71640 = n71649 & n225;
  assign n71624 = ~n71650;
  assign n71637 = n71666 ^ n68920;
  assign n71651 = n71667 & n71668;
  assign n71658 = ~n71666;
  assign n71683 = n71580 & n68880;
  assign n71685 = ~n71580;
  assign n71654 = n71721 & n71715;
  assign n71643 = n71730 ^ n71731;
  assign n71709 = n71756 & n71757;
  assign n71753 = n71777 & n71778;
  assign n67826 = n71787 ^ n71788;
  assign n71627 = n71789 & n71790;
  assign n71806 = ~n71821;
  assign n69479 = n71600 ^ n71601;
  assign n71513 = n71601 & n71600;
  assign n71619 = n71624 & n71625;
  assign n67628 = n71636 ^ n71637;
  assign n71588 = ~n71582;
  assign n71613 = ~n71640;
  assign n71630 = ~n71651;
  assign n71644 = n71658 & n71659;
  assign n71616 = ~n71683;
  assign n71675 = n71685 & n68878;
  assign n71697 = n71643 & n7394;
  assign n71682 = n71709 ^ n71710;
  assign n71703 = ~n71643;
  assign n71711 = ~n71709;
  assign n71728 = ~n71753;
  assign n71764 = n67826 & n70270;
  assign n71761 = n67826 & n69297;
  assign n71760 = n71627 & n71774;
  assign n67832 = ~n67826;
  assign n71759 = ~n71627;
  assign n71770 = n71806 & n71807;
  assign n70399 = ~n69479;
  assign n71611 = n67628 & n70514;
  assign n71612 = ~n71619;
  assign n67640 = ~n67628;
  assign n71607 = n71630 & n71631;
  assign n71634 = ~n71644;
  assign n71571 = ~n71675;
  assign n71655 = n221 ^ n71682;
  assign n71648 = ~n71697;
  assign n71684 = n71703 & n220;
  assign n71704 = n71711 & n71712;
  assign n71695 = n71728 & n71729;
  assign n71739 = n67832 & n70016;
  assign n71738 = n67832 & n71758;
  assign n71736 = n71759 & n71606;
  assign n71629 = ~n71760;
  assign n71708 = ~n71761;
  assign n70262 = ~n71764;
  assign n67957 = n71770 ^ n71771;
  assign n71595 = n67640 & n68920;
  assign n71583 = n71607 ^ n71608;
  assign n71585 = ~n71611;
  assign n71577 = n71612 & n71613;
  assign n71614 = n71607 & n71608;
  assign n71609 = ~n71607;
  assign n71604 = n71634 & n71635;
  assign n71518 = n71654 ^ n71655;
  assign n71596 = n71655 & n71654;
  assign n71621 = ~n71684;
  assign n71661 = n71695 ^ n71696;
  assign n71677 = ~n71704;
  assign n71690 = ~n71695;
  assign n71603 = ~n71736;
  assign n71727 = n67957 & n69315;
  assign n70303 = ~n71738;
  assign n71707 = ~n71739;
  assign n69368 = ~n67957;
  assign n71541 = n71577 ^ n71556;
  assign n71494 = n71582 ^ n71583;
  assign n71578 = n71577 & n19565;
  assign n71579 = ~n71577;
  assign n71584 = ~n71595;
  assign n71581 = n71604 ^ n68880;
  assign n71592 = n71609 & n71610;
  assign n71587 = ~n71614;
  assign n71615 = ~n71604;
  assign n71591 = ~n71596;
  assign n71565 = n71660 ^ n71661;
  assign n71642 = n71677 & n71678;
  assign n71676 = n71690 & n71691;
  assign n71575 = n71707 & n71708;
  assign n71722 = n69368 & n70079;
  assign n71694 = ~n71727;
  assign n71514 = n224 ^ n71541;
  assign n71546 = n71494 & n19533;
  assign n71548 = ~n71494;
  assign n71555 = ~n71578;
  assign n71563 = n71579 & n224;
  assign n67595 = n71580 ^ n71581;
  assign n71491 = n71584 & n71585;
  assign n71569 = n71587 & n71588;
  assign n71559 = ~n71592;
  assign n71598 = n71615 & n71616;
  assign n71639 = n71565 & n219;
  assign n71617 = n71642 ^ n71643;
  assign n71638 = ~n71565;
  assign n71647 = ~n71642;
  assign n71664 = ~n71676;
  assign n71687 = n71575 & n71692;
  assign n71681 = ~n71575;
  assign n71693 = ~n71722;
  assign n69459 = n71513 ^ n71514;
  assign n71517 = ~n71514;
  assign n71498 = ~n71546;
  assign n71530 = n71548 & n239;
  assign n71549 = n67595 & n70407;
  assign n71545 = n71555 & n71556;
  assign n71540 = n71491 & n71557;
  assign n71522 = ~n71563;
  assign n71550 = ~n71491;
  assign n67591 = ~n67595;
  assign n71558 = ~n71569;
  assign n71570 = ~n71598;
  assign n71597 = n220 ^ n71617;
  assign n71622 = n71638 & n7342;
  assign n71562 = ~n71639;
  assign n71641 = n71647 & n71648;
  assign n71626 = n71664 & n71665;
  assign n71674 = n71681 & n71553;
  assign n71573 = ~n71687;
  assign n71656 = n71693 & n71694;
  assign n70309 = ~n69459;
  assign n71439 = n71517 & n71513;
  assign n71467 = ~n71530;
  assign n71525 = ~n71540;
  assign n71521 = ~n71545;
  assign n71531 = n67591 & n68878;
  assign n71508 = ~n71549;
  assign n71532 = n71550 & n71524;
  assign n71523 = n71558 & n71559;
  assign n71551 = n71570 & n71571;
  assign n71441 = n71596 ^ n71597;
  assign n71590 = ~n71597;
  assign n71594 = ~n71622;
  assign n71605 = n71626 ^ n71627;
  assign n71620 = ~n71641;
  assign n71628 = ~n71626;
  assign n71487 = n71656 ^ n71657;
  assign n71544 = ~n71674;
  assign n71438 = ~n71439;
  assign n71493 = n71521 & n71522;
  assign n71492 = n71523 ^ n71524;
  assign n71509 = ~n71531;
  assign n71501 = ~n71532;
  assign n71526 = ~n71523;
  assign n71519 = n71551 ^ n68823;
  assign n71542 = n71551 & n68823;
  assign n71547 = ~n71551;
  assign n71560 = n71441 & n68786;
  assign n71566 = ~n71441;
  assign n71535 = n71590 & n71591;
  assign n71538 = n71605 ^ n71606;
  assign n71599 = n71620 & n71621;
  assign n71618 = n71628 & n71629;
  assign n71446 = n71491 ^ n71492;
  assign n71472 = n71493 ^ n71494;
  assign n71451 = n71508 & n71509;
  assign n71499 = ~n71493;
  assign n67545 = n71518 ^ n71519;
  assign n71515 = n71525 & n71526;
  assign n71520 = ~n71542;
  assign n71539 = n71547 & n68845;
  assign n71475 = ~n71560;
  assign n71554 = n71566 & n68814;
  assign n71586 = n71538 & n218;
  assign n71529 = ~n71535;
  assign n71576 = ~n71538;
  assign n71564 = n219 ^ n71599;
  assign n71593 = ~n71599;
  assign n71602 = ~n71618;
  assign n71440 = n239 ^ n71472;
  assign n71478 = n71446 & n238;
  assign n71473 = ~n71446;
  assign n71489 = n67545 & n68845;
  assign n71490 = n71498 & n71499;
  assign n67568 = ~n67545;
  assign n71459 = ~n71451;
  assign n71500 = ~n71515;
  assign n71510 = n71520 & n71518;
  assign n71497 = ~n71539;
  assign n71444 = ~n71554;
  assign n71536 = n71564 ^ n71565;
  assign n71567 = n71576 & n7252;
  assign n71505 = ~n71586;
  assign n71589 = n71593 & n71594;
  assign n71574 = n71602 & n71603;
  assign n69395 = n71439 ^ n71440;
  assign n71437 = ~n71440;
  assign n71461 = n71473 & n19483;
  assign n71416 = ~n71478;
  assign n71480 = n67568 & n70313;
  assign n71464 = ~n71489;
  assign n71466 = ~n71490;
  assign n71477 = n71500 & n71501;
  assign n71496 = ~n71510;
  assign n71395 = n71535 ^ n71536;
  assign n71528 = ~n71536;
  assign n71534 = ~n71567;
  assign n71552 = n71574 ^ n71575;
  assign n71561 = ~n71589;
  assign n71572 = ~n71574;
  assign n70234 = ~n69395;
  assign n70118 = n71437 & n71438;
  assign n71447 = ~n71461;
  assign n71445 = n71466 & n71467;
  assign n71452 = n71477 ^ n71469;
  assign n71463 = ~n71480;
  assign n71476 = n71477 & n71485;
  assign n71468 = ~n71477;
  assign n71470 = n71496 & n71497;
  assign n71507 = n71395 & n68748;
  assign n71502 = ~n71395;
  assign n71483 = n71528 & n71529;
  assign n71457 = n71552 ^ n71553;
  assign n71537 = n71561 & n71562;
  assign n71568 = n71572 & n71573;
  assign n71403 = ~n70118;
  assign n71417 = n71445 ^ n71446;
  assign n71392 = n71451 ^ n71452;
  assign n71386 = n71463 & n71464;
  assign n71448 = ~n71445;
  assign n71462 = n71468 & n71469;
  assign n71442 = n71470 ^ n68786;
  assign n71458 = ~n71476;
  assign n71474 = ~n71470;
  assign n71495 = n71502 & n68780;
  assign n71394 = ~n71507;
  assign n71488 = ~n71483;
  assign n71512 = n71457 & n217;
  assign n71516 = ~n71457;
  assign n71506 = n71537 ^ n71538;
  assign n71533 = ~n71537;
  assign n71543 = ~n71568;
  assign n70149 = n238 ^ n71417;
  assign n71422 = n71392 & n237;
  assign n71419 = ~n71392;
  assign n71435 = n71386 & n71407;
  assign n67514 = n71441 ^ n71442;
  assign n71436 = n71447 & n71448;
  assign n71433 = ~n71386;
  assign n71450 = n71458 & n71459;
  assign n71432 = ~n71462;
  assign n71465 = n71474 & n71475;
  assign n71421 = ~n71495;
  assign n71484 = n218 ^ n71506;
  assign n71455 = ~n71512;
  assign n71503 = n71516 & n7185;
  assign n71527 = n71533 & n71534;
  assign n71511 = n71543 & n71544;
  assign n71402 = ~n70149;
  assign n71414 = n71419 & n19432;
  assign n71377 = ~n71422;
  assign n71423 = n67514 & n70252;
  assign n71424 = n71433 & n71434;
  assign n71405 = ~n71435;
  assign n71415 = ~n71436;
  assign n67516 = ~n67514;
  assign n71431 = ~n71450;
  assign n71443 = ~n71465;
  assign n71358 = n71483 ^ n71484;
  assign n71425 = n71484 & n71488;
  assign n71482 = ~n71503;
  assign n71486 = n216 ^ n71511;
  assign n71504 = ~n71527;
  assign n71361 = n71402 & n71403;
  assign n71399 = ~n71414;
  assign n71391 = n71415 & n71416;
  assign n71412 = n67516 & n68814;
  assign n71400 = ~n71423;
  assign n71384 = ~n71424;
  assign n71406 = n71431 & n71432;
  assign n71418 = n71443 & n71444;
  assign n71453 = n71358 & n68740;
  assign n71460 = ~n71358;
  assign n71430 = ~n71425;
  assign n71428 = n71486 ^ n71487;
  assign n71479 = n71504 & n71505;
  assign n71369 = ~n71361;
  assign n71381 = n71391 ^ n71392;
  assign n71387 = n71406 ^ n71407;
  assign n71401 = ~n71412;
  assign n71398 = ~n71391;
  assign n71396 = n71418 ^ n68748;
  assign n71404 = ~n71406;
  assign n71420 = ~n71418;
  assign n71366 = ~n71453;
  assign n71449 = n71460 & n68706;
  assign n71456 = n217 ^ n71479;
  assign n71481 = ~n71479;
  assign n71362 = n237 ^ n71381;
  assign n71355 = n71386 ^ n71387;
  assign n67459 = n71395 ^ n71396;
  assign n71389 = n71398 & n71399;
  assign n71347 = n71400 & n71401;
  assign n71390 = n71404 & n71405;
  assign n71413 = n71420 & n71421;
  assign n71380 = ~n71449;
  assign n71426 = n71456 ^ n71457;
  assign n71471 = n71481 & n71482;
  assign n71345 = n71361 ^ n71362;
  assign n71324 = n71362 & n71369;
  assign n71350 = ~n71355;
  assign n71375 = n67459 & n70144;
  assign n71352 = ~n71347;
  assign n71376 = ~n71389;
  assign n67486 = ~n67459;
  assign n71383 = ~n71390;
  assign n71393 = ~n71413;
  assign n71320 = n71425 ^ n71426;
  assign n71429 = ~n71426;
  assign n71454 = ~n71471;
  assign n67220 = n71345 ^ n68287;
  assign n71241 = n71345 & n68277;
  assign n71344 = ~n71345;
  assign n71328 = ~n71324;
  assign n71357 = ~n71375;
  assign n71373 = n67486 & n68748;
  assign n71354 = n71376 & n71377;
  assign n71367 = n71383 & n71384;
  assign n71378 = n71393 & n71394;
  assign n71410 = n71320 & n68695;
  assign n71411 = ~n71320;
  assign n71408 = n71429 & n71430;
  assign n71427 = n71454 & n71455;
  assign n71317 = n67220 & n69344;
  assign n67222 = ~n67220;
  assign n71329 = n71344 & n68277;
  assign n71335 = n71354 ^ n71355;
  assign n71363 = n71354 & n19414;
  assign n71348 = n71367 ^ n71368;
  assign n71356 = ~n71373;
  assign n71370 = n71367 & n71368;
  assign n71360 = ~n71354;
  assign n71371 = ~n71367;
  assign n71359 = n71378 ^ n68706;
  assign n71379 = ~n71378;
  assign n71323 = ~n71410;
  assign n71397 = n71411 & n68661;
  assign n71409 = n71427 ^ n71428;
  assign n71310 = ~n71317;
  assign n71311 = ~n71329;
  assign n71325 = n236 ^ n71335;
  assign n71309 = n71347 ^ n71348;
  assign n71296 = n71356 & n71357;
  assign n67429 = n71358 ^ n71359;
  assign n71353 = n71360 & n236;
  assign n71349 = ~n71363;
  assign n71351 = ~n71370;
  assign n71364 = n71371 & n71372;
  assign n71374 = n71379 & n71380;
  assign n71340 = ~n71397;
  assign n71277 = n71408 ^ n71409;
  assign n71287 = n71310 & n71311;
  assign n71305 = n71324 ^ n71325;
  assign n71260 = n71325 & n71328;
  assign n71295 = ~n71309;
  assign n71336 = n71349 & n71350;
  assign n71338 = n67429 & n68740;
  assign n71341 = n71296 & n71316;
  assign n71342 = ~n71296;
  assign n71346 = n71351 & n71352;
  assign n67438 = ~n67429;
  assign n71327 = ~n71353;
  assign n71333 = ~n71364;
  assign n71365 = ~n71374;
  assign n71385 = n71277 & n68621;
  assign n71388 = ~n71277;
  assign n71265 = n71287 ^ n71288;
  assign n71283 = ~n71287;
  assign n71299 = n71305 & n68262;
  assign n71304 = ~n71305;
  assign n71274 = ~n71260;
  assign n71326 = ~n71336;
  assign n71319 = ~n71338;
  assign n71331 = n67438 & n70058;
  assign n71314 = ~n71341;
  assign n71330 = n71342 & n71343;
  assign n71332 = ~n71346;
  assign n71337 = n71365 & n71366;
  assign n71281 = ~n71385;
  assign n71382 = n71388 & n68658;
  assign n69068 = n263 ^ n71265;
  assign n70990 = n71265 & n263;
  assign n71102 = n71283 & n71284;
  assign n71282 = ~n71299;
  assign n71289 = n71304 & n68251;
  assign n71308 = n71326 & n71327;
  assign n71291 = ~n71330;
  assign n71318 = ~n71331;
  assign n71315 = n71332 & n71333;
  assign n71321 = n71337 ^ n68661;
  assign n71339 = ~n71337;
  assign n71301 = ~n71382;
  assign n70769 = ~n69068;
  assign n71279 = n71282 & n71241;
  assign n71264 = ~n71289;
  assign n71286 = n71308 ^ n71309;
  assign n71306 = n71308 & n19360;
  assign n71297 = n71315 ^ n71316;
  assign n71245 = n71318 & n71319;
  assign n67382 = n71320 ^ n71321;
  assign n71312 = ~n71308;
  assign n71313 = ~n71315;
  assign n71334 = n71339 & n71340;
  assign n71263 = ~n71279;
  assign n71273 = n71282 & n71264;
  assign n71261 = n71286 ^ n19360;
  assign n71249 = n71296 ^ n71297;
  assign n71294 = ~n71306;
  assign n71303 = n67382 & n68695;
  assign n71298 = n71312 & n235;
  assign n71252 = ~n71245;
  assign n71307 = n71313 & n71314;
  assign n67418 = ~n67382;
  assign n71322 = ~n71334;
  assign n71223 = n71260 ^ n71261;
  assign n71238 = n71263 & n71264;
  assign n71242 = ~n71273;
  assign n71191 = n71261 & n71274;
  assign n71226 = ~n71249;
  assign n71285 = n71294 & n71295;
  assign n71267 = ~n71298;
  assign n71293 = n67418 & n70020;
  assign n71275 = ~n71303;
  assign n71290 = ~n71307;
  assign n71302 = n71322 & n71323;
  assign n71222 = n71238 ^ n71223;
  assign n67099 = n71241 ^ n71242;
  assign n71234 = n71238 & n68068;
  assign n71236 = ~n71238;
  assign n71202 = ~n71191;
  assign n71266 = ~n71285;
  assign n71268 = n71290 & n71291;
  assign n71276 = ~n71293;
  assign n71278 = n71302 ^ n68621;
  assign n71300 = ~n71302;
  assign n71215 = n71222 & n68083;
  assign n71216 = n67099 & n69260;
  assign n71201 = ~n71222;
  assign n71224 = ~n71234;
  assign n67080 = ~n67099;
  assign n71232 = n71236 & n68083;
  assign n71248 = n71266 & n71267;
  assign n71246 = n71268 ^ n71269;
  assign n71181 = n71275 & n71276;
  assign n67351 = n71277 ^ n71278;
  assign n71272 = n71268 & n71269;
  assign n71270 = ~n71268;
  assign n71292 = n71300 & n71301;
  assign n67010 = n71201 ^ n68083;
  assign n71150 = ~n71215;
  assign n71210 = n67080 & n68251;
  assign n71197 = ~n71216;
  assign n71214 = n71223 & n71224;
  assign n71190 = ~n71232;
  assign n71180 = n71245 ^ n71246;
  assign n71218 = n71248 ^ n71249;
  assign n71244 = n71248 & n19316;
  assign n71254 = n71181 & n71259;
  assign n71250 = ~n71248;
  assign n71255 = n67351 & n69950;
  assign n67346 = ~n67351;
  assign n71257 = ~n71181;
  assign n71258 = n71270 & n71271;
  assign n71251 = ~n71272;
  assign n71280 = ~n71292;
  assign n67000 = ~n67010;
  assign n71198 = ~n71210;
  assign n71189 = ~n71214;
  assign n71192 = n234 ^ n71218;
  assign n71219 = n71180 & n19279;
  assign n71221 = ~n71180;
  assign n71225 = ~n71244;
  assign n71235 = n71250 & n234;
  assign n71243 = n71251 & n71252;
  assign n71239 = n67346 & n68621;
  assign n71206 = ~n71254;
  assign n71231 = ~n71255;
  assign n71240 = n71257 & n71200;
  assign n71228 = ~n71258;
  assign n71262 = n71280 & n71281;
  assign n71167 = n67000 & n69218;
  assign n71188 = n71189 & n71190;
  assign n71133 = n71191 ^ n71192;
  assign n71174 = n71197 & n71198;
  assign n71122 = n71192 & n71202;
  assign n71184 = ~n71219;
  assign n71213 = n71221 & n233;
  assign n71217 = n71225 & n71226;
  assign n71208 = ~n71235;
  assign n71230 = ~n71239;
  assign n71177 = ~n71240;
  assign n71227 = ~n71243;
  assign n71256 = n71262 & n68622;
  assign n71253 = ~n71262;
  assign n71149 = ~n71167;
  assign n71168 = n71174 & n71175;
  assign n71173 = n71133 & n67991;
  assign n71171 = ~n71174;
  assign n71169 = ~n71133;
  assign n71153 = ~n71188;
  assign n71155 = ~n71213;
  assign n71207 = ~n71217;
  assign n71199 = n71227 & n71228;
  assign n71157 = n71230 & n71231;
  assign n71247 = n71253 & n68565;
  assign n71233 = ~n71256;
  assign n71061 = n71149 & n71150;
  assign n71134 = n71153 ^ n68013;
  assign n71145 = ~n71168;
  assign n71162 = n71169 & n68013;
  assign n71163 = n71171 & n71172;
  assign n71152 = ~n71173;
  assign n71182 = n71199 ^ n71200;
  assign n71179 = n71207 & n71208;
  assign n71209 = n71157 & n71127;
  assign n71203 = ~n71157;
  assign n71205 = ~n71199;
  assign n71229 = n71233 & n71237;
  assign n71212 = ~n71247;
  assign n71116 = n71061 & n71089;
  assign n66925 = n71133 ^ n71134;
  assign n71117 = ~n71061;
  assign n71144 = n71152 & n71153;
  assign n71142 = n71145 & n71102;
  assign n71125 = ~n71162;
  assign n71120 = ~n71163;
  assign n71151 = n71179 ^ n71180;
  assign n71115 = n71181 ^ n71182;
  assign n71183 = ~n71179;
  assign n71193 = n71203 & n71204;
  assign n71194 = n71205 & n71206;
  assign n71148 = ~n71209;
  assign n71211 = ~n71229;
  assign n71220 = n71212 & n71233;
  assign n71101 = n66925 & n69170;
  assign n71086 = ~n71116;
  assign n71111 = n71117 & n71118;
  assign n66901 = ~n66925;
  assign n71119 = ~n71142;
  assign n71124 = ~n71144;
  assign n71137 = n71120 & n71145;
  assign n71123 = n233 ^ n71151;
  assign n71146 = n71115 & n232;
  assign n71158 = ~n71115;
  assign n71166 = n71183 & n71184;
  assign n71131 = ~n71193;
  assign n71176 = ~n71194;
  assign n71187 = n71211 & n71212;
  assign n71195 = ~n71220;
  assign n71070 = ~n71101;
  assign n71092 = n66901 & n68013;
  assign n71060 = ~n71111;
  assign n71088 = n71119 & n71120;
  assign n71048 = n71122 ^ n71123;
  assign n71110 = n71124 & n71125;
  assign n71103 = ~n71137;
  assign n71052 = n71123 & n71122;
  assign n71094 = ~n71146;
  assign n71141 = n71158 & n19255;
  assign n71154 = ~n71166;
  assign n71156 = n71176 & n71177;
  assign n71161 = n71187 ^ n68543;
  assign n67271 = n71195 ^ n71196;
  assign n71185 = ~n71187;
  assign n71062 = n71088 ^ n71089;
  assign n71069 = ~n71092;
  assign n71090 = n71048 & n67930;
  assign n71082 = n71102 ^ n71103;
  assign n71056 = ~n71110;
  assign n71087 = ~n71088;
  assign n71095 = ~n71048;
  assign n71071 = ~n71052;
  assign n71129 = ~n71141;
  assign n71114 = n71154 & n71155;
  assign n71126 = n71156 ^ n71157;
  assign n67249 = n71160 ^ n71161;
  assign n71147 = ~n71156;
  assign n71170 = n67271 & n68565;
  assign n71178 = n71185 & n71186;
  assign n67348 = ~n67271;
  assign n70976 = n71061 ^ n71062;
  assign n70987 = n71069 & n71070;
  assign n71047 = n71056 ^ n67930;
  assign n71073 = n71082 & n11627;
  assign n71072 = ~n71082;
  assign n71080 = n71086 & n71087;
  assign n71025 = ~n71090;
  assign n71081 = n71095 & n67937;
  assign n71096 = n71114 ^ n71115;
  assign n71022 = n71126 ^ n71127;
  assign n71128 = ~n71114;
  assign n71138 = n67249 & n68574;
  assign n71143 = n71147 & n71148;
  assign n67305 = ~n67249;
  assign n71159 = n67348 & n69893;
  assign n71139 = ~n71170;
  assign n71164 = ~n71178;
  assign n71031 = n70976 & n11492;
  assign n66796 = n71047 ^ n71048;
  assign n71038 = n70987 & n71049;
  assign n71028 = ~n70976;
  assign n71033 = ~n70987;
  assign n71054 = n71072 & n262;
  assign n71037 = ~n71073;
  assign n71059 = ~n71080;
  assign n71055 = ~n71081;
  assign n71053 = n232 ^ n71096;
  assign n71085 = n71022 & n19197;
  assign n71084 = ~n71022;
  assign n71112 = n71128 & n71129;
  assign n71113 = n67305 & n69839;
  assign n71106 = ~n71138;
  assign n71130 = ~n71143;
  assign n71140 = ~n71159;
  assign n71132 = n71164 & n71165;
  assign n71016 = n66796 & n67930;
  assign n71011 = n71028 & n261;
  assign n70969 = ~n71031;
  assign n71023 = n71033 & n71030;
  assign n66852 = ~n66796;
  assign n71013 = ~n71038;
  assign n71034 = n71037 & n70990;
  assign n70950 = n71052 ^ n71053;
  assign n71015 = ~n71054;
  assign n71046 = n71055 & n71056;
  assign n71029 = n71059 & n71060;
  assign n70992 = n71053 & n71071;
  assign n71079 = n71084 & n247;
  assign n71058 = ~n71085;
  assign n71093 = ~n71112;
  assign n71107 = ~n71113;
  assign n71099 = n71130 & n71131;
  assign n71105 = n71132 ^ n68496;
  assign n71063 = n71139 & n71140;
  assign n71135 = ~n71132;
  assign n70939 = ~n71011;
  assign n71001 = n66852 & n69115;
  assign n70978 = ~n71016;
  assign n70974 = ~n71023;
  assign n70988 = n71029 ^ n71030;
  assign n71014 = ~n71034;
  assign n71020 = n71037 & n71015;
  assign n71012 = ~n71029;
  assign n71024 = ~n71046;
  assign n71003 = ~n70992;
  assign n71027 = ~n71079;
  assign n71065 = n71093 & n71094;
  assign n71064 = n71099 ^ n71100;
  assign n71091 = n71099 & n71100;
  assign n67200 = n71104 ^ n71105;
  assign n70964 = n71106 & n71107;
  assign n71097 = ~n71099;
  assign n71121 = n71135 & n71136;
  assign n71075 = ~n71063;
  assign n70900 = n70987 ^ n70988;
  assign n70977 = ~n71001;
  assign n71000 = n71012 & n71013;
  assign n70975 = n71014 & n71015;
  assign n70991 = ~n71020;
  assign n70985 = n71024 & n71025;
  assign n70995 = n71063 ^ n71064;
  assign n71021 = n247 ^ n71065;
  assign n71057 = ~n71065;
  assign n71078 = n67200 & n68504;
  assign n70968 = ~n70964;
  assign n67264 = ~n67200;
  assign n71074 = ~n71091;
  assign n71083 = n71097 & n71098;
  assign n71108 = ~n71121;
  assign n70949 = n70900 & n260;
  assign n70948 = ~n70900;
  assign n70942 = n70975 ^ n70976;
  assign n70902 = n70977 & n70978;
  assign n70951 = n70985 ^ n67852;
  assign n69027 = n70990 ^ n70991;
  assign n70984 = n70985 & n67876;
  assign n70973 = ~n71000;
  assign n70970 = ~n70975;
  assign n70989 = ~n70985;
  assign n70993 = n71021 ^ n71022;
  assign n71019 = n70995 & n19179;
  assign n71032 = ~n70995;
  assign n71045 = n71057 & n71058;
  assign n71051 = n67264 & n69793;
  assign n71050 = n71074 & n71075;
  assign n71040 = ~n71078;
  assign n71036 = ~n71083;
  assign n71076 = n71108 & n71109;
  assign n68992 = n261 ^ n70942;
  assign n70936 = n70948 & n11437;
  assign n70871 = ~n70949;
  assign n66731 = n70950 ^ n70951;
  assign n70944 = n70902 & n70953;
  assign n70937 = ~n70902;
  assign n70966 = n70969 & n70970;
  assign n70933 = n70973 & n70974;
  assign n70683 = ~n69027;
  assign n70960 = ~n70984;
  assign n70979 = n70989 & n67852;
  assign n70855 = n70992 ^ n70993;
  assign n70912 = n70993 & n71003;
  assign n70982 = ~n71019;
  assign n71017 = n71032 & n246;
  assign n71026 = ~n71045;
  assign n71035 = ~n71050;
  assign n71039 = ~n71051;
  assign n71041 = n71076 ^ n71077;
  assign n71067 = ~n71076;
  assign n70914 = n66731 & n69077;
  assign n70598 = ~n68992;
  assign n70903 = n70933 ^ n70934;
  assign n66762 = ~n66731;
  assign n70905 = ~n70936;
  assign n70930 = n70937 & n70934;
  assign n70916 = ~n70944;
  assign n70952 = n70960 & n70950;
  assign n70915 = ~n70933;
  assign n70954 = n70855 & n67796;
  assign n70938 = ~n70966;
  assign n70928 = ~n70979;
  assign n70947 = ~n70855;
  assign n70921 = ~n70912;
  assign n70957 = ~n71017;
  assign n70994 = n71026 & n71027;
  assign n71008 = n71035 & n71036;
  assign n70875 = n71039 & n71040;
  assign n67145 = n68450 ^ n71041;
  assign n71044 = n71041 & n68450;
  assign n71066 = n71067 & n71068;
  assign n70838 = n70902 ^ n70903;
  assign n70884 = ~n70914;
  assign n70904 = n70915 & n70916;
  assign n70901 = n66762 & n67852;
  assign n70883 = ~n70930;
  assign n70899 = n70938 & n70939;
  assign n70935 = n70947 & n67782;
  assign n70927 = ~n70952;
  assign n70892 = ~n70954;
  assign n70955 = n70994 ^ n70995;
  assign n70965 = n71008 ^ n70999;
  assign n70981 = ~n70994;
  assign n71009 = n70875 & n70908;
  assign n71002 = n71008 & n71018;
  assign n70997 = n67145 & n69745;
  assign n71004 = ~n70875;
  assign n67204 = ~n67145;
  assign n70998 = ~n71008;
  assign n70972 = ~n71044;
  assign n71042 = ~n71066;
  assign n70872 = n70838 & n259;
  assign n70868 = ~n70838;
  assign n70869 = n70899 ^ n70900;
  assign n70885 = ~n70901;
  assign n70882 = ~n70904;
  assign n70906 = ~n70899;
  assign n70886 = n70927 & n70928;
  assign n70862 = ~n70935;
  assign n70913 = n246 ^ n70955;
  assign n70919 = n70964 ^ n70965;
  assign n70980 = n70981 & n70982;
  assign n70971 = ~n70997;
  assign n70986 = n70998 & n70999;
  assign n70967 = ~n71002;
  assign n70996 = n71004 & n71005;
  assign n70910 = ~n71009;
  assign n71010 = n71042 & n71043;
  assign n70860 = n70868 & n11347;
  assign n68929 = n260 ^ n70869;
  assign n70799 = ~n70872;
  assign n70844 = n70882 & n70883;
  assign n70813 = n70884 & n70885;
  assign n70856 = n70886 ^ n67782;
  assign n70890 = n70905 & n70906;
  assign n70891 = ~n70886;
  assign n70784 = n70912 ^ n70913;
  assign n70920 = ~n70913;
  assign n70929 = n70919 & n245;
  assign n70932 = ~n70919;
  assign n70961 = n70967 & n70968;
  assign n70803 = n70971 & n70972;
  assign n70956 = ~n70980;
  assign n70946 = ~n70986;
  assign n70874 = ~n70996;
  assign n70959 = n71010 ^ n68405;
  assign n71006 = ~n71010;
  assign n70814 = n70844 ^ n70845;
  assign n70846 = n70813 & n70845;
  assign n66648 = n70855 ^ n70856;
  assign n70840 = ~n70860;
  assign n70819 = ~n70844;
  assign n70850 = ~n70813;
  assign n70870 = ~n70890;
  assign n70881 = n70891 & n70892;
  assign n70878 = n70784 & n67720;
  assign n70877 = ~n70784;
  assign n70847 = n70920 & n70921;
  assign n70864 = ~n70929;
  assign n70917 = n70932 & n19125;
  assign n70918 = n70956 & n70957;
  assign n70943 = n70803 & n70833;
  assign n70940 = ~n70803;
  assign n67089 = n70958 ^ n70959;
  assign n70945 = ~n70961;
  assign n70983 = n71006 & n71007;
  assign n70768 = n70813 ^ n70814;
  assign n70827 = n66648 & n67782;
  assign n66688 = ~n66648;
  assign n70820 = ~n70846;
  assign n70836 = n70850 & n70851;
  assign n70837 = n70870 & n70871;
  assign n70867 = n70877 & n67747;
  assign n70830 = ~n70878;
  assign n70861 = ~n70881;
  assign n70887 = ~n70917;
  assign n70879 = n70918 ^ n70919;
  assign n70931 = n67089 & n68411;
  assign n70888 = ~n70918;
  assign n70924 = n70940 & n70941;
  assign n70835 = ~n70943;
  assign n70907 = n70945 & n70946;
  assign n67163 = ~n67089;
  assign n70962 = ~n70983;
  assign n70772 = n70768 & n11226;
  assign n70776 = ~n70768;
  assign n70810 = n70819 & n70820;
  assign n70806 = n66688 & n69048;
  assign n70783 = ~n70827;
  assign n70794 = ~n70836;
  assign n70795 = n70837 ^ n70838;
  assign n70818 = n70861 & n70862;
  assign n70841 = ~n70837;
  assign n70787 = ~n70867;
  assign n70848 = n245 ^ n70879;
  assign n70880 = n70887 & n70888;
  assign n70876 = n70907 ^ n70908;
  assign n70909 = ~n70907;
  assign n70802 = ~n70924;
  assign n70895 = ~n70931;
  assign n70922 = n67163 & n69707;
  assign n70923 = n70962 & n70963;
  assign n70738 = ~n70772;
  assign n70762 = n70776 & n258;
  assign n70761 = n259 ^ n70795;
  assign n70782 = ~n70806;
  assign n70793 = ~n70810;
  assign n70785 = n70818 ^ n67720;
  assign n70815 = n70840 & n70841;
  assign n70698 = n70847 ^ n70848;
  assign n70831 = ~n70818;
  assign n70746 = n70848 & n70847;
  assign n70817 = n70875 ^ n70876;
  assign n70863 = ~n70880;
  assign n70889 = n70909 & n70910;
  assign n70896 = ~n70922;
  assign n70894 = n70923 ^ n68354;
  assign n70925 = ~n70923;
  assign n68897 = n70761 ^ n68929;
  assign n70704 = ~n70762;
  assign n70685 = n70761 & n68929;
  assign n70710 = n70782 & n70783;
  assign n66559 = n70784 ^ n70785;
  assign n70744 = n70793 & n70794;
  assign n70798 = ~n70815;
  assign n70809 = n70698 & n67688;
  assign n70808 = n70830 & n70831;
  assign n70807 = ~n70698;
  assign n70757 = ~n70746;
  assign n70842 = n70817 & n19082;
  assign n70816 = n70863 & n70864;
  assign n70839 = ~n70817;
  assign n70873 = ~n70889;
  assign n67026 = n70893 ^ n70894;
  assign n70718 = n70895 & n70896;
  assign n70911 = n70925 & n70926;
  assign n70422 = ~n68897;
  assign n70711 = n70744 ^ n70745;
  assign n70739 = n66559 & n69008;
  assign n70690 = ~n70685;
  assign n70751 = n70710 & n70745;
  assign n70756 = n66559 & n70769;
  assign n70742 = ~n70710;
  assign n70721 = ~n70744;
  assign n66594 = ~n66559;
  assign n70767 = n70798 & n70799;
  assign n70797 = n70807 & n67678;
  assign n70786 = ~n70808;
  assign n70749 = ~n70809;
  assign n70789 = n70816 ^ n70817;
  assign n70821 = n70839 & n244;
  assign n70811 = ~n70842;
  assign n70812 = ~n70816;
  assign n70866 = n67026 & n69653;
  assign n70832 = n70873 & n70874;
  assign n70857 = n70718 & n70760;
  assign n70858 = ~n70718;
  assign n67109 = ~n67026;
  assign n70897 = ~n70911;
  assign n70669 = n70710 ^ n70711;
  assign n70700 = ~n70739;
  assign n70732 = n70742 & n70743;
  assign n70728 = n66594 & n67747;
  assign n70720 = ~n70751;
  assign n70727 = n66594 & n69068;
  assign n69084 = ~n70756;
  assign n70717 = n70767 ^ n70768;
  assign n70737 = ~n70767;
  assign n70754 = n70786 & n70787;
  assign n70747 = n244 ^ n70789;
  assign n70713 = ~n70797;
  assign n70796 = n70811 & n70812;
  assign n70771 = ~n70821;
  assign n70804 = n70832 ^ n70833;
  assign n70849 = n67109 & n68354;
  assign n70765 = ~n70857;
  assign n70843 = n70858 & n70859;
  assign n70834 = ~n70832;
  assign n70823 = ~n70866;
  assign n70865 = n70897 & n70898;
  assign n70661 = n70669 & n11154;
  assign n70666 = ~n70669;
  assign n70686 = n258 ^ n70717;
  assign n70697 = n70720 & n70721;
  assign n69064 = ~n70727;
  assign n70701 = ~n70728;
  assign n70676 = ~n70732;
  assign n70724 = n70737 & n70738;
  assign n70629 = n70746 ^ n70747;
  assign n70699 = n70754 ^ n67678;
  assign n70646 = n70747 & n70757;
  assign n70750 = ~n70754;
  assign n70770 = ~n70796;
  assign n70726 = n70803 ^ n70804;
  assign n70822 = n70834 & n70835;
  assign n70723 = ~n70843;
  assign n70824 = ~n70849;
  assign n70829 = n70865 ^ n68315;
  assign n70853 = ~n70865;
  assign n70632 = ~n70661;
  assign n70642 = n70666 & n257;
  assign n68865 = n70685 ^ n70686;
  assign n70583 = n70686 & n70690;
  assign n70675 = ~n70697;
  assign n66492 = n70698 ^ n70699;
  assign n70601 = n70700 & n70701;
  assign n70702 = n70629 & n67628;
  assign n70703 = ~n70724;
  assign n70694 = ~n70629;
  assign n70731 = n70749 & n70750;
  assign n70725 = n70770 & n70771;
  assign n70758 = n70726 & n19042;
  assign n70763 = ~n70726;
  assign n70801 = ~n70822;
  assign n70635 = n70823 & n70824;
  assign n66948 = n70828 ^ n70829;
  assign n70852 = n70853 & n70854;
  assign n70597 = ~n70642;
  assign n70349 = ~n68865;
  assign n70671 = n66492 & n67678;
  assign n70633 = n70675 & n70676;
  assign n70670 = n66492 & n70683;
  assign n70582 = ~n70583;
  assign n70672 = n70601 & n70684;
  assign n70667 = ~n70601;
  assign n66521 = ~n66492;
  assign n70693 = n70694 & n67640;
  assign n70664 = ~n70702;
  assign n70668 = n70703 & n70704;
  assign n70689 = n70725 ^ n70726;
  assign n70712 = ~n70731;
  assign n70730 = ~n70725;
  assign n70729 = ~n70758;
  assign n70748 = n70763 & n243;
  assign n70781 = n70635 & n70800;
  assign n70759 = n70801 & n70802;
  assign n70780 = n66948 & n70805;
  assign n70792 = n66948 & n68315;
  assign n67053 = ~n66948;
  assign n70788 = ~n70635;
  assign n70825 = ~n70852;
  assign n70602 = n70633 ^ n70634;
  assign n70645 = n66521 & n69027;
  assign n70650 = n66521 & n68972;
  assign n70649 = n70667 & n70634;
  assign n70628 = n70668 ^ n70669;
  assign n69030 = ~n70670;
  assign n70622 = ~n70671;
  assign n70641 = ~n70633;
  assign n70640 = ~n70672;
  assign n70631 = ~n70668;
  assign n70647 = n243 ^ n70689;
  assign n70617 = ~n70693;
  assign n70658 = n70712 & n70713;
  assign n70716 = n70729 & n70730;
  assign n70688 = ~n70748;
  assign n70719 = n70759 ^ n70760;
  assign n69674 = ~n70780;
  assign n70679 = ~n70781;
  assign n70773 = n67053 & n69614;
  assign n70775 = n67053 & n69676;
  assign n70774 = n70788 & n70682;
  assign n70764 = ~n70759;
  assign n70753 = ~n70792;
  assign n70791 = n70825 & n70826;
  assign n70562 = n70601 ^ n70602;
  assign n70584 = n257 ^ n70628;
  assign n70619 = n70631 & n70632;
  assign n70618 = n70640 & n70641;
  assign n69052 = ~n70645;
  assign n70538 = n70646 ^ n70647;
  assign n70606 = ~n70649;
  assign n70621 = ~n70650;
  assign n70630 = n70658 ^ n67628;
  assign n70571 = n70647 & n70646;
  assign n70663 = ~n70658;
  assign n70687 = ~n70716;
  assign n70653 = n70718 ^ n70719;
  assign n70755 = n70764 & n70765;
  assign n70752 = ~n70773;
  assign n70639 = ~n70774;
  assign n69692 = ~n70775;
  assign n66838 = n70790 ^ n70791;
  assign n70778 = ~n70791;
  assign n70557 = n70562 & n256;
  assign n68830 = n70583 ^ n70584;
  assign n70560 = ~n70562;
  assign n70581 = ~n70584;
  assign n70605 = ~n70618;
  assign n70596 = ~n70619;
  assign n70527 = n70621 & n70622;
  assign n66420 = n70629 ^ n70630;
  assign n70614 = n70538 & n67591;
  assign n70609 = ~n70538;
  assign n70648 = n70663 & n70664;
  assign n70652 = n70687 & n70688;
  assign n70680 = n70653 & n19000;
  assign n70677 = ~n70653;
  assign n70558 = n70752 & n70753;
  assign n70722 = ~n70755;
  assign n70741 = n66838 & n69581;
  assign n70740 = n66838 & n70766;
  assign n66973 = ~n66838;
  assign n70777 = n70778 & n70779;
  assign n70477 = ~n70557;
  assign n70548 = n70560 & n11085;
  assign n70217 = ~n68830;
  assign n70485 = n70581 & n70582;
  assign n70561 = n70596 & n70597;
  assign n70586 = n66420 & n70598;
  assign n70587 = n66420 & n68920;
  assign n70579 = n70527 & n70603;
  assign n70553 = n70605 & n70606;
  assign n70585 = ~n70527;
  assign n70595 = n70609 & n67595;
  assign n66440 = ~n66420;
  assign n70532 = ~n70614;
  assign n70616 = ~n70648;
  assign n70611 = n70652 ^ n70653;
  assign n70644 = ~n70652;
  assign n70662 = n70677 & n242;
  assign n70643 = ~n70680;
  assign n70707 = n70558 & n70594;
  assign n70681 = n70722 & n70723;
  assign n70695 = ~n70558;
  assign n70734 = n66973 & n69631;
  assign n69655 = ~n70740;
  assign n70705 = ~n70741;
  assign n70733 = n66973 & n68212;
  assign n70735 = ~n70777;
  assign n70522 = ~n70548;
  assign n70528 = n70553 ^ n70554;
  assign n70524 = n70561 ^ n70562;
  assign n70523 = ~n70561;
  assign n70552 = ~n70553;
  assign n70551 = ~n70579;
  assign n70570 = n70585 & n70554;
  assign n69013 = ~n70586;
  assign n70567 = n66440 & n68992;
  assign n70546 = ~n70587;
  assign n70566 = n66440 & n67640;
  assign n70569 = ~n70595;
  assign n70572 = n242 ^ n70611;
  assign n70615 = n70616 & n70617;
  assign n70637 = n70643 & n70644;
  assign n70608 = ~n70662;
  assign n70636 = n70681 ^ n70682;
  assign n70691 = n70695 & n70696;
  assign n70678 = ~n70681;
  assign n70600 = ~n70707;
  assign n70706 = ~n70733;
  assign n69634 = ~n70734;
  assign n70708 = n70735 & n70736;
  assign n70504 = n70522 & n70523;
  assign n70486 = n256 ^ n70524;
  assign n70444 = n70527 ^ n70528;
  assign n70547 = n70551 & n70552;
  assign n70545 = ~n70566;
  assign n68989 = ~n70567;
  assign n70521 = ~n70570;
  assign n70457 = n70571 ^ n70572;
  assign n70497 = n70572 & n70571;
  assign n70568 = ~n70615;
  assign n70574 = n70635 ^ n70636;
  assign n70607 = ~n70637;
  assign n70657 = n70678 & n70679;
  assign n70564 = ~n70691;
  assign n70516 = n70705 & n70706;
  assign n70659 = n70708 ^ n70709;
  assign n70714 = ~n70708;
  assign n68796 = n70485 ^ n70486;
  assign n70362 = n70486 & n70485;
  assign n70494 = n70444 & n271;
  assign n70476 = ~n70504;
  assign n70482 = ~n70444;
  assign n70450 = n70545 & n70546;
  assign n70520 = ~n70547;
  assign n70539 = n70457 & n67545;
  assign n70533 = ~n70457;
  assign n70512 = ~n70497;
  assign n70565 = n70568 & n70569;
  assign n70537 = n70568 ^ n67591;
  assign n70592 = n70574 & n241;
  assign n70573 = n70607 & n70608;
  assign n70604 = ~n70574;
  assign n70638 = ~n70657;
  assign n66766 = n68191 ^ n70659;
  assign n70665 = n70516 & n70479;
  assign n70655 = ~n70516;
  assign n70660 = ~n70659;
  assign n70692 = n70714 & n70715;
  assign n70165 = ~n68796;
  assign n70443 = n70476 & n70477;
  assign n70472 = n70482 & n10976;
  assign n70367 = ~n70362;
  assign n70395 = ~n70494;
  assign n70502 = n70450 & n70491;
  assign n70490 = n70520 & n70521;
  assign n70526 = n70533 & n67568;
  assign n70513 = ~n70450;
  assign n66357 = n70537 ^ n70538;
  assign n70456 = ~n70539;
  assign n70531 = ~n70565;
  assign n70540 = n70573 ^ n70574;
  assign n70519 = ~n70592;
  assign n70580 = n70604 & n18956;
  assign n70555 = ~n70573;
  assign n70623 = n66766 & n69620;
  assign n70593 = n70638 & n70639;
  assign n66910 = ~n66766;
  assign n70654 = n70655 & n70656;
  assign n70651 = n70660 & n68191;
  assign n70530 = ~n70665;
  assign n70673 = ~n70692;
  assign n70393 = n70443 ^ n70444;
  assign n70438 = ~n70443;
  assign n70437 = ~n70472;
  assign n70451 = n70490 ^ n70491;
  assign n70487 = ~n70502;
  assign n70488 = ~n70490;
  assign n70501 = n66357 & n67591;
  assign n70495 = n70513 & n70514;
  assign n66382 = ~n66357;
  assign n70500 = ~n70526;
  assign n70496 = n70531 & n70532;
  assign n70498 = n241 ^ n70540;
  assign n70556 = ~n70580;
  assign n70559 = n70593 ^ n70594;
  assign n70612 = n66910 & n70620;
  assign n70613 = n66910 & n69517;
  assign n69598 = ~n70623;
  assign n70599 = ~n70593;
  assign n70590 = ~n70651;
  assign n70484 = ~n70654;
  assign n70626 = n70673 & n70674;
  assign n70363 = n271 ^ n70393;
  assign n70425 = n70437 & n70438;
  assign n70369 = n70450 ^ n70451;
  assign n70467 = n70487 & n70488;
  assign n70481 = n66382 & n68878;
  assign n70436 = ~n70495;
  assign n70458 = n70496 ^ n67545;
  assign n70376 = n70497 ^ n70498;
  assign n70453 = ~n70501;
  assign n70404 = n70498 & n70512;
  assign n70499 = ~n70496;
  assign n70544 = n70555 & n70556;
  assign n70475 = n70558 ^ n70559;
  assign n70588 = n70599 & n70600;
  assign n69625 = ~n70612;
  assign n70589 = ~n70613;
  assign n70591 = n70626 ^ n70627;
  assign n70624 = ~n70626;
  assign n68757 = n70362 ^ n70363;
  assign n70366 = ~n70363;
  assign n70412 = n70369 & n10896;
  assign n70394 = ~n70425;
  assign n70408 = ~n70369;
  assign n66320 = n70457 ^ n70458;
  assign n70435 = ~n70467;
  assign n70454 = ~n70481;
  assign n70421 = ~n70404;
  assign n70480 = n70499 & n70500;
  assign n70517 = n70475 & n18899;
  assign n70525 = ~n70475;
  assign n70518 = ~n70544;
  assign n70563 = ~n70588;
  assign n70400 = n70589 & n70590;
  assign n66681 = n68111 ^ n70591;
  assign n70578 = ~n70591;
  assign n70610 = n70624 & n70625;
  assign n70096 = ~n68757;
  assign n70278 = n70366 & n70367;
  assign n70368 = n70394 & n70395;
  assign n70387 = n70408 & n270;
  assign n70360 = ~n70412;
  assign n70417 = n66320 & n68897;
  assign n70416 = n66320 & n68845;
  assign n70406 = n70435 & n70436;
  assign n66308 = ~n66320;
  assign n70364 = n70453 & n70454;
  assign n70455 = ~n70480;
  assign n70493 = ~n70517;
  assign n70474 = n70518 & n70519;
  assign n70503 = n70525 & n240;
  assign n70549 = n66681 & n69559;
  assign n70515 = n70563 & n70564;
  assign n66823 = ~n66681;
  assign n70420 = ~n70400;
  assign n70575 = n70578 & n68111;
  assign n70576 = ~n70610;
  assign n70325 = n70368 ^ n70369;
  assign n70316 = ~n70387;
  assign n70361 = ~n70368;
  assign n70365 = n70406 ^ n70407;
  assign n70379 = ~n70416;
  assign n68928 = ~n70417;
  assign n70396 = n66308 & n67545;
  assign n70411 = n66308 & n70422;
  assign n70418 = n70364 & n70430;
  assign n70383 = ~n70406;
  assign n70423 = ~n70364;
  assign n70414 = n70455 & n70456;
  assign n70446 = n70474 ^ n70475;
  assign n70448 = ~n70503;
  assign n70492 = ~n70474;
  assign n70478 = n70515 ^ n70516;
  assign n70535 = n66823 & n69467;
  assign n69563 = ~n70549;
  assign n70536 = n66823 & n70550;
  assign n70529 = ~n70515;
  assign n70511 = ~n70575;
  assign n70541 = n70576 & n70577;
  assign n70279 = n270 ^ n70325;
  assign n70345 = n70360 & n70361;
  assign n70277 = n70364 ^ n70365;
  assign n70378 = ~n70396;
  assign n68909 = ~n70411;
  assign n70377 = n70414 ^ n67514;
  assign n70384 = ~n70418;
  assign n70397 = n70423 & n70407;
  assign n70415 = n70414 & n67514;
  assign n70424 = ~n70414;
  assign n70405 = n240 ^ n70446;
  assign n70410 = n70478 ^ n70479;
  assign n70469 = n70492 & n70493;
  assign n70505 = n70529 & n70530;
  assign n70510 = ~n70535;
  assign n69583 = ~n70536;
  assign n70507 = n70541 ^ n68036;
  assign n70542 = ~n70541;
  assign n68714 = n70278 ^ n70279;
  assign n70198 = n70279 & n70278;
  assign n70331 = n70277 & n269;
  assign n70326 = ~n70277;
  assign n70315 = ~n70345;
  assign n66225 = n70376 ^ n70377;
  assign n70266 = n70378 & n70379;
  assign n70372 = n70383 & n70384;
  assign n70342 = ~n70397;
  assign n70264 = n70404 ^ n70405;
  assign n70386 = ~n70415;
  assign n70317 = n70405 & n70421;
  assign n70398 = n70424 & n67516;
  assign n70439 = n70410 & n18888;
  assign n70442 = ~n70410;
  assign n70447 = ~n70469;
  assign n70483 = ~n70505;
  assign n66637 = n70506 ^ n70507;
  assign n70335 = n70510 & n70511;
  assign n70534 = n70542 & n70543;
  assign n70021 = ~n68714;
  assign n70276 = n70315 & n70316;
  assign n70308 = n70326 & n10806;
  assign n70242 = ~n70331;
  assign n70332 = n70266 & n70340;
  assign n70333 = n66225 & n67516;
  assign n70337 = n66225 & n70349;
  assign n70336 = ~n70266;
  assign n66271 = ~n66225;
  assign n70341 = ~n70372;
  assign n70370 = n70264 & n67459;
  assign n70380 = n70386 & n70376;
  assign n70359 = ~n70264;
  assign n70353 = ~n70398;
  assign n70322 = ~n70317;
  assign n70403 = ~n70439;
  assign n70432 = n70442 & n255;
  assign n70409 = n70447 & n70448;
  assign n70468 = n66637 & n69549;
  assign n70440 = n70483 & n70484;
  assign n70465 = n70335 & n70489;
  assign n70473 = n66637 & n69472;
  assign n70463 = ~n70335;
  assign n66743 = ~n66637;
  assign n70508 = ~n70534;
  assign n70240 = n70276 ^ n70277;
  assign n70284 = ~n70276;
  assign n70283 = ~n70308;
  assign n70307 = ~n70332;
  assign n70323 = n66271 & n68814;
  assign n70292 = ~n70333;
  assign n70330 = n66271 & n68865;
  assign n70324 = n70336 & n70313;
  assign n68873 = ~n70337;
  assign n70312 = n70341 & n70342;
  assign n70354 = n70359 & n67486;
  assign n70311 = ~n70370;
  assign n70352 = ~n70380;
  assign n70357 = n70409 ^ n70410;
  assign n70402 = ~n70409;
  assign n70356 = ~n70432;
  assign n70401 = n70440 ^ n70441;
  assign n70445 = n70440 & n70460;
  assign n70459 = n70463 & n70296;
  assign n70452 = n66743 & n70464;
  assign n70339 = ~n70465;
  assign n70461 = n66743 & n68038;
  assign n70449 = ~n70440;
  assign n69540 = ~n70468;
  assign n70433 = ~n70473;
  assign n70466 = n70508 & n70509;
  assign n70199 = n269 ^ n70240;
  assign n70260 = n70283 & n70284;
  assign n70267 = n70312 ^ n70313;
  assign n70293 = ~n70323;
  assign n70269 = ~n70324;
  assign n68885 = ~n70330;
  assign n70306 = ~n70312;
  assign n70299 = n70352 & n70353;
  assign n70259 = ~n70354;
  assign n70318 = n255 ^ n70357;
  assign n70320 = n70400 ^ n70401;
  assign n70388 = n70402 & n70403;
  assign n70419 = ~n70445;
  assign n70431 = n70449 & n70441;
  assign n69528 = ~n70452;
  assign n70286 = ~n70459;
  assign n70434 = ~n70461;
  assign n70429 = n70466 ^ n67963;
  assign n70470 = ~n70466;
  assign n68687 = n70198 ^ n70199;
  assign n70197 = ~n70199;
  assign n70241 = ~n70260;
  assign n70194 = n70266 ^ n70267;
  assign n70174 = n70292 & n70293;
  assign n70265 = n70299 ^ n67459;
  assign n70294 = n70306 & n70307;
  assign n70176 = n70317 ^ n70318;
  assign n70310 = ~n70299;
  assign n70321 = ~n70318;
  assign n70358 = n70320 & n254;
  assign n70371 = ~n70320;
  assign n70355 = ~n70388;
  assign n70413 = n70419 & n70420;
  assign n66564 = n70428 ^ n70429;
  assign n70375 = ~n70431;
  assign n70207 = n70433 & n70434;
  assign n70462 = n70470 & n70471;
  assign n69948 = ~n68687;
  assign n70124 = n70197 & n70198;
  assign n70193 = n70241 & n70242;
  assign n70220 = n70194 & n268;
  assign n70228 = ~n70194;
  assign n70253 = n70174 & n70216;
  assign n66193 = n70264 ^ n70265;
  assign n70251 = ~n70174;
  assign n70274 = n70176 & n67438;
  assign n70268 = ~n70294;
  assign n70289 = n70310 & n70311;
  assign n70280 = ~n70176;
  assign n70246 = n70321 & n70322;
  assign n70319 = n70355 & n70356;
  assign n70282 = ~n70358;
  assign n70346 = n70371 & n18839;
  assign n70385 = n66564 & n70399;
  assign n70392 = n66564 & n69381;
  assign n70374 = ~n70413;
  assign n66658 = ~n66564;
  assign n70225 = ~n70207;
  assign n70426 = ~n70462;
  assign n70130 = ~n70124;
  assign n70167 = n70193 ^ n70194;
  assign n70185 = ~n70193;
  assign n70160 = ~n70220;
  assign n70211 = n70228 & n10723;
  assign n70231 = n66193 & n68748;
  assign n70218 = n66193 & n68830;
  assign n66209 = ~n66193;
  assign n70237 = n70251 & n70252;
  assign n70233 = ~n70253;
  assign n70215 = n70268 & n70269;
  assign n70226 = ~n70274;
  assign n70263 = n70280 & n67429;
  assign n70258 = ~n70289;
  assign n70244 = ~n70246;
  assign n70275 = n70319 ^ n70320;
  assign n70327 = ~n70319;
  assign n70328 = ~n70346;
  assign n70334 = n70374 & n70375;
  assign n70382 = n66658 & n67963;
  assign n70381 = n66658 & n69479;
  assign n69499 = ~n70385;
  assign n70343 = ~n70392;
  assign n70389 = n70426 & n70427;
  assign n70125 = n268 ^ n70167;
  assign n70184 = ~n70211;
  assign n70175 = n70215 ^ n70216;
  assign n70203 = n66209 & n70217;
  assign n68847 = ~n70218;
  assign n70204 = n66209 & n67486;
  assign n70187 = ~n70231;
  assign n70192 = ~n70237;
  assign n70232 = ~n70215;
  assign n70221 = n70258 & n70259;
  assign n70189 = ~n70263;
  assign n70247 = n254 ^ n70275;
  assign n70300 = n70327 & n70328;
  assign n70295 = n70334 ^ n70335;
  assign n70338 = ~n70334;
  assign n69482 = ~n70381;
  assign n70344 = ~n70382;
  assign n70348 = n70389 ^ n67905;
  assign n70390 = ~n70389;
  assign n68630 = n70124 ^ n70125;
  assign n70046 = n70125 & n70130;
  assign n70121 = n70174 ^ n70175;
  assign n70171 = n70184 & n70185;
  assign n68833 = ~n70203;
  assign n70186 = ~n70204;
  assign n70177 = n70221 ^ n67429;
  assign n70210 = n70232 & n70233;
  assign n70109 = n70246 ^ n70247;
  assign n70227 = ~n70221;
  assign n70243 = ~n70247;
  assign n70236 = n70295 ^ n70296;
  assign n70281 = ~n70300;
  assign n70329 = n70338 & n70339;
  assign n70103 = n70343 & n70344;
  assign n66481 = n70347 ^ n70348;
  assign n70373 = n70390 & n70391;
  assign n69890 = ~n68630;
  assign n70153 = n70121 & n10627;
  assign n70159 = ~n70171;
  assign n70142 = ~n70121;
  assign n66152 = n70176 ^ n70177;
  assign n70116 = n70186 & n70187;
  assign n70200 = n70109 & n67382;
  assign n70191 = ~n70210;
  assign n70202 = n70226 & n70227;
  assign n70201 = ~n70109;
  assign n70163 = n70243 & n70244;
  assign n70250 = n70236 & n253;
  assign n70235 = n70281 & n70282;
  assign n70254 = ~n70236;
  assign n70305 = n70103 & n70158;
  assign n70314 = n66481 & n69459;
  assign n70301 = n66481 & n69336;
  assign n70285 = ~n70329;
  assign n66571 = ~n66481;
  assign n70297 = ~n70103;
  assign n70350 = ~n70373;
  assign n70138 = n70142 & n267;
  assign n70115 = ~n70153;
  assign n70120 = n70159 & n70160;
  assign n70156 = n66152 & n70165;
  assign n70161 = n70116 & n70166;
  assign n70145 = n66152 & n67429;
  assign n70152 = ~n70116;
  assign n66175 = ~n66152;
  assign n70143 = n70191 & n70192;
  assign n70102 = ~n70200;
  assign n70190 = n70201 & n67418;
  assign n70188 = ~n70202;
  assign n70170 = ~n70163;
  assign n70195 = n70235 ^ n70236;
  assign n70173 = ~n70250;
  assign n70245 = n70254 & n18788;
  assign n70206 = ~n70235;
  assign n70248 = n70285 & n70286;
  assign n70290 = n70297 & n70298;
  assign n70273 = ~n70301;
  assign n70287 = n66571 & n67899;
  assign n70151 = ~n70305;
  assign n70291 = n66571 & n70309;
  assign n69457 = ~n70314;
  assign n70304 = n70350 & n70351;
  assign n70087 = n70120 ^ n70121;
  assign n70114 = ~n70120;
  assign n70086 = ~n70138;
  assign n70117 = n70143 ^ n70144;
  assign n70113 = ~n70145;
  assign n70135 = n66175 & n68740;
  assign n70141 = n70152 & n70144;
  assign n70136 = n66175 & n68796;
  assign n68799 = ~n70156;
  assign n70126 = ~n70161;
  assign n70127 = ~n70143;
  assign n70146 = n70188 & n70189;
  assign n70155 = ~n70190;
  assign n70164 = n253 ^ n70195;
  assign n70205 = ~n70245;
  assign n70208 = n70248 ^ n70249;
  assign n70255 = n70248 & n70249;
  assign n70256 = ~n70248;
  assign n70272 = ~n70287;
  assign n70108 = ~n70290;
  assign n69442 = ~n70291;
  assign n70271 = n70304 ^ n67826;
  assign n70302 = ~n70304;
  assign n70047 = n267 ^ n70087;
  assign n70099 = n70114 & n70115;
  assign n70043 = n70116 ^ n70117;
  assign n70111 = n70126 & n70127;
  assign n70112 = ~n70135;
  assign n68818 = ~n70136;
  assign n70095 = ~n70141;
  assign n70110 = n70146 ^ n67382;
  assign n70051 = n70163 ^ n70164;
  assign n70154 = ~n70146;
  assign n70063 = n70164 & n70170;
  assign n70196 = n70205 & n70206;
  assign n70132 = n70207 ^ n70208;
  assign n70224 = ~n70255;
  assign n70238 = n70256 & n70257;
  assign n66410 = n70270 ^ n70271;
  assign n70040 = n70272 & n70273;
  assign n70288 = n70302 & n70303;
  assign n68586 = n70046 ^ n70047;
  assign n70050 = ~n70047;
  assign n70074 = n70043 & n266;
  assign n70085 = ~n70099;
  assign n70073 = ~n70043;
  assign n66096 = n70109 ^ n70110;
  assign n70094 = ~n70111;
  assign n70027 = n70112 & n70113;
  assign n70123 = n70051 & n67346;
  assign n70137 = n70154 & n70155;
  assign n70128 = ~n70051;
  assign n70168 = n70132 & n18712;
  assign n70169 = ~n70132;
  assign n70172 = ~n70196;
  assign n70214 = n70224 & n70225;
  assign n70230 = n66410 & n69395;
  assign n70183 = ~n70238;
  assign n70229 = n70040 & n70239;
  assign n70222 = n66410 & n69297;
  assign n70219 = ~n70040;
  assign n66499 = ~n66410;
  assign n70261 = ~n70288;
  assign n69837 = ~n68586;
  assign n69970 = n70050 & n70046;
  assign n70072 = n70073 & n10589;
  assign n70009 = ~n70074;
  assign n70042 = n70085 & n70086;
  assign n70081 = n70027 & n70093;
  assign n70057 = n70094 & n70095;
  assign n70075 = n66096 & n68695;
  assign n70091 = n66096 & n70096;
  assign n66112 = ~n66096;
  assign n70092 = ~n70027;
  assign n70036 = ~n70123;
  assign n70122 = n70128 & n67351;
  assign n70101 = ~n70137;
  assign n70140 = ~n70168;
  assign n70162 = n70169 & n252;
  assign n70131 = n70172 & n70173;
  assign n70182 = ~n70214;
  assign n70212 = n66499 & n67826;
  assign n70213 = n70219 & n70084;
  assign n70181 = ~n70222;
  assign n70077 = ~n70229;
  assign n69402 = ~n70230;
  assign n70209 = n66499 & n70234;
  assign n70223 = n70261 & n70262;
  assign n69983 = ~n69970;
  assign n70011 = n70042 ^ n70043;
  assign n70028 = n70057 ^ n70058;
  assign n70044 = ~n70042;
  assign n70045 = ~n70072;
  assign n70037 = ~n70075;
  assign n70055 = ~n70081;
  assign n70070 = n66112 & n68757;
  assign n70056 = ~n70057;
  assign n68771 = ~n70091;
  assign n70061 = n66112 & n67382;
  assign n70065 = n70092 & n70058;
  assign n70082 = n70101 & n70102;
  assign n70090 = ~n70122;
  assign n70100 = n70131 ^ n70132;
  assign n70098 = ~n70162;
  assign n70139 = ~n70131;
  assign n70157 = n70182 & n70183;
  assign n69432 = ~n70209;
  assign n70180 = ~n70212;
  assign n70049 = ~n70213;
  assign n70179 = n70223 ^ n67957;
  assign n69971 = n266 ^ n70011;
  assign n69987 = n70027 ^ n70028;
  assign n70034 = n70044 & n70045;
  assign n70039 = n70055 & n70056;
  assign n70038 = ~n70061;
  assign n70030 = ~n70065;
  assign n68756 = ~n70070;
  assign n70052 = n70082 ^ n67351;
  assign n70089 = ~n70082;
  assign n70064 = n252 ^ n70100;
  assign n70129 = n70139 & n70140;
  assign n70104 = n70157 ^ n70158;
  assign n70150 = ~n70157;
  assign n66460 = n70178 ^ n70179;
  assign n69974 = n70180 & n70181;
  assign n68546 = n69970 ^ n69971;
  assign n69982 = ~n69971;
  assign n69989 = n69987 & n265;
  assign n69992 = ~n69987;
  assign n70008 = ~n70034;
  assign n69965 = n70037 & n70038;
  assign n70029 = ~n70039;
  assign n66020 = n70051 ^ n70052;
  assign n69980 = n70063 ^ n70064;
  assign n70062 = n70089 & n70090;
  assign n70071 = ~n70064;
  assign n70068 = n70103 ^ n70104;
  assign n70097 = ~n70129;
  assign n70119 = n70149 ^ n66460;
  assign n70133 = n70150 & n70151;
  assign n70147 = n66460 & n69315;
  assign n70148 = ~n66460;
  assign n69991 = ~n69974;
  assign n69786 = ~n68546;
  assign n69913 = n69982 & n69983;
  assign n69927 = ~n69989;
  assign n69976 = n69992 & n10522;
  assign n69986 = n70008 & n70009;
  assign n70013 = n66020 & n68714;
  assign n70024 = n69965 & n69994;
  assign n69993 = n70029 & n70030;
  assign n70012 = n66020 & n67346;
  assign n70019 = ~n69965;
  assign n66069 = ~n66020;
  assign n70035 = ~n70062;
  assign n70001 = n70071 & n70063;
  assign n70088 = n70068 & n18693;
  assign n70067 = n70097 & n70098;
  assign n70080 = ~n70068;
  assign n69393 = n70118 ^ n70119;
  assign n70107 = ~n70133;
  assign n70105 = ~n70147;
  assign n70134 = n70148 & n69368;
  assign n69961 = ~n69976;
  assign n69946 = n69986 ^ n69987;
  assign n69966 = n69993 ^ n69994;
  assign n69962 = ~n69986;
  assign n69978 = ~n70012;
  assign n68711 = ~n70013;
  assign n70003 = n70019 & n70020;
  assign n70004 = n66069 & n68621;
  assign n69996 = ~n69993;
  assign n70005 = n66069 & n70021;
  assign n69995 = ~n70024;
  assign n70014 = n70035 & n70036;
  assign n70033 = n70067 ^ n70068;
  assign n70069 = n70080 & n251;
  assign n70059 = ~n70088;
  assign n70060 = ~n70067;
  assign n70083 = n70107 & n70108;
  assign n70106 = ~n70134;
  assign n69920 = n265 ^ n69946;
  assign n69951 = n69961 & n69962;
  assign n69902 = n69965 ^ n69966;
  assign n69972 = n69995 & n69996;
  assign n69964 = ~n70003;
  assign n69979 = ~n70004;
  assign n68734 = ~n70005;
  assign n69981 = n70014 ^ n67271;
  assign n70010 = n70014 & n67348;
  assign n70007 = n251 ^ n70033;
  assign n70023 = ~n70014;
  assign n70053 = n70059 & n70060;
  assign n70032 = ~n70069;
  assign n70041 = n70083 ^ n70084;
  assign n70076 = ~n70083;
  assign n70078 = n70105 & n70106;
  assign n68505 = n69913 ^ n69920;
  assign n69912 = ~n69920;
  assign n69937 = n69902 & n10470;
  assign n69926 = ~n69951;
  assign n69928 = ~n69902;
  assign n69963 = ~n69972;
  assign n69932 = n69978 & n69979;
  assign n65954 = n69980 ^ n69981;
  assign n69907 = n70001 ^ n70007;
  assign n69988 = ~n70010;
  assign n70002 = n70023 & n67271;
  assign n70000 = ~n70007;
  assign n69998 = n70040 ^ n70041;
  assign n70031 = ~n70053;
  assign n70066 = n70076 & n70077;
  assign n70054 = n70078 ^ n70079;
  assign n69748 = ~n68505;
  assign n69848 = n69912 & n69913;
  assign n69901 = n69926 & n69927;
  assign n69916 = n69928 & n264;
  assign n69909 = ~n69937;
  assign n69947 = n65954 & n68687;
  assign n69952 = n65954 & n68565;
  assign n69931 = n69963 & n69964;
  assign n69945 = n69932 & n69904;
  assign n66006 = ~n65954;
  assign n69949 = ~n69932;
  assign n69967 = n69907 & n67249;
  assign n69973 = n69988 & n69980;
  assign n69969 = ~n69907;
  assign n69924 = n70000 & n70001;
  assign n69959 = ~n70002;
  assign n70022 = n69998 & n250;
  assign n69997 = n70031 & n70032;
  assign n70017 = ~n69998;
  assign n69936 = n248 ^ n70054;
  assign n70048 = ~n70066;
  assign n69886 = n69901 ^ n69902;
  assign n69859 = ~n69848;
  assign n69877 = ~n69916;
  assign n69910 = ~n69901;
  assign n69903 = n69931 ^ n69932;
  assign n69930 = ~n69945;
  assign n68692 = ~n69947;
  assign n69939 = n66006 & n69948;
  assign n69940 = n69949 & n69950;
  assign n69929 = ~n69931;
  assign n69942 = n66006 & n67271;
  assign n69922 = ~n69952;
  assign n69900 = ~n69967;
  assign n69955 = n69969 & n67305;
  assign n69958 = ~n69973;
  assign n69960 = n69997 ^ n69998;
  assign n70006 = n70017 & n18624;
  assign n69985 = ~n69997;
  assign n69954 = ~n70022;
  assign n70025 = n70048 & n70049;
  assign n69849 = n264 ^ n69886;
  assign n69857 = n69903 ^ n69904;
  assign n69897 = n69909 & n69910;
  assign n69923 = n69929 & n69930;
  assign n68674 = ~n69939;
  assign n69906 = ~n69940;
  assign n69921 = ~n69942;
  assign n69934 = ~n69955;
  assign n69938 = n69958 & n69959;
  assign n69925 = n250 ^ n69960;
  assign n69984 = ~n70006;
  assign n69975 = n70025 ^ n70016;
  assign n70018 = n70025 & n70026;
  assign n70015 = ~n70025;
  assign n68461 = n69848 ^ n69849;
  assign n69858 = ~n69849;
  assign n69889 = n69857 & n10418;
  assign n69880 = ~n69857;
  assign n69876 = ~n69897;
  assign n69863 = n69921 & n69922;
  assign n69905 = ~n69923;
  assign n69852 = n69924 ^ n69925;
  assign n69908 = n69938 ^ n67249;
  assign n69870 = n69925 & n69924;
  assign n69933 = ~n69938;
  assign n69919 = n69974 ^ n69975;
  assign n69968 = n69984 & n69985;
  assign n69999 = n70015 & n70016;
  assign n69990 = ~n70018;
  assign n69695 = ~n68461;
  assign n69802 = n69858 & n69859;
  assign n69856 = n69876 & n69877;
  assign n69872 = n69880 & n279;
  assign n69854 = ~n69889;
  assign n69898 = n69863 & n69888;
  assign n69887 = n69905 & n69906;
  assign n65909 = n69907 ^ n69908;
  assign n69892 = ~n69863;
  assign n69866 = ~n69852;
  assign n69917 = n69933 & n69934;
  assign n69944 = n69919 & n249;
  assign n69953 = ~n69968;
  assign n69943 = ~n69919;
  assign n69977 = n69990 & n69991;
  assign n69957 = ~n69999;
  assign n69819 = ~n69802;
  assign n69835 = n69856 ^ n69857;
  assign n69834 = ~n69872;
  assign n69855 = ~n69856;
  assign n69864 = n69887 ^ n69888;
  assign n69878 = n65909 & n69890;
  assign n69882 = n65909 & n68574;
  assign n69891 = n69892 & n69893;
  assign n65935 = ~n65909;
  assign n69884 = ~n69898;
  assign n69883 = ~n69887;
  assign n69899 = ~n69917;
  assign n69941 = n69943 & n18560;
  assign n69895 = ~n69944;
  assign n69918 = n69953 & n69954;
  assign n69956 = ~n69977;
  assign n69803 = n279 ^ n69835;
  assign n69845 = n69854 & n69855;
  assign n69811 = n69863 ^ n69864;
  assign n68650 = ~n69878;
  assign n69873 = n65935 & n68630;
  assign n69851 = ~n69882;
  assign n69867 = n69883 & n69884;
  assign n69868 = n65935 & n67249;
  assign n69861 = ~n69891;
  assign n69879 = n69899 & n69900;
  assign n69896 = n69918 ^ n69919;
  assign n69914 = ~n69918;
  assign n69915 = ~n69941;
  assign n69935 = n69956 & n69957;
  assign n68426 = n69802 ^ n69803;
  assign n69765 = n69803 & n69819;
  assign n69829 = n69811 & n10398;
  assign n69836 = ~n69811;
  assign n69833 = ~n69845;
  assign n69860 = ~n69867;
  assign n69850 = ~n69868;
  assign n68629 = ~n69873;
  assign n69853 = n69879 ^ n67200;
  assign n69885 = n69879 & n67264;
  assign n69871 = n249 ^ n69896;
  assign n69881 = ~n69879;
  assign n69911 = n69914 & n69915;
  assign n69875 = n69935 ^ n69936;
  assign n69666 = ~n68426;
  assign n69806 = ~n69829;
  assign n69810 = n69833 & n69834;
  assign n69825 = n69836 & n278;
  assign n69812 = n69850 & n69851;
  assign n65839 = n69852 ^ n69853;
  assign n69830 = n69860 & n69861;
  assign n69799 = n69870 ^ n69871;
  assign n69846 = n69871 & n69870;
  assign n69869 = n69881 & n67200;
  assign n69865 = ~n69885;
  assign n69894 = ~n69911;
  assign n69794 = n69810 ^ n69811;
  assign n69788 = ~n69825;
  assign n69807 = ~n69810;
  assign n69813 = n69830 ^ n69831;
  assign n69827 = n65839 & n67200;
  assign n69832 = n69812 & n69831;
  assign n69828 = n65839 & n68586;
  assign n69838 = ~n69812;
  assign n69818 = ~n69830;
  assign n65885 = ~n65839;
  assign n69843 = n69799 & n67145;
  assign n69844 = ~n69799;
  assign n69862 = n69865 & n69866;
  assign n69841 = ~n69869;
  assign n69874 = n69894 & n69895;
  assign n69766 = n278 ^ n69794;
  assign n69801 = n69806 & n69807;
  assign n69770 = n69812 ^ n69813;
  assign n69809 = ~n69827;
  assign n68589 = ~n69828;
  assign n69826 = n65885 & n68504;
  assign n69817 = ~n69832;
  assign n69823 = n65885 & n69837;
  assign n69824 = n69838 & n69839;
  assign n69815 = ~n69843;
  assign n69842 = n69844 & n67204;
  assign n69840 = ~n69862;
  assign n69847 = n69874 ^ n69875;
  assign n68388 = n69765 ^ n69766;
  assign n69735 = n69766 & n69765;
  assign n69791 = n69770 & n10372;
  assign n69787 = ~n69801;
  assign n69789 = ~n69770;
  assign n69804 = n69817 & n69818;
  assign n68612 = ~n69823;
  assign n69798 = ~n69824;
  assign n69808 = ~n69826;
  assign n69820 = n69840 & n69841;
  assign n69796 = ~n69842;
  assign n69754 = n69846 ^ n69847;
  assign n69621 = ~n68388;
  assign n69769 = n69787 & n69788;
  assign n69785 = n69789 & n277;
  assign n69773 = ~n69791;
  assign n69797 = ~n69804;
  assign n69760 = n69808 & n69809;
  assign n69800 = n69820 ^ n67145;
  assign n69814 = ~n69820;
  assign n69822 = n69754 & n67163;
  assign n69821 = ~n69754;
  assign n69753 = n69769 ^ n69770;
  assign n69772 = ~n69769;
  assign n69752 = ~n69785;
  assign n69790 = n69760 & n69781;
  assign n69780 = n69797 & n69798;
  assign n65775 = n69799 ^ n69800;
  assign n69792 = ~n69760;
  assign n69805 = n69814 & n69815;
  assign n69816 = n69821 & n67089;
  assign n69779 = ~n69822;
  assign n69736 = n277 ^ n69753;
  assign n69764 = n69772 & n69773;
  assign n69761 = n69780 ^ n69781;
  assign n69782 = n65775 & n68450;
  assign n69777 = n65775 & n69786;
  assign n69776 = ~n69790;
  assign n69784 = n69792 & n69793;
  assign n69775 = ~n69780;
  assign n65797 = ~n65775;
  assign n69795 = ~n69805;
  assign n69763 = ~n69816;
  assign n68372 = n69735 ^ n69736;
  assign n69701 = n69736 & n69735;
  assign n69730 = n69760 ^ n69761;
  assign n69751 = ~n69764;
  assign n69768 = n69775 & n69776;
  assign n68572 = ~n69777;
  assign n69758 = ~n69782;
  assign n69771 = n65797 & n68546;
  assign n69774 = n65797 & n67204;
  assign n69757 = ~n69784;
  assign n69783 = n69795 & n69796;
  assign n69586 = ~n68372;
  assign n69739 = n69730 & n10334;
  assign n69729 = n69751 & n69752;
  assign n69740 = ~n69730;
  assign n69756 = ~n69768;
  assign n68545 = ~n69771;
  assign n69759 = ~n69774;
  assign n69755 = n69783 ^ n67089;
  assign n69778 = ~n69783;
  assign n69716 = n69729 ^ n69730;
  assign n69725 = ~n69739;
  assign n69737 = n69740 & n276;
  assign n69726 = ~n69729;
  assign n65644 = n69754 ^ n69755;
  assign n69744 = n69756 & n69757;
  assign n69723 = n69758 & n69759;
  assign n69767 = n69778 & n69779;
  assign n69702 = n276 ^ n69716;
  assign n69717 = n69725 & n69726;
  assign n69715 = ~n69737;
  assign n69724 = n69744 ^ n69745;
  assign n69743 = n65644 & n69748;
  assign n69747 = n69723 & n69750;
  assign n69738 = n65644 & n67089;
  assign n69728 = ~n69744;
  assign n69746 = ~n69723;
  assign n65736 = ~n65644;
  assign n69762 = ~n69767;
  assign n68305 = n69701 ^ n69702;
  assign n69658 = n69702 & n69701;
  assign n69714 = ~n69717;
  assign n69698 = n69723 ^ n69724;
  assign n69720 = ~n69738;
  assign n69732 = n65736 & n68505;
  assign n68510 = ~n69743;
  assign n69734 = n69746 & n69745;
  assign n69731 = n65736 & n68411;
  assign n69727 = ~n69747;
  assign n69749 = n69762 & n69763;
  assign n69552 = ~n68305;
  assign n69705 = n69698 & n275;
  assign n69697 = n69714 & n69715;
  assign n69703 = ~n69698;
  assign n69722 = n69727 & n69728;
  assign n69719 = ~n69731;
  assign n68530 = ~n69732;
  assign n69713 = ~n69734;
  assign n69741 = n69749 & n67026;
  assign n69742 = ~n69749;
  assign n69677 = n69697 ^ n69698;
  assign n69700 = n69703 & n10269;
  assign n69670 = ~n69705;
  assign n69685 = ~n69697;
  assign n69678 = n69719 & n69720;
  assign n69712 = ~n69722;
  assign n69721 = ~n69741;
  assign n69733 = n69742 & n67109;
  assign n69659 = n275 ^ n69677;
  assign n69686 = ~n69700;
  assign n69704 = n69678 & n69690;
  assign n69689 = n69712 & n69713;
  assign n69706 = ~n69678;
  assign n69718 = n69721 & n69708;
  assign n69711 = ~n69733;
  assign n68282 = n69658 ^ n69659;
  assign n69664 = ~n69659;
  assign n69680 = n69685 & n69686;
  assign n69679 = n69689 ^ n69690;
  assign n69693 = ~n69704;
  assign n69699 = n69706 & n69707;
  assign n69694 = ~n69689;
  assign n69710 = ~n69718;
  assign n69709 = n69711 & n69721;
  assign n69505 = ~n68282;
  assign n69610 = n69664 & n69658;
  assign n69646 = n69678 ^ n69679;
  assign n69669 = ~n69680;
  assign n69688 = n69693 & n69694;
  assign n69672 = ~n69699;
  assign n65601 = n69708 ^ n69709;
  assign n69696 = n69710 & n69711;
  assign n69660 = n69646 & n10216;
  assign n69645 = n69669 & n69670;
  assign n69662 = ~n69646;
  assign n69671 = ~n69688;
  assign n69687 = n65601 & n67109;
  assign n69683 = n65601 & n69695;
  assign n69675 = n69696 ^ n66948;
  assign n65649 = ~n65601;
  assign n69691 = ~n69696;
  assign n69630 = n69645 ^ n69646;
  assign n69643 = ~n69660;
  assign n69650 = n69662 & n274;
  assign n69644 = ~n69645;
  assign n69661 = n69671 & n69672;
  assign n65473 = n69675 ^ n69676;
  assign n68460 = ~n69683;
  assign n69682 = n65649 & n68354;
  assign n69681 = n65649 & n68461;
  assign n69668 = ~n69687;
  assign n69684 = n69691 & n69692;
  assign n69611 = n274 ^ n69630;
  assign n69639 = n69643 & n69644;
  assign n69628 = ~n69650;
  assign n69641 = n69661 ^ n69656;
  assign n69665 = n65473 & n66948;
  assign n69657 = n65473 & n69666;
  assign n65568 = ~n65473;
  assign n69636 = ~n69661;
  assign n68484 = ~n69681;
  assign n69667 = ~n69682;
  assign n69673 = ~n69684;
  assign n68197 = n69610 ^ n69611;
  assign n69567 = n69611 & n69610;
  assign n69627 = ~n69639;
  assign n69648 = n65568 & n68315;
  assign n69647 = n65568 & n68426;
  assign n68423 = ~n69657;
  assign n69638 = ~n69665;
  assign n69640 = n69667 & n69668;
  assign n69663 = n69673 & n69674;
  assign n69460 = ~n68197;
  assign n69602 = n69627 & n69628;
  assign n69603 = n69640 ^ n69641;
  assign n68448 = ~n69647;
  assign n69637 = ~n69648;
  assign n69649 = n69640 & n69656;
  assign n69632 = n69663 ^ n66838;
  assign n69652 = ~n69640;
  assign n69654 = ~n69663;
  assign n69589 = n69602 ^ n69603;
  assign n69605 = ~n69602;
  assign n69616 = n69603 & n10199;
  assign n69626 = ~n69603;
  assign n65389 = n69631 ^ n69632;
  assign n69575 = n69637 & n69638;
  assign n69635 = ~n69649;
  assign n69642 = n69652 & n69653;
  assign n69651 = n69654 & n69655;
  assign n69568 = n273 ^ n69589;
  assign n69604 = ~n69616;
  assign n69606 = n69626 & n273;
  assign n69617 = n65389 & n66973;
  assign n69615 = n65389 & n68388;
  assign n69618 = n69575 & n69600;
  assign n65482 = ~n65389;
  assign n69613 = ~n69575;
  assign n69629 = n69635 & n69636;
  assign n69623 = ~n69642;
  assign n69633 = ~n69651;
  assign n68146 = n69567 ^ n69568;
  assign n69529 = n69568 & n69567;
  assign n69596 = n69604 & n69605;
  assign n69588 = ~n69606;
  assign n69607 = n69613 & n69614;
  assign n68384 = ~n69615;
  assign n69594 = ~n69617;
  assign n69591 = ~n69618;
  assign n69612 = n65482 & n68212;
  assign n69609 = n65482 & n69621;
  assign n69622 = ~n69629;
  assign n69619 = n69633 & n69634;
  assign n69429 = ~n68146;
  assign n69524 = ~n69529;
  assign n69587 = ~n69596;
  assign n69579 = ~n69607;
  assign n68413 = ~n69609;
  assign n69593 = ~n69612;
  assign n69595 = n69619 ^ n69620;
  assign n69599 = n69622 & n69623;
  assign n69624 = ~n69619;
  assign n69555 = n69587 & n69588;
  assign n69558 = n69593 & n69594;
  assign n65307 = n69595 ^ n66766;
  assign n69576 = n69599 ^ n69600;
  assign n69601 = n69595 & n66766;
  assign n69592 = ~n69599;
  assign n69608 = n69624 & n69625;
  assign n69556 = n69575 ^ n69576;
  assign n69551 = ~n69555;
  assign n69577 = n65307 & n69586;
  assign n69574 = n69558 & n69544;
  assign n69585 = n65307 & n68191;
  assign n65381 = ~n65307;
  assign n69580 = ~n69558;
  assign n69590 = n69591 & n69592;
  assign n69570 = ~n69601;
  assign n69597 = ~n69608;
  assign n69545 = n69555 ^ n69556;
  assign n69564 = n69556 & n10140;
  assign n69561 = ~n69556;
  assign n69572 = n65381 & n68372;
  assign n69565 = ~n69574;
  assign n68370 = ~n69577;
  assign n69573 = n69580 & n69581;
  assign n69569 = ~n69585;
  assign n69578 = ~n69590;
  assign n69584 = n69597 & n69598;
  assign n69530 = n272 ^ n69545;
  assign n69553 = n69561 & n272;
  assign n69550 = ~n69564;
  assign n69500 = n69569 & n69570;
  assign n68352 = ~n69572;
  assign n69547 = ~n69573;
  assign n69557 = n69578 & n69579;
  assign n69560 = n69584 ^ n66681;
  assign n69582 = ~n69584;
  assign n68072 = n69529 ^ n69530;
  assign n69523 = ~n69530;
  assign n69541 = n69550 & n69551;
  assign n69534 = ~n69553;
  assign n69543 = n69557 ^ n69558;
  assign n65215 = n69559 ^ n69560;
  assign n69512 = ~n69500;
  assign n69566 = ~n69557;
  assign n69571 = n69582 & n69583;
  assign n69372 = ~n68072;
  assign n69464 = n69523 & n69524;
  assign n69533 = ~n69541;
  assign n69507 = n69543 ^ n69544;
  assign n69542 = n65215 & n68111;
  assign n69538 = n65215 & n69552;
  assign n65282 = ~n65215;
  assign n69554 = n69565 & n69566;
  assign n69562 = ~n69571;
  assign n69506 = n69533 & n69534;
  assign n69526 = n69507 & n10097;
  assign n69525 = ~n69507;
  assign n68326 = ~n69538;
  assign n69520 = ~n69542;
  assign n69536 = n65282 & n68305;
  assign n69535 = n65282 & n66681;
  assign n69546 = ~n69554;
  assign n69548 = n69562 & n69563;
  assign n69488 = n69506 ^ n69507;
  assign n69515 = n69525 & n287;
  assign n69508 = ~n69526;
  assign n69509 = ~n69506;
  assign n69521 = ~n69535;
  assign n68308 = ~n69536;
  assign n69531 = n69546 & n69547;
  assign n69518 = n69548 ^ n69549;
  assign n69539 = ~n69548;
  assign n69465 = n287 ^ n69488;
  assign n69496 = n69508 & n69509;
  assign n69485 = ~n69515;
  assign n65136 = n66637 ^ n69518;
  assign n69443 = n69520 & n69521;
  assign n69501 = n69531 ^ n69532;
  assign n69522 = n69531 & n69532;
  assign n69519 = ~n69518;
  assign n69516 = ~n69531;
  assign n69537 = n69539 & n69540;
  assign n69355 = n69464 ^ n69465;
  assign n69470 = ~n69465;
  assign n69484 = ~n69496;
  assign n69450 = n69500 ^ n69501;
  assign n69494 = n69443 & n69510;
  assign n69504 = n65136 & n68282;
  assign n69503 = n65136 & n68038;
  assign n65207 = ~n65136;
  assign n69497 = ~n69443;
  assign n69514 = n69516 & n69517;
  assign n69513 = n69519 & n66743;
  assign n69511 = ~n69522;
  assign n69527 = ~n69537;
  assign n69423 = n69470 & n69464;
  assign n69474 = n69484 & n69485;
  assign n69478 = n69450 & n10065;
  assign n69483 = ~n69450;
  assign n69476 = ~n69494;
  assign n69491 = n69497 & n69467;
  assign n69486 = ~n69503;
  assign n68285 = ~n69504;
  assign n69493 = n65207 & n69505;
  assign n69495 = n69511 & n69512;
  assign n69487 = ~n69513;
  assign n69490 = ~n69514;
  assign n69502 = n69527 & n69528;
  assign n69435 = ~n69423;
  assign n69449 = n286 ^ n69474;
  assign n69468 = ~n69478;
  assign n69469 = ~n69474;
  assign n69477 = n69483 & n286;
  assign n69410 = n69486 & n69487;
  assign n69446 = ~n69491;
  assign n68257 = ~n69493;
  assign n69489 = ~n69495;
  assign n69480 = n69502 ^ n66564;
  assign n69498 = ~n69502;
  assign n69424 = n69449 ^ n69450;
  assign n69454 = n69468 & n69469;
  assign n69473 = n69410 & n69427;
  assign n69448 = ~n69477;
  assign n69471 = ~n69410;
  assign n65084 = n69479 ^ n69480;
  assign n69466 = n69489 & n69490;
  assign n69492 = n69498 & n69499;
  assign n69412 = n69423 ^ n69424;
  assign n69388 = n69424 & n69435;
  assign n69447 = ~n69454;
  assign n69463 = n65084 & n68197;
  assign n69444 = n69466 ^ n69467;
  assign n69461 = n69471 & n69472;
  assign n69462 = n65084 & n66658;
  assign n69433 = ~n69473;
  assign n65128 = ~n65084;
  assign n69475 = ~n69466;
  assign n69481 = ~n69492;
  assign n66125 = n69412 ^ n67220;
  assign n69400 = n69412 & n67222;
  assign n69409 = ~n69412;
  assign n69406 = n69443 ^ n69444;
  assign n69425 = n69447 & n69448;
  assign n69452 = n65128 & n67963;
  assign n69451 = n65128 & n69460;
  assign n69408 = ~n69461;
  assign n69437 = ~n69462;
  assign n68201 = ~n69463;
  assign n69455 = n69475 & n69476;
  assign n69458 = n69481 & n69482;
  assign n69378 = ~n66125;
  assign n69354 = ~n69400;
  assign n69317 = n69409 & n67222;
  assign n69405 = n285 ^ n69425;
  assign n69431 = n69406 & n285;
  assign n69404 = ~n69425;
  assign n69428 = ~n69406;
  assign n68227 = ~n69451;
  assign n69438 = ~n69452;
  assign n69445 = ~n69455;
  assign n69439 = n69458 ^ n69459;
  assign n69456 = ~n69458;
  assign n69376 = n69378 & n68277;
  assign n69389 = n69405 ^ n69406;
  assign n69420 = n69428 & n10044;
  assign n69391 = ~n69431;
  assign n69360 = n69437 & n69438;
  assign n65009 = n66481 ^ n69439;
  assign n69426 = n69445 & n69446;
  assign n69440 = ~n69439;
  assign n69453 = n69456 & n69457;
  assign n69353 = ~n69376;
  assign n69367 = n69388 ^ n69389;
  assign n69387 = ~n69389;
  assign n69403 = ~n69420;
  assign n69415 = n65009 & n67899;
  assign n69411 = n69426 ^ n69427;
  assign n69421 = n65009 & n69429;
  assign n69418 = n69360 & n69430;
  assign n65024 = ~n65009;
  assign n69419 = ~n69360;
  assign n69436 = n69440 & n66571;
  assign n69434 = ~n69426;
  assign n69441 = ~n69453;
  assign n69341 = n69353 & n69354;
  assign n69364 = n69367 & n67099;
  assign n69356 = ~n69367;
  assign n69310 = n69387 & n69388;
  assign n69397 = n69403 & n69404;
  assign n69359 = n69410 ^ n69411;
  assign n69398 = ~n69415;
  assign n69383 = ~n69418;
  assign n69413 = n65024 & n68146;
  assign n69414 = n69419 & n69381;
  assign n68169 = ~n69421;
  assign n69422 = n69433 & n69434;
  assign n69399 = ~n69436;
  assign n69416 = n69441 & n69442;
  assign n69321 = n69341 ^ n69342;
  assign n69343 = ~n69341;
  assign n69351 = n69356 & n67080;
  assign n69330 = ~n69364;
  assign n69309 = ~n69310;
  assign n69379 = n69359 & n9976;
  assign n69390 = ~n69397;
  assign n69385 = ~n69359;
  assign n69318 = n69398 & n69399;
  assign n68139 = ~n69413;
  assign n69366 = ~n69414;
  assign n69396 = n69416 ^ n66410;
  assign n69407 = ~n69422;
  assign n69417 = n69416 & n69432;
  assign n67559 = n295 ^ n69321;
  assign n69146 = n69321 & n295;
  assign n69210 = n69343 & n69344;
  assign n69338 = n69330 & n69317;
  assign n69327 = ~n69351;
  assign n69363 = ~n69379;
  assign n69373 = n69385 & n284;
  assign n69358 = n69390 & n69391;
  assign n69386 = n69318 & n69394;
  assign n64928 = n69395 ^ n69396;
  assign n69384 = ~n69318;
  assign n69380 = n69407 & n69408;
  assign n69401 = ~n69417;
  assign n67584 = ~n67559;
  assign n69316 = n69330 & n69327;
  assign n69326 = ~n69338;
  assign n69337 = n69358 ^ n69359;
  assign n69332 = ~n69373;
  assign n69362 = ~n69358;
  assign n69361 = n69380 ^ n69381;
  assign n69371 = n69384 & n69336;
  assign n69374 = n64928 & n67826;
  assign n69345 = ~n69386;
  assign n69375 = n64928 & n68072;
  assign n64942 = ~n64928;
  assign n69382 = ~n69380;
  assign n69392 = n69401 & n69402;
  assign n65997 = n69316 ^ n69317;
  assign n69320 = n69326 & n69327;
  assign n69311 = n284 ^ n69337;
  assign n69325 = n69360 ^ n69361;
  assign n69347 = n69362 & n69363;
  assign n69313 = ~n69371;
  assign n69370 = n64942 & n69372;
  assign n69369 = n64942 & n66499;
  assign n69348 = ~n69374;
  assign n68087 = ~n69375;
  assign n69377 = n69382 & n69383;
  assign n64875 = n69392 ^ n69393;
  assign n69294 = n65997 & n67080;
  assign n66016 = ~n65997;
  assign n69273 = n69310 ^ n69311;
  assign n69287 = ~n69320;
  assign n69308 = ~n69311;
  assign n69333 = n69325 & n283;
  assign n69331 = ~n69347;
  assign n69334 = ~n69325;
  assign n68059 = n69355 ^ n64875;
  assign n69357 = n64875 & n69368;
  assign n69349 = ~n69369;
  assign n68128 = ~n69370;
  assign n69352 = ~n64875;
  assign n69365 = ~n69377;
  assign n69282 = ~n69294;
  assign n69274 = n69287 ^ n67010;
  assign n69291 = n66016 & n68251;
  assign n69301 = n69273 & n67000;
  assign n69305 = ~n69273;
  assign n69270 = n69308 & n69309;
  assign n69324 = n69331 & n69332;
  assign n69300 = ~n69333;
  assign n69329 = n69334 & n9936;
  assign n69275 = n69348 & n69349;
  assign n69350 = n69352 & n66460;
  assign n69340 = ~n69357;
  assign n69335 = n69365 & n69366;
  assign n65915 = n69273 ^ n69274;
  assign n69281 = ~n69291;
  assign n69286 = ~n69301;
  assign n69292 = n69305 & n67010;
  assign n69285 = ~n69270;
  assign n69303 = n69324 ^ n69325;
  assign n69322 = ~n69324;
  assign n69323 = ~n69329;
  assign n69319 = n69335 ^ n69336;
  assign n69289 = ~n69275;
  assign n69346 = ~n69335;
  assign n69339 = ~n69350;
  assign n69252 = n65915 & n68083;
  assign n65966 = ~n65915;
  assign n69265 = n69281 & n69282;
  assign n69283 = n69286 & n69287;
  assign n69268 = ~n69292;
  assign n69271 = n283 ^ n69303;
  assign n69280 = n69318 ^ n69319;
  assign n69307 = n69322 & n69323;
  assign n69314 = n69339 & n69340;
  assign n69328 = n69345 & n69346;
  assign n69238 = ~n69252;
  assign n69248 = n65966 & n67010;
  assign n69253 = n69265 & n69266;
  assign n69259 = ~n69265;
  assign n69224 = n69270 ^ n69271;
  assign n69267 = ~n69283;
  assign n69284 = ~n69271;
  assign n69295 = n69280 & n282;
  assign n69299 = ~n69307;
  assign n69302 = ~n69280;
  assign n69229 = n69314 ^ n69315;
  assign n69312 = ~n69328;
  assign n69237 = ~n69248;
  assign n69239 = ~n69253;
  assign n69249 = n69259 & n69260;
  assign n69246 = n69267 & n69268;
  assign n69258 = n69224 & n66901;
  assign n69262 = ~n69224;
  assign n69240 = n69284 & n69285;
  assign n69255 = ~n69295;
  assign n69279 = n69299 & n69300;
  assign n69290 = n69302 & n9908;
  assign n69296 = n69312 & n69313;
  assign n69206 = n69237 & n69238;
  assign n69225 = n69246 ^ n66925;
  assign n69244 = n69239 & n69210;
  assign n69227 = ~n69249;
  assign n69233 = ~n69246;
  assign n69223 = ~n69258;
  assign n69251 = n69262 & n66925;
  assign n69247 = ~n69240;
  assign n69256 = n69279 ^ n69280;
  assign n69278 = ~n69290;
  assign n69277 = ~n69279;
  assign n69276 = n69296 ^ n69297;
  assign n69298 = n69296 & n69306;
  assign n69304 = ~n69296;
  assign n69214 = n69206 & n69191;
  assign n65835 = n69224 ^ n69225;
  assign n69217 = ~n69206;
  assign n69232 = n69227 & n69239;
  assign n69226 = ~n69244;
  assign n69234 = ~n69251;
  assign n69241 = n282 ^ n69256;
  assign n69236 = n69275 ^ n69276;
  assign n69269 = n69277 & n69278;
  assign n69288 = ~n69298;
  assign n69293 = n69304 & n69297;
  assign n69207 = n65835 & n66901;
  assign n69208 = ~n69214;
  assign n69212 = n69217 & n69218;
  assign n65892 = ~n65835;
  assign n69205 = n69226 & n69227;
  assign n69211 = ~n69232;
  assign n69231 = n69233 & n69234;
  assign n69180 = n69240 ^ n69241;
  assign n69198 = n69241 & n69247;
  assign n69257 = n69236 & n281;
  assign n69254 = ~n69269;
  assign n69261 = ~n69236;
  assign n69272 = n69288 & n69289;
  assign n69264 = ~n69293;
  assign n69190 = n69205 ^ n69206;
  assign n69188 = ~n69207;
  assign n69201 = n65892 & n68013;
  assign n69202 = n69210 ^ n69211;
  assign n69187 = ~n69212;
  assign n69209 = ~n69205;
  assign n69219 = n69180 & n66796;
  assign n69220 = ~n69180;
  assign n69222 = ~n69231;
  assign n69235 = n69254 & n69255;
  assign n69216 = ~n69257;
  assign n69250 = n69261 & n9894;
  assign n69263 = ~n69272;
  assign n69141 = n69190 ^ n69191;
  assign n69189 = ~n69201;
  assign n69192 = n69202 & n2545;
  assign n69194 = ~n69202;
  assign n69195 = n69208 & n69209;
  assign n69183 = ~n69219;
  assign n69213 = n69220 & n66852;
  assign n69200 = n69222 & n69223;
  assign n69221 = n69235 ^ n69236;
  assign n69243 = ~n69235;
  assign n69242 = ~n69250;
  assign n69245 = n69263 & n69264;
  assign n69168 = n69141 & n2430;
  assign n69173 = ~n69141;
  assign n69148 = n69188 & n69189;
  assign n69176 = ~n69192;
  assign n69185 = n69194 & n294;
  assign n69186 = ~n69195;
  assign n69181 = n69200 ^ n66796;
  assign n69204 = ~n69213;
  assign n69203 = ~n69200;
  assign n69199 = n281 ^ n69221;
  assign n69230 = n69242 & n69243;
  assign n69228 = n280 ^ n69245;
  assign n69142 = ~n69168;
  assign n69163 = n69173 & n293;
  assign n69166 = n69148 & n69172;
  assign n69169 = ~n69148;
  assign n69174 = n69176 & n69146;
  assign n65771 = n69180 ^ n69181;
  assign n69158 = ~n69185;
  assign n69171 = n69186 & n69187;
  assign n69138 = n69198 ^ n69199;
  assign n69193 = n69203 & n69204;
  assign n69178 = n69199 & n69198;
  assign n69197 = n69228 ^ n69229;
  assign n69215 = ~n69230;
  assign n69120 = ~n69163;
  assign n69153 = ~n69166;
  assign n69156 = n65771 & n67930;
  assign n69164 = n69169 & n69170;
  assign n69149 = n69171 ^ n69172;
  assign n69157 = ~n69174;
  assign n65799 = ~n65771;
  assign n69167 = n69176 & n69158;
  assign n69154 = ~n69171;
  assign n69184 = n69138 & n66731;
  assign n69182 = ~n69193;
  assign n69177 = ~n69138;
  assign n69196 = n69215 & n69216;
  assign n69103 = n69148 ^ n69149;
  assign n69150 = n69153 & n69154;
  assign n69145 = ~n69156;
  assign n69140 = n69157 & n69158;
  assign n69135 = ~n69164;
  assign n69155 = n65799 & n66796;
  assign n69147 = ~n69167;
  assign n69175 = n69177 & n66762;
  assign n69159 = n69182 & n69183;
  assign n69162 = ~n69184;
  assign n69179 = n69196 ^ n69197;
  assign n69132 = n69103 & n2338;
  assign n69130 = ~n69103;
  assign n69125 = n69140 ^ n69141;
  assign n69129 = n69146 ^ n69147;
  assign n69134 = ~n69150;
  assign n69143 = ~n69140;
  assign n69144 = ~n69155;
  assign n69139 = n69159 ^ n66731;
  assign n69161 = ~n69159;
  assign n69137 = ~n69175;
  assign n69098 = n69178 ^ n69179;
  assign n69109 = n293 ^ n69125;
  assign n68820 = n69129 ^ n67584;
  assign n69127 = n69130 & n292;
  assign n69106 = ~n69132;
  assign n69108 = n69129 & n67584;
  assign n69114 = n69134 & n69135;
  assign n65681 = n69138 ^ n69139;
  assign n69133 = n69142 & n69143;
  assign n69096 = n69144 & n69145;
  assign n69151 = n69161 & n69162;
  assign n69160 = n69098 & n66648;
  assign n69165 = ~n69098;
  assign n67497 = n69108 ^ n69109;
  assign n69111 = ~n69109;
  assign n69097 = n69114 ^ n69115;
  assign n67552 = ~n68820;
  assign n69088 = ~n69127;
  assign n69128 = n69096 & n69131;
  assign n69121 = n65681 & n67852;
  assign n69112 = ~n69114;
  assign n69119 = ~n69133;
  assign n65701 = ~n65681;
  assign n69126 = ~n69096;
  assign n69136 = ~n69151;
  assign n69105 = ~n69160;
  assign n69152 = n69165 & n66688;
  assign n68772 = ~n67497;
  assign n69066 = n69096 ^ n69097;
  assign n69061 = n69111 & n69108;
  assign n69102 = n69119 & n69120;
  assign n69101 = ~n69121;
  assign n69116 = n69126 & n69115;
  assign n69118 = n65701 & n66762;
  assign n69113 = ~n69128;
  assign n69122 = n69136 & n69137;
  assign n69124 = ~n69152;
  assign n69078 = n69066 & n291;
  assign n69081 = ~n69066;
  assign n69089 = n69102 ^ n69103;
  assign n69110 = n69112 & n69113;
  assign n69093 = ~n69116;
  assign n69107 = ~n69102;
  assign n69100 = ~n69118;
  assign n69099 = n69122 ^ n66648;
  assign n69123 = ~n69122;
  assign n69044 = ~n69078;
  assign n69073 = n69081 & n2210;
  assign n69062 = n292 ^ n69089;
  assign n65586 = n69098 ^ n69099;
  assign n69057 = n69100 & n69101;
  assign n69095 = n69106 & n69107;
  assign n69092 = ~n69110;
  assign n69117 = n69123 & n69124;
  assign n67466 = n69061 ^ n69062;
  assign n69059 = ~n69073;
  assign n69067 = ~n69062;
  assign n69076 = n69092 & n69093;
  assign n69090 = n65586 & n67782;
  assign n69091 = n69057 & n69094;
  assign n69086 = ~n69057;
  assign n65619 = ~n65586;
  assign n69087 = ~n69095;
  assign n69104 = ~n69117;
  assign n68738 = ~n67466;
  assign n69032 = n69067 & n69061;
  assign n69058 = n69076 ^ n69077;
  assign n69074 = ~n69076;
  assign n69079 = n69086 & n69077;
  assign n69065 = n69087 & n69088;
  assign n69082 = n65619 & n66648;
  assign n69070 = ~n69090;
  assign n69075 = ~n69091;
  assign n69085 = n69104 & n69105;
  assign n69022 = n69057 ^ n69058;
  assign n69026 = ~n69032;
  assign n69046 = n69065 ^ n69066;
  assign n69072 = n69074 & n69075;
  assign n69056 = ~n69079;
  assign n69060 = ~n69065;
  assign n69071 = ~n69082;
  assign n69069 = n69085 ^ n66559;
  assign n69083 = ~n69085;
  assign n69037 = n69022 & n290;
  assign n69040 = ~n69022;
  assign n69033 = n291 ^ n69046;
  assign n69054 = n69059 & n69060;
  assign n65502 = n69068 ^ n69069;
  assign n69019 = n69070 & n69071;
  assign n69055 = ~n69072;
  assign n69080 = n69083 & n69084;
  assign n67430 = n69032 ^ n69033;
  assign n68996 = ~n69037;
  assign n69031 = n69040 & n2109;
  assign n69025 = ~n69033;
  assign n69049 = n65502 & n66594;
  assign n69043 = ~n69054;
  assign n69038 = n69055 & n69056;
  assign n69053 = n69019 & n69039;
  assign n65555 = ~n65502;
  assign n69047 = ~n69019;
  assign n69063 = ~n69080;
  assign n68702 = ~n67430;
  assign n68984 = n69025 & n69026;
  assign n69017 = ~n69031;
  assign n69020 = n69038 ^ n69039;
  assign n69021 = n69043 & n69044;
  assign n69035 = ~n69038;
  assign n69041 = n69047 & n69048;
  assign n69024 = ~n69049;
  assign n69045 = n65555 & n67747;
  assign n69036 = ~n69053;
  assign n69050 = n69063 & n69064;
  assign n68983 = n69019 ^ n69020;
  assign n69004 = n69021 ^ n69022;
  assign n68991 = ~n68984;
  assign n69034 = n69035 & n69036;
  assign n69018 = ~n69021;
  assign n69016 = ~n69041;
  assign n69023 = ~n69045;
  assign n69028 = n69050 ^ n66492;
  assign n69051 = ~n69050;
  assign n68997 = n68983 & n2069;
  assign n68985 = n290 ^ n69004;
  assign n69002 = ~n68983;
  assign n69014 = n69017 & n69018;
  assign n68980 = n69023 & n69024;
  assign n65408 = n69027 ^ n69028;
  assign n69015 = ~n69034;
  assign n69042 = n69051 & n69052;
  assign n67406 = n68984 ^ n68985;
  assign n68939 = n68985 & n68991;
  assign n68979 = ~n68997;
  assign n68990 = n69002 & n289;
  assign n68995 = ~n69014;
  assign n69011 = n65408 & n66492;
  assign n69009 = n68980 & n68999;
  assign n68998 = n69015 & n69016;
  assign n69007 = ~n68980;
  assign n65454 = ~n65408;
  assign n69029 = ~n69042;
  assign n68657 = ~n67406;
  assign n68948 = ~n68939;
  assign n68957 = ~n68990;
  assign n68982 = n68995 & n68996;
  assign n68981 = n68998 ^ n68999;
  assign n69003 = n69007 & n69008;
  assign n69001 = ~n69009;
  assign n68987 = ~n69011;
  assign n69005 = n65454 & n67678;
  assign n69000 = ~n68998;
  assign n69010 = n69029 & n69030;
  assign n68936 = n68980 ^ n68981;
  assign n68961 = n68982 ^ n68983;
  assign n68978 = ~n68982;
  assign n68994 = n69000 & n69001;
  assign n68977 = ~n69003;
  assign n68986 = ~n69005;
  assign n68993 = n69010 ^ n66420;
  assign n69012 = ~n69010;
  assign n68940 = n289 ^ n68961;
  assign n68960 = n68936 & n2009;
  assign n68964 = ~n68936;
  assign n68974 = n68978 & n68979;
  assign n68945 = n68986 & n68987;
  assign n65328 = n68992 ^ n68993;
  assign n68976 = ~n68994;
  assign n69006 = n69012 & n69013;
  assign n67352 = n68939 ^ n68940;
  assign n68898 = n68940 & n68948;
  assign n68938 = ~n68960;
  assign n68950 = n68964 & n288;
  assign n68956 = ~n68974;
  assign n68969 = n68945 & n68963;
  assign n68973 = n65328 & n66440;
  assign n68962 = n68976 & n68977;
  assign n65373 = ~n65328;
  assign n68971 = ~n68945;
  assign n68988 = ~n69006;
  assign n68614 = ~n67352;
  assign n68905 = ~n68898;
  assign n68924 = ~n68950;
  assign n68935 = n68956 & n68957;
  assign n68946 = n68962 ^ n68963;
  assign n68959 = ~n68969;
  assign n68958 = ~n68962;
  assign n68967 = n68971 & n68972;
  assign n68952 = ~n68973;
  assign n68965 = n65373 & n67640;
  assign n68975 = n68988 & n68989;
  assign n68918 = n68935 ^ n68936;
  assign n68903 = n68945 ^ n68946;
  assign n68937 = ~n68935;
  assign n68955 = n68958 & n68959;
  assign n68953 = ~n68965;
  assign n68942 = ~n68967;
  assign n68968 = n68975 & n66382;
  assign n68970 = ~n68975;
  assign n68899 = n288 ^ n68918;
  assign n68921 = n68903 & n1922;
  assign n68922 = ~n68903;
  assign n68934 = n68937 & n68938;
  assign n68906 = n68952 & n68953;
  assign n68941 = ~n68955;
  assign n68954 = ~n68968;
  assign n68966 = n68970 & n66357;
  assign n67319 = n68898 ^ n68899;
  assign n68904 = ~n68899;
  assign n68912 = ~n68921;
  assign n68915 = n68922 & n303;
  assign n68923 = ~n68934;
  assign n68919 = n68941 & n68942;
  assign n68932 = n68906 & n68947;
  assign n68933 = ~n68906;
  assign n68951 = n68954 & n68929;
  assign n68944 = ~n68966;
  assign n68569 = ~n67319;
  assign n68867 = n68904 & n68905;
  assign n68887 = ~n68915;
  assign n68907 = n68919 ^ n68920;
  assign n68902 = n68923 & n68924;
  assign n68926 = ~n68932;
  assign n68931 = n68933 & n68920;
  assign n68925 = ~n68919;
  assign n68943 = ~n68951;
  assign n68949 = n68944 & n68954;
  assign n68892 = n68902 ^ n68903;
  assign n68861 = n68906 ^ n68907;
  assign n68911 = ~n68902;
  assign n68916 = n68925 & n68926;
  assign n68901 = ~n68931;
  assign n68917 = n68943 & n68944;
  assign n68930 = ~n68949;
  assign n68868 = n303 ^ n68892;
  assign n68891 = n68861 & n302;
  assign n68888 = ~n68861;
  assign n68895 = n68911 & n68912;
  assign n68900 = ~n68916;
  assign n68896 = n68917 ^ n66320;
  assign n65240 = n68929 ^ n68930;
  assign n68927 = ~n68917;
  assign n67276 = n68867 ^ n68868;
  assign n68871 = ~n68868;
  assign n68882 = n68888 & n1874;
  assign n68849 = ~n68891;
  assign n68886 = ~n68895;
  assign n65162 = n68896 ^ n68897;
  assign n68883 = n68900 & n68901;
  assign n68913 = n65240 & n67591;
  assign n65268 = ~n65240;
  assign n68914 = n68927 & n68928;
  assign n68528 = ~n67276;
  assign n68834 = n68871 & n68867;
  assign n68875 = ~n68882;
  assign n68870 = n68883 ^ n68880;
  assign n68860 = n68886 & n68887;
  assign n68890 = n65162 & n67545;
  assign n65183 = ~n65162;
  assign n68858 = ~n68883;
  assign n68894 = ~n68913;
  assign n68910 = n65268 & n66357;
  assign n68908 = ~n68914;
  assign n68854 = n68860 ^ n68861;
  assign n68874 = ~n68860;
  assign n68879 = n65183 & n66308;
  assign n68862 = ~n68890;
  assign n68889 = n68908 & n68909;
  assign n68893 = ~n68910;
  assign n68835 = n302 ^ n68854;
  assign n68859 = n68874 & n68875;
  assign n68863 = ~n68879;
  assign n68866 = n68889 ^ n66225;
  assign n68869 = n68893 & n68894;
  assign n68884 = ~n68889;
  assign n67232 = n68834 ^ n68835;
  assign n68794 = n68835 & n68834;
  assign n68848 = ~n68859;
  assign n68806 = n68862 & n68863;
  assign n65061 = n68865 ^ n68866;
  assign n68827 = n68869 ^ n68870;
  assign n68876 = n68869 & n68880;
  assign n68881 = n68884 & n68885;
  assign n68877 = ~n68869;
  assign n68491 = ~n67232;
  assign n68826 = n68848 & n68849;
  assign n68855 = n68827 & n1851;
  assign n68852 = n68806 & n68823;
  assign n68850 = n65061 & n66225;
  assign n68844 = ~n68806;
  assign n68851 = ~n68827;
  assign n65125 = ~n65061;
  assign n68857 = ~n68876;
  assign n68864 = n68877 & n68878;
  assign n68872 = ~n68881;
  assign n68812 = n68826 ^ n68827;
  assign n68828 = ~n68826;
  assign n68842 = n68844 & n68845;
  assign n68837 = ~n68850;
  assign n68843 = n68851 & n301;
  assign n68824 = ~n68852;
  assign n68841 = n65125 & n67516;
  assign n68829 = ~n68855;
  assign n68856 = n68857 & n68858;
  assign n68839 = ~n68864;
  assign n68853 = n68872 & n68873;
  assign n68795 = n301 ^ n68812;
  assign n68821 = n68828 & n68829;
  assign n68836 = ~n68841;
  assign n68804 = ~n68842;
  assign n68809 = ~n68843;
  assign n68831 = n68853 ^ n66193;
  assign n68838 = ~n68856;
  assign n68846 = ~n68853;
  assign n67178 = n68794 ^ n68795;
  assign n68793 = ~n68795;
  assign n68808 = ~n68821;
  assign n64979 = n68830 ^ n68831;
  assign n68766 = n68836 & n68837;
  assign n68822 = n68838 & n68839;
  assign n68840 = n68846 & n68847;
  assign n68451 = ~n67178;
  assign n68744 = n68793 & n68794;
  assign n68783 = n68808 & n68809;
  assign n68815 = n64979 & n68820;
  assign n68816 = n64979 & n67486;
  assign n68811 = n68766 & n68786;
  assign n68813 = ~n68766;
  assign n68807 = n68822 ^ n68823;
  assign n65013 = ~n64979;
  assign n68825 = ~n68822;
  assign n68832 = ~n68840;
  assign n68759 = ~n68744;
  assign n68777 = ~n68783;
  assign n68784 = n68806 ^ n68807;
  assign n68788 = ~n68811;
  assign n68802 = n65013 & n67552;
  assign n68801 = n65013 & n66209;
  assign n68800 = n68813 & n68814;
  assign n67555 = ~n68815;
  assign n68791 = ~n68816;
  assign n68819 = n68824 & n68825;
  assign n68810 = n68832 & n68833;
  assign n68761 = n68783 ^ n68784;
  assign n68787 = n68784 & n1797;
  assign n68790 = ~n68784;
  assign n68769 = ~n68800;
  assign n68792 = ~n68801;
  assign n67535 = ~n68802;
  assign n68797 = n68810 ^ n66152;
  assign n68803 = ~n68819;
  assign n68817 = ~n68810;
  assign n68745 = n300 ^ n68761;
  assign n68776 = ~n68787;
  assign n68782 = n68790 & n300;
  assign n68724 = n68791 & n68792;
  assign n64906 = n68796 ^ n68797;
  assign n68785 = n68803 & n68804;
  assign n68805 = n68817 & n68818;
  assign n67132 = n68744 ^ n68745;
  assign n68688 = n68745 & n68759;
  assign n68763 = n68776 & n68777;
  assign n68773 = n64906 & n67497;
  assign n68775 = n68724 & n68780;
  assign n68752 = ~n68782;
  assign n68779 = n64906 & n66152;
  assign n68778 = ~n68724;
  assign n68767 = n68785 ^ n68786;
  assign n64944 = ~n64906;
  assign n68789 = ~n68785;
  assign n68798 = ~n68805;
  assign n68416 = ~n67132;
  assign n68700 = ~n68688;
  assign n68751 = ~n68763;
  assign n68717 = n68766 ^ n68767;
  assign n68760 = n64944 & n68772;
  assign n68762 = n64944 & n67429;
  assign n67502 = ~n68773;
  assign n68749 = ~n68775;
  assign n68765 = n68778 & n68748;
  assign n68754 = ~n68779;
  assign n68781 = n68788 & n68789;
  assign n68774 = n68798 & n68799;
  assign n68731 = n68751 & n68752;
  assign n68743 = n68717 & n1764;
  assign n68746 = ~n68717;
  assign n67520 = ~n68760;
  assign n68753 = ~n68762;
  assign n68728 = ~n68765;
  assign n68758 = n68774 ^ n66096;
  assign n68768 = ~n68781;
  assign n68770 = ~n68774;
  assign n68716 = n299 ^ n68731;
  assign n68736 = ~n68743;
  assign n68742 = n68746 & n299;
  assign n68737 = ~n68731;
  assign n68676 = n68753 & n68754;
  assign n64851 = n68757 ^ n68758;
  assign n68747 = n68768 & n68769;
  assign n68764 = n68770 & n68771;
  assign n68689 = n68716 ^ n68717;
  assign n68721 = n68736 & n68737;
  assign n68735 = n68676 & n68706;
  assign n68713 = ~n68742;
  assign n68730 = n64851 & n67466;
  assign n68732 = n64851 & n66112;
  assign n68725 = n68747 ^ n68748;
  assign n68739 = ~n68676;
  assign n64865 = ~n64851;
  assign n68750 = ~n68747;
  assign n68755 = ~n68764;
  assign n67068 = n68688 ^ n68689;
  assign n68699 = ~n68689;
  assign n68712 = ~n68721;
  assign n68698 = n68724 ^ n68725;
  assign n67461 = ~n68730;
  assign n68726 = n64865 & n67382;
  assign n68719 = ~n68732;
  assign n68708 = ~n68735;
  assign n68723 = n64865 & n68738;
  assign n68720 = n68739 & n68740;
  assign n68741 = n68749 & n68750;
  assign n68729 = n68755 & n68756;
  assign n68364 = ~n67068;
  assign n68651 = n68699 & n68700;
  assign n68697 = n68712 & n68713;
  assign n68707 = n68698 & n298;
  assign n68704 = ~n68698;
  assign n68679 = ~n68720;
  assign n67484 = ~n68723;
  assign n68718 = ~n68726;
  assign n68715 = n68729 ^ n66020;
  assign n68727 = ~n68741;
  assign n68733 = ~n68729;
  assign n68669 = n68697 ^ n68698;
  assign n68701 = n68704 & n1703;
  assign n68667 = ~n68707;
  assign n68680 = ~n68697;
  assign n64755 = n68714 ^ n68715;
  assign n68635 = n68718 & n68719;
  assign n68705 = n68727 & n68728;
  assign n68722 = n68733 & n68734;
  assign n68652 = n298 ^ n68669;
  assign n68681 = ~n68701;
  assign n68690 = n64755 & n68702;
  assign n68693 = n68635 & n68661;
  assign n68696 = n64755 & n67346;
  assign n68677 = n68705 ^ n68706;
  assign n68694 = ~n68635;
  assign n64793 = ~n64755;
  assign n68709 = ~n68705;
  assign n68710 = ~n68722;
  assign n67041 = n68651 ^ n68652;
  assign n68597 = n68652 & n68651;
  assign n68645 = n68676 ^ n68677;
  assign n68675 = n68680 & n68681;
  assign n67447 = ~n68690;
  assign n68685 = n64793 & n67430;
  assign n68684 = n64793 & n66020;
  assign n68662 = ~n68693;
  assign n68683 = n68694 & n68695;
  assign n68671 = ~n68696;
  assign n68703 = n68708 & n68709;
  assign n68686 = n68710 & n68711;
  assign n68337 = ~n67041;
  assign n68659 = n68645 & n1678;
  assign n68665 = ~n68645;
  assign n68666 = ~n68675;
  assign n68641 = ~n68683;
  assign n68670 = ~n68684;
  assign n67436 = ~n68685;
  assign n68672 = n68686 ^ n68687;
  assign n68678 = ~n68703;
  assign n68691 = ~n68686;
  assign n68638 = ~n68659;
  assign n68655 = n68665 & n297;
  assign n68644 = n68666 & n68667;
  assign n68603 = n68670 & n68671;
  assign n64707 = n65954 ^ n68672;
  assign n68668 = ~n68672;
  assign n68660 = n68678 & n68679;
  assign n68682 = n68691 & n68692;
  assign n68619 = n68644 ^ n68645;
  assign n68624 = ~n68655;
  assign n68637 = ~n68644;
  assign n68647 = n64707 & n68657;
  assign n68654 = n64707 & n67271;
  assign n68646 = n68603 & n68658;
  assign n64745 = ~n64707;
  assign n68636 = n68660 ^ n68661;
  assign n68648 = ~n68603;
  assign n68664 = n68668 & n66006;
  assign n68663 = ~n68660;
  assign n68673 = ~n68682;
  assign n68598 = n297 ^ n68619;
  assign n68594 = n68635 ^ n68636;
  assign n68632 = n68637 & n68638;
  assign n68626 = ~n68646;
  assign n67408 = ~n68647;
  assign n68643 = n68648 & n68621;
  assign n68642 = n64745 & n67406;
  assign n68633 = ~n68654;
  assign n68656 = n68662 & n68663;
  assign n68634 = ~n68664;
  assign n68653 = n68673 & n68674;
  assign n66929 = n68597 ^ n68598;
  assign n68606 = ~n68598;
  assign n68625 = n68594 & n1618;
  assign n68623 = ~n68632;
  assign n68618 = ~n68594;
  assign n68582 = n68633 & n68634;
  assign n67394 = ~n68642;
  assign n68601 = ~n68643;
  assign n68631 = n68653 ^ n65909;
  assign n68640 = ~n68656;
  assign n68649 = ~n68653;
  assign n68288 = ~n66929;
  assign n68553 = n68606 & n68597;
  assign n68615 = n68618 & n296;
  assign n68617 = n68582 & n68622;
  assign n68593 = n68623 & n68624;
  assign n68596 = ~n68625;
  assign n68616 = ~n68582;
  assign n64689 = n68630 ^ n68631;
  assign n68620 = n68640 & n68641;
  assign n68639 = n68649 & n68650;
  assign n68580 = n68593 ^ n68594;
  assign n68608 = n64689 & n68614;
  assign n68595 = ~n68593;
  assign n68609 = n64689 & n65935;
  assign n68584 = ~n68615;
  assign n68607 = n68616 & n68565;
  assign n68577 = ~n68617;
  assign n68604 = n68620 ^ n68621;
  assign n64697 = ~n64689;
  assign n68627 = ~n68620;
  assign n68628 = ~n68639;
  assign n68554 = n296 ^ n68580;
  assign n68592 = n68595 & n68596;
  assign n68552 = n68603 ^ n68604;
  assign n68556 = ~n68607;
  assign n67355 = ~n68608;
  assign n68590 = ~n68609;
  assign n68602 = n64697 & n67352;
  assign n68599 = n64697 & n67249;
  assign n68613 = n68626 & n68627;
  assign n68610 = n68628 & n68629;
  assign n66896 = n68553 ^ n68554;
  assign n68557 = ~n68554;
  assign n68585 = n68552 & n311;
  assign n68583 = ~n68592;
  assign n68579 = ~n68552;
  assign n68591 = ~n68599;
  assign n67375 = ~n68602;
  assign n68587 = n68610 ^ n65839;
  assign n68600 = ~n68613;
  assign n68611 = ~n68610;
  assign n68232 = ~n66896;
  assign n68516 = n68557 & n68553;
  assign n68575 = n68579 & n1559;
  assign n68551 = n68583 & n68584;
  assign n68536 = ~n68585;
  assign n64634 = n68586 ^ n68587;
  assign n68523 = n68590 & n68591;
  assign n68581 = n68600 & n68601;
  assign n68605 = n68611 & n68612;
  assign n68526 = ~n68516;
  assign n68537 = n68551 ^ n68552;
  assign n68568 = n68523 & n68543;
  assign n68566 = n64634 & n67200;
  assign n68560 = ~n68551;
  assign n68567 = n64634 & n67319;
  assign n68561 = ~n68575;
  assign n68573 = ~n68523;
  assign n68564 = n68581 ^ n68582;
  assign n64653 = ~n64634;
  assign n68578 = ~n68581;
  assign n68588 = ~n68605;
  assign n68517 = n311 ^ n68537;
  assign n68550 = n68560 & n68561;
  assign n68521 = n68564 ^ n68565;
  assign n68563 = n64653 & n65839;
  assign n68548 = ~n68566;
  assign n67335 = ~n68567;
  assign n68540 = ~n68568;
  assign n68559 = n64653 & n68569;
  assign n68558 = n68573 & n68574;
  assign n68576 = n68577 & n68578;
  assign n68570 = n68588 & n68589;
  assign n66772 = n68516 ^ n68517;
  assign n68525 = ~n68517;
  assign n68538 = n68521 & n310;
  assign n68541 = ~n68521;
  assign n68535 = ~n68550;
  assign n68519 = ~n68558;
  assign n67317 = ~n68559;
  assign n68549 = ~n68563;
  assign n68547 = n68570 ^ n65775;
  assign n68555 = ~n68576;
  assign n68571 = ~n68570;
  assign n68185 = ~n66772;
  assign n68475 = n68525 & n68526;
  assign n68520 = n68535 & n68536;
  assign n68500 = ~n68538;
  assign n68534 = n68541 & n1507;
  assign n64596 = n68546 ^ n68547;
  assign n68478 = n68548 & n68549;
  assign n68542 = n68555 & n68556;
  assign n68562 = n68571 & n68572;
  assign n68497 = n68520 ^ n68521;
  assign n68515 = ~n68520;
  assign n68531 = n64596 & n67276;
  assign n68532 = n64596 & n65797;
  assign n68514 = ~n68534;
  assign n68487 = ~n68478;
  assign n64620 = ~n64596;
  assign n68524 = n68542 ^ n68543;
  assign n68539 = ~n68542;
  assign n68544 = ~n68562;
  assign n68476 = n310 ^ n68497;
  assign n68511 = n68514 & n68515;
  assign n68474 = n68523 ^ n68524;
  assign n68522 = n64620 & n68528;
  assign n67274 = ~n68531;
  assign n68512 = n64620 & n67204;
  assign n68508 = ~n68532;
  assign n68533 = n68539 & n68540;
  assign n68527 = n68544 & n68545;
  assign n66691 = n68475 ^ n68476;
  assign n68477 = ~n68476;
  assign n68502 = n68474 & n1450;
  assign n68499 = ~n68511;
  assign n68501 = ~n68474;
  assign n68507 = ~n68512;
  assign n67303 = ~n68522;
  assign n68506 = n68527 ^ n65644;
  assign n68518 = ~n68533;
  assign n68529 = ~n68527;
  assign n68124 = ~n66691;
  assign n68436 = n68477 & n68475;
  assign n68473 = n68499 & n68500;
  assign n68492 = n68501 & n309;
  assign n68468 = ~n68502;
  assign n64559 = n68505 ^ n68506;
  assign n68424 = n68507 & n68508;
  assign n68495 = n68518 & n68519;
  assign n68513 = n68529 & n68530;
  assign n68441 = ~n68436;
  assign n68458 = n68473 ^ n68474;
  assign n68489 = n64559 & n68491;
  assign n68455 = ~n68492;
  assign n68488 = n64559 & n65644;
  assign n68469 = ~n68473;
  assign n68490 = n68424 & n68494;
  assign n68479 = n68495 ^ n68496;
  assign n64578 = ~n64559;
  assign n68485 = ~n68424;
  assign n68498 = n68495 & n68496;
  assign n68503 = ~n68495;
  assign n68509 = ~n68513;
  assign n68437 = n309 ^ n68458;
  assign n68467 = n68468 & n68469;
  assign n68439 = n68478 ^ n68479;
  assign n68480 = n64578 & n67089;
  assign n68470 = n68485 & n68450;
  assign n68463 = ~n68488;
  assign n68471 = n64578 & n67232;
  assign n67231 = ~n68489;
  assign n68446 = ~n68490;
  assign n68486 = ~n68498;
  assign n68493 = n68503 & n68504;
  assign n68482 = n68509 & n68510;
  assign n66610 = n68436 ^ n68437;
  assign n68440 = ~n68437;
  assign n68457 = n68439 & n1423;
  assign n68454 = ~n68467;
  assign n68456 = ~n68439;
  assign n68421 = ~n68470;
  assign n67258 = ~n68471;
  assign n68464 = ~n68480;
  assign n68462 = n68482 ^ n65601;
  assign n68481 = n68486 & n68487;
  assign n68466 = ~n68493;
  assign n68483 = ~n68482;
  assign n68052 = ~n66610;
  assign n68022 = n68440 & n68441;
  assign n68438 = n68454 & n68455;
  assign n68453 = n68456 & n308;
  assign n68434 = ~n68457;
  assign n64527 = n68461 ^ n68462;
  assign n68381 = n68463 & n68464;
  assign n68465 = ~n68481;
  assign n68472 = n68483 & n68484;
  assign n68400 = ~n68022;
  assign n68419 = n68438 ^ n68439;
  assign n68433 = ~n68438;
  assign n68443 = n64527 & n67178;
  assign n68444 = n64527 & n65601;
  assign n68418 = ~n68453;
  assign n64539 = ~n64527;
  assign n68391 = ~n68381;
  assign n68449 = n68465 & n68466;
  assign n68459 = ~n68472;
  assign n67981 = n308 ^ n68419;
  assign n68430 = n68433 & n68434;
  assign n67181 = ~n68443;
  assign n68428 = ~n68444;
  assign n68425 = n68449 ^ n68450;
  assign n68435 = n64539 & n68451;
  assign n68431 = n64539 & n67109;
  assign n68445 = ~n68449;
  assign n68452 = n68459 & n68460;
  assign n68357 = n67981 & n68400;
  assign n68398 = n68424 ^ n68425;
  assign n68417 = ~n68430;
  assign n68429 = ~n68431;
  assign n67209 = ~n68435;
  assign n68442 = n68445 & n68446;
  assign n68427 = n68452 ^ n65473;
  assign n68447 = ~n68452;
  assign n68402 = n68398 & n307;
  assign n68403 = ~n68398;
  assign n68397 = n68417 & n68418;
  assign n64471 = n68426 ^ n68427;
  assign n68332 = n68428 & n68429;
  assign n68420 = ~n68442;
  assign n68432 = n68447 & n68448;
  assign n68378 = n68397 ^ n68398;
  assign n68367 = ~n68402;
  assign n68395 = n68403 & n1356;
  assign n68407 = n68332 & n68415;
  assign n68406 = n64471 & n65473;
  assign n68414 = n64471 & n68416;
  assign n68387 = ~n68397;
  assign n64476 = ~n64471;
  assign n68408 = ~n68332;
  assign n68404 = n68420 & n68421;
  assign n68422 = ~n68432;
  assign n68358 = n307 ^ n68378;
  assign n68386 = ~n68395;
  assign n68382 = n68404 ^ n68405;
  assign n68392 = n64476 & n67132;
  assign n68379 = ~n68406;
  assign n68356 = ~n68407;
  assign n68393 = n68408 & n68354;
  assign n68394 = n64476 & n66948;
  assign n67128 = ~n68414;
  assign n68409 = n68404 & n68405;
  assign n68410 = ~n68404;
  assign n68401 = n68422 & n68423;
  assign n68338 = n68357 ^ n68358;
  assign n68363 = ~n68358;
  assign n68343 = n68381 ^ n68382;
  assign n68377 = n68386 & n68387;
  assign n67158 = ~n68392;
  assign n68335 = ~n68393;
  assign n68380 = ~n68394;
  assign n68389 = n68401 ^ n65389;
  assign n68390 = ~n68409;
  assign n68396 = n68410 & n68411;
  assign n68412 = ~n68401;
  assign n64198 = n68338 ^ n66125;
  assign n68339 = n68338 & n66125;
  assign n68341 = ~n68338;
  assign n68299 = n68363 & n68357;
  assign n68373 = n68343 & n1286;
  assign n68368 = ~n68343;
  assign n68366 = ~n68377;
  assign n68291 = n68379 & n68380;
  assign n64408 = n68388 ^ n68389;
  assign n68385 = n68390 & n68391;
  assign n68376 = ~n68396;
  assign n68399 = n68412 & n68413;
  assign n68317 = n64198 & n67222;
  assign n64200 = ~n64198;
  assign n68310 = ~n68339;
  assign n68220 = n68341 & n66125;
  assign n68342 = n68366 & n68367;
  assign n68359 = n68368 & n306;
  assign n68350 = ~n68373;
  assign n68374 = n64408 & n67068;
  assign n68365 = n64408 & n66973;
  assign n68296 = ~n68291;
  assign n64457 = ~n64408;
  assign n68375 = ~n68385;
  assign n68383 = ~n68399;
  assign n68309 = ~n68317;
  assign n68323 = n68342 ^ n68343;
  assign n68349 = ~n68342;
  assign n68328 = ~n68359;
  assign n68362 = n64457 & n68364;
  assign n68360 = n64457 & n65389;
  assign n68348 = ~n68365;
  assign n67101 = ~n68374;
  assign n68353 = n68375 & n68376;
  assign n68371 = n68383 & n68384;
  assign n68286 = n68309 & n68310;
  assign n68300 = n306 ^ n68323;
  assign n68340 = n68349 & n68350;
  assign n68333 = n68353 ^ n68354;
  assign n68347 = ~n68360;
  assign n67066 = ~n68362;
  assign n68355 = ~n68353;
  assign n68346 = n68371 ^ n68372;
  assign n68369 = ~n68371;
  assign n68249 = n68286 ^ n68287;
  assign n68276 = ~n68286;
  assign n68294 = n68299 ^ n68300;
  assign n68258 = n68300 & n68299;
  assign n68304 = n68332 ^ n68333;
  assign n68327 = ~n68340;
  assign n64361 = n65307 ^ n68346;
  assign n68241 = n68347 & n68348;
  assign n68344 = n68355 & n68356;
  assign n68345 = n68346 & n65381;
  assign n68361 = n68369 & n68370;
  assign n66116 = n327 ^ n68249;
  assign n68104 = n68249 & n327;
  assign n68250 = n68276 & n68277;
  assign n68275 = n68294 & n65997;
  assign n68279 = ~n68294;
  assign n68267 = ~n68258;
  assign n68312 = n68304 & n305;
  assign n68303 = n68327 & n68328;
  assign n68313 = ~n68304;
  assign n68324 = n68241 & n68336;
  assign n68331 = n64361 & n68337;
  assign n68329 = ~n68241;
  assign n64410 = ~n64361;
  assign n68334 = ~n68344;
  assign n68302 = ~n68345;
  assign n68351 = ~n68361;
  assign n67378 = ~n66116;
  assign n68234 = n68104 & n326;
  assign n68235 = ~n68104;
  assign n68141 = n68250 ^ n68251;
  assign n68247 = n68250 & n68251;
  assign n68261 = ~n68250;
  assign n68217 = ~n68275;
  assign n68270 = n68279 & n66016;
  assign n68283 = n68303 ^ n68304;
  assign n68264 = ~n68312;
  assign n68297 = n68313 & n1201;
  assign n68290 = ~n68303;
  assign n68245 = ~n68324;
  assign n68318 = n68329 & n68212;
  assign n68322 = n64410 & n67041;
  assign n68319 = n64410 & n66766;
  assign n67008 = ~n68331;
  assign n68316 = n68334 & n68335;
  assign n68330 = n68351 & n68352;
  assign n68071 = ~n68234;
  assign n68223 = n68235 & n13593;
  assign n68116 = ~n68247;
  assign n68243 = n68261 & n68262;
  assign n68254 = ~n68270;
  assign n68259 = n305 ^ n68283;
  assign n68289 = ~n68297;
  assign n68292 = n68316 ^ n68315;
  assign n68210 = ~n68318;
  assign n68301 = ~n68319;
  assign n68311 = n68316 & n68320;
  assign n67043 = ~n68322;
  assign n68306 = n68330 ^ n65215;
  assign n68314 = ~n68316;
  assign n68325 = ~n68330;
  assign n68103 = ~n68223;
  assign n68145 = ~n68243;
  assign n68242 = n68254 & n68220;
  assign n68170 = n68258 ^ n68259;
  assign n68219 = n68254 & n68217;
  assign n68183 = n68259 & n68267;
  assign n68278 = n68289 & n68290;
  assign n68237 = n68291 ^ n68292;
  assign n68162 = n68301 & n68302;
  assign n64340 = n68305 ^ n68306;
  assign n68295 = ~n68311;
  assign n68298 = n68314 & n68315;
  assign n68321 = n68325 & n68326;
  assign n64106 = n68219 ^ n68220;
  assign n68218 = n68170 & n65966;
  assign n68216 = ~n68242;
  assign n68222 = ~n68170;
  assign n68180 = ~n68183;
  assign n68266 = n68237 & n304;
  assign n68265 = ~n68237;
  assign n68263 = ~n68278;
  assign n68274 = n64340 & n66929;
  assign n68280 = n64340 & n65282;
  assign n68165 = ~n68162;
  assign n64370 = ~n64340;
  assign n68293 = n68295 & n68296;
  assign n68272 = ~n68298;
  assign n68307 = ~n68321;
  assign n68202 = n64106 & n65997;
  assign n64109 = ~n64106;
  assign n68199 = n68216 & n68217;
  assign n68174 = ~n68218;
  assign n68214 = n68222 & n65915;
  assign n68236 = n68263 & n68264;
  assign n68248 = n68265 & n1168;
  assign n68204 = ~n68266;
  assign n66932 = ~n68274;
  assign n68252 = ~n68280;
  assign n68268 = n64370 & n66681;
  assign n68273 = n64370 & n68288;
  assign n68271 = ~n68293;
  assign n68281 = n68307 & n68308;
  assign n68171 = n68199 ^ n65915;
  assign n68188 = n64109 & n67080;
  assign n68176 = ~n68202;
  assign n68195 = ~n68199;
  assign n68194 = ~n68214;
  assign n68205 = n68236 ^ n68237;
  assign n68239 = ~n68248;
  assign n68238 = ~n68236;
  assign n68253 = ~n68268;
  assign n68240 = n68271 & n68272;
  assign n66967 = ~n68273;
  assign n68260 = n68281 ^ n68282;
  assign n68284 = ~n68281;
  assign n64051 = n68170 ^ n68171;
  assign n68175 = ~n68188;
  assign n68186 = n68194 & n68195;
  assign n68184 = n304 ^ n68205;
  assign n68225 = n68238 & n68239;
  assign n68211 = n68240 ^ n68241;
  assign n68079 = n68252 & n68253;
  assign n64296 = n68260 ^ n65136;
  assign n68244 = ~n68240;
  assign n68255 = ~n68260;
  assign n68269 = n68284 & n68285;
  assign n68149 = n64051 & n65966;
  assign n64082 = ~n64051;
  assign n68140 = n68175 & n68176;
  assign n68106 = n68183 ^ n68184;
  assign n68173 = ~n68186;
  assign n68179 = ~n68184;
  assign n68182 = n68211 ^ n68212;
  assign n68203 = ~n68225;
  assign n68228 = n64296 & n68232;
  assign n68221 = n68079 & n68233;
  assign n68229 = n64296 & n66743;
  assign n64320 = ~n64296;
  assign n68231 = n68244 & n68245;
  assign n68224 = ~n68079;
  assign n68246 = n68255 & n65207;
  assign n68256 = ~n68269;
  assign n68105 = n68140 ^ n68141;
  assign n68134 = n64082 & n67010;
  assign n68120 = ~n68149;
  assign n68153 = n68106 & n65835;
  assign n68144 = ~n68140;
  assign n68154 = ~n68106;
  assign n68137 = n68173 & n68174;
  assign n68125 = n68179 & n68180;
  assign n68193 = n68182 & n319;
  assign n68181 = n68203 & n68204;
  assign n68189 = ~n68182;
  assign n68119 = ~n68221;
  assign n68215 = n64320 & n66896;
  assign n68213 = n68224 & n68111;
  assign n66891 = ~n68228;
  assign n68206 = ~n68229;
  assign n68209 = ~n68231;
  assign n68207 = ~n68246;
  assign n68230 = n68256 & n68257;
  assign n68081 = n68104 ^ n68105;
  assign n68102 = ~n68105;
  assign n68121 = ~n68134;
  assign n68107 = n68137 ^ n65835;
  assign n68133 = n68144 & n68145;
  assign n68089 = ~n68153;
  assign n68148 = n68154 & n65892;
  assign n68122 = ~n68137;
  assign n68136 = ~n68125;
  assign n68152 = n68181 ^ n68182;
  assign n68177 = n68189 & n1118;
  assign n68131 = ~n68193;
  assign n68157 = ~n68181;
  assign n68007 = n68206 & n68207;
  assign n68190 = n68209 & n68210;
  assign n68077 = ~n68213;
  assign n66856 = ~n68215;
  assign n68198 = n68230 ^ n65084;
  assign n68226 = ~n68230;
  assign n68053 = n326 ^ n68081;
  assign n68100 = n68102 & n68103;
  assign n64018 = n68106 ^ n68107;
  assign n68040 = n68120 & n68121;
  assign n68115 = ~n68133;
  assign n68123 = ~n68148;
  assign n68126 = n319 ^ n68152;
  assign n68156 = ~n68177;
  assign n68163 = n68190 ^ n68191;
  assign n68015 = ~n68007;
  assign n68187 = n68190 & n68196;
  assign n64253 = n68197 ^ n68198;
  assign n68192 = ~n68190;
  assign n68208 = n68226 & n68227;
  assign n66064 = n68053 ^ n66116;
  assign n68034 = ~n68053;
  assign n68084 = n64018 & n66901;
  assign n64041 = ~n64018;
  assign n68056 = ~n68040;
  assign n68070 = ~n68100;
  assign n68067 = n68115 & n68116;
  assign n68108 = n68122 & n68123;
  assign n68061 = n68125 ^ n68126;
  assign n68028 = n68126 & n68136;
  assign n68155 = n68156 & n68157;
  assign n68098 = n68162 ^ n68163;
  assign n68172 = n64253 & n66658;
  assign n68166 = n64253 & n68185;
  assign n68164 = ~n68187;
  assign n64287 = ~n64253;
  assign n68178 = n68192 & n68191;
  assign n68200 = ~n68208;
  assign n67347 = ~n66064;
  assign n67948 = n68034 & n66116;
  assign n68041 = n68067 ^ n68068;
  assign n67999 = n68070 & n68071;
  assign n68044 = ~n68084;
  assign n68065 = n64041 & n65835;
  assign n68069 = n68067 & n68068;
  assign n68082 = ~n68067;
  assign n68090 = n68061 & n65799;
  assign n68091 = ~n68061;
  assign n68088 = ~n68108;
  assign n68135 = n68098 & n318;
  assign n68132 = ~n68098;
  assign n68130 = ~n68155;
  assign n68159 = n68164 & n68165;
  assign n66817 = ~n68166;
  assign n68158 = n64287 & n66772;
  assign n68150 = ~n68172;
  assign n68161 = n64287 & n65084;
  assign n68143 = ~n68178;
  assign n68167 = n68200 & n68201;
  assign n68000 = n68040 ^ n68041;
  assign n68043 = n67999 & n13543;
  assign n68051 = ~n67999;
  assign n68045 = ~n68065;
  assign n68057 = ~n68069;
  assign n68066 = n68082 & n68083;
  assign n68060 = n68088 & n68089;
  assign n68021 = ~n68090;
  assign n68078 = n68091 & n65771;
  assign n68097 = n68130 & n68131;
  assign n68129 = n68132 & n1025;
  assign n68063 = ~n68135;
  assign n66775 = ~n68158;
  assign n68142 = ~n68159;
  assign n68151 = ~n68161;
  assign n68147 = n68167 ^ n65009;
  assign n68168 = ~n68167;
  assign n67972 = n67999 ^ n68000;
  assign n68010 = ~n68000;
  assign n68011 = ~n68043;
  assign n67960 = n68044 & n68045;
  assign n68025 = n68051 & n325;
  assign n68050 = n68056 & n68057;
  assign n68016 = n68060 ^ n68061;
  assign n68024 = ~n68066;
  assign n68055 = ~n68060;
  assign n68054 = ~n68078;
  assign n68064 = n68097 ^ n68098;
  assign n68096 = ~n68097;
  assign n68095 = ~n68129;
  assign n68110 = n68142 & n68143;
  assign n64212 = n68146 ^ n68147;
  assign n67933 = n68150 & n68151;
  assign n68160 = n68168 & n68169;
  assign n67949 = n325 ^ n67972;
  assign n67992 = n68010 & n68011;
  assign n68009 = n67960 & n67991;
  assign n63982 = n65771 ^ n68016;
  assign n68012 = ~n67960;
  assign n67977 = ~n68025;
  assign n68017 = n68016 & n65799;
  assign n68023 = ~n68050;
  assign n68047 = n68054 & n68055;
  assign n68029 = n318 ^ n68064;
  assign n68085 = n68095 & n68096;
  assign n68080 = n68110 ^ n68111;
  assign n68112 = n64212 & n68124;
  assign n68117 = n64212 & n65024;
  assign n68113 = n67933 & n68127;
  assign n68101 = ~n67933;
  assign n64247 = ~n64212;
  assign n68118 = ~n68110;
  assign n68138 = ~n68160;
  assign n65970 = n67948 ^ n67949;
  assign n67870 = n67949 & n67948;
  assign n67976 = ~n67992;
  assign n64005 = ~n63982;
  assign n67987 = ~n68009;
  assign n67997 = n68012 & n68013;
  assign n67953 = ~n68017;
  assign n67990 = n68023 & n68024;
  assign n67951 = n68028 ^ n68029;
  assign n67968 = n68029 & n68028;
  assign n68020 = ~n68047;
  assign n68032 = n68079 ^ n68080;
  assign n68062 = ~n68085;
  assign n68092 = n68101 & n67963;
  assign n68099 = n64247 & n66571;
  assign n66695 = ~n68112;
  assign n68093 = n64247 & n66691;
  assign n67955 = ~n68113;
  assign n68075 = ~n68117;
  assign n68094 = n68118 & n68119;
  assign n68114 = n68138 & n68139;
  assign n67310 = ~n65970;
  assign n67931 = n67976 & n67977;
  assign n67980 = n64005 & n66796;
  assign n67961 = n67990 ^ n67991;
  assign n67959 = ~n67997;
  assign n67988 = ~n67990;
  assign n67993 = n67951 & n65681;
  assign n67996 = ~n67951;
  assign n67998 = n68020 & n68021;
  assign n67966 = ~n67968;
  assign n68046 = n68032 & n317;
  assign n68031 = n68062 & n68063;
  assign n68048 = ~n68032;
  assign n67927 = ~n68092;
  assign n66733 = ~n68093;
  assign n68076 = ~n68094;
  assign n68074 = ~n68099;
  assign n68073 = n68114 ^ n64928;
  assign n68109 = n68114 & n68128;
  assign n67932 = n67960 ^ n67961;
  assign n67916 = ~n67931;
  assign n67952 = ~n67980;
  assign n67979 = n67987 & n67988;
  assign n67970 = ~n67993;
  assign n67989 = n67996 & n65701;
  assign n67971 = ~n67998;
  assign n67995 = n68031 ^ n68032;
  assign n67974 = ~n68046;
  assign n68026 = n68048 & n970;
  assign n68006 = ~n68031;
  assign n64166 = n68072 ^ n68073;
  assign n67867 = n68074 & n68075;
  assign n68035 = n68076 & n68077;
  assign n68086 = ~n68109;
  assign n67909 = n67931 ^ n67932;
  assign n67928 = n67932 & n13481;
  assign n67935 = ~n67932;
  assign n67907 = n67952 & n67953;
  assign n67967 = n67970 & n67971;
  assign n67950 = n67971 ^ n65701;
  assign n67958 = ~n67979;
  assign n67947 = ~n67989;
  assign n67969 = n317 ^ n67995;
  assign n68005 = ~n68026;
  assign n68008 = n68035 ^ n68036;
  assign n68039 = n64166 & n66610;
  assign n68042 = n64166 & n66499;
  assign n68049 = n68035 & n68036;
  assign n64168 = ~n64166;
  assign n67880 = ~n67867;
  assign n68037 = ~n68035;
  assign n68058 = n68086 & n68087;
  assign n67871 = n324 ^ n67909;
  assign n67915 = ~n67928;
  assign n67921 = n67935 & n324;
  assign n67911 = ~n67907;
  assign n63934 = n67950 ^ n67951;
  assign n67936 = n67958 & n67959;
  assign n67946 = ~n67967;
  assign n67887 = n67968 ^ n67969;
  assign n67965 = ~n67969;
  assign n67994 = n68005 & n68006;
  assign n67942 = n68007 ^ n68008;
  assign n68033 = n68037 & n68038;
  assign n66661 = ~n68039;
  assign n68001 = ~n68042;
  assign n68030 = n64168 & n64942;
  assign n68014 = ~n68049;
  assign n68027 = n64168 & n68052;
  assign n64171 = n68058 ^ n68059;
  assign n65938 = n67870 ^ n67871;
  assign n67798 = n67871 & n67870;
  assign n67901 = n67915 & n67916;
  assign n67884 = ~n67921;
  assign n67923 = n63934 & n66762;
  assign n67908 = n67936 ^ n67937;
  assign n63959 = ~n63934;
  assign n67924 = n67936 & n67937;
  assign n67929 = ~n67936;
  assign n67920 = n67946 & n67947;
  assign n67938 = n67887 & n65619;
  assign n67940 = ~n67887;
  assign n67895 = n67965 & n67966;
  assign n67978 = n67942 & n901;
  assign n67973 = ~n67994;
  assign n67975 = ~n67942;
  assign n68003 = n68014 & n68015;
  assign n67982 = n68022 ^ n64171;
  assign n66614 = ~n68027;
  assign n68002 = ~n68030;
  assign n68018 = n64171 & n66460;
  assign n67986 = ~n68033;
  assign n68019 = ~n64171;
  assign n67265 = ~n65938;
  assign n67790 = ~n67798;
  assign n67883 = ~n67901;
  assign n67857 = n67907 ^ n67908;
  assign n67912 = n63959 & n65701;
  assign n67888 = n67920 ^ n65586;
  assign n67886 = ~n67923;
  assign n67910 = ~n67924;
  assign n67922 = n67929 & n67930;
  assign n67913 = ~n67920;
  assign n67878 = ~n67938;
  assign n67925 = n67940 & n65586;
  assign n67893 = ~n67895;
  assign n67941 = n67973 & n67974;
  assign n67964 = n67975 & n316;
  assign n67944 = ~n67978;
  assign n66580 = n67981 ^ n67982;
  assign n67801 = n68001 & n68002;
  assign n67985 = ~n68003;
  assign n67983 = ~n68018;
  assign n68004 = n68019 & n64875;
  assign n67856 = n67883 & n67884;
  assign n67874 = n67857 & n13439;
  assign n63899 = n67887 ^ n67888;
  assign n67875 = ~n67857;
  assign n67903 = n67910 & n67911;
  assign n67885 = ~n67912;
  assign n67882 = ~n67922;
  assign n67914 = ~n67925;
  assign n67917 = n67941 ^ n67942;
  assign n67919 = ~n67964;
  assign n67943 = ~n67941;
  assign n67962 = n67985 & n67986;
  assign n67805 = ~n67801;
  assign n67984 = ~n68004;
  assign n67822 = n67856 ^ n67857;
  assign n67848 = ~n67874;
  assign n67866 = n67875 & n323;
  assign n67849 = ~n67856;
  assign n67865 = n63899 & n65619;
  assign n63935 = ~n63899;
  assign n67817 = n67885 & n67886;
  assign n67881 = ~n67903;
  assign n67902 = n67913 & n67914;
  assign n67896 = n316 ^ n67917;
  assign n67939 = n67943 & n67944;
  assign n67934 = n67962 ^ n67963;
  assign n67954 = ~n67962;
  assign n67956 = n67983 & n67984;
  assign n67799 = n323 ^ n67822;
  assign n67846 = n67848 & n67849;
  assign n67853 = n63935 & n66648;
  assign n67831 = ~n67865;
  assign n67824 = ~n67866;
  assign n67860 = n67817 & n67876;
  assign n67864 = ~n67817;
  assign n67851 = n67881 & n67882;
  assign n67820 = n67895 ^ n67896;
  assign n67877 = ~n67902;
  assign n67892 = ~n67896;
  assign n67891 = n67933 ^ n67934;
  assign n67918 = ~n67939;
  assign n67945 = n67954 & n67955;
  assign n67726 = n67956 ^ n67957;
  assign n65821 = n67798 ^ n67799;
  assign n67789 = ~n67799;
  assign n67823 = ~n67846;
  assign n67818 = n67851 ^ n67852;
  assign n67830 = ~n67853;
  assign n67845 = ~n67860;
  assign n67850 = n67864 & n67852;
  assign n67844 = ~n67851;
  assign n67862 = n67820 & n65555;
  assign n67847 = n67877 & n67878;
  assign n67861 = ~n67820;
  assign n67833 = n67892 & n67893;
  assign n67897 = n67891 & n315;
  assign n67890 = n67918 & n67919;
  assign n67900 = ~n67891;
  assign n67926 = ~n67945;
  assign n67215 = ~n65821;
  assign n67740 = n67789 & n67790;
  assign n67794 = n67817 ^ n67818;
  assign n67793 = n67823 & n67824;
  assign n67758 = n67830 & n67831;
  assign n67828 = n67844 & n67845;
  assign n67821 = n67847 ^ n65502;
  assign n67810 = ~n67850;
  assign n67858 = n67861 & n65502;
  assign n67838 = ~n67862;
  assign n67839 = ~n67847;
  assign n67837 = ~n67833;
  assign n67863 = n67890 ^ n67891;
  assign n67842 = ~n67897;
  assign n67894 = n67900 & n840;
  assign n67873 = ~n67890;
  assign n67904 = n67926 & n67927;
  assign n67766 = n67793 ^ n67794;
  assign n67792 = n67794 & n322;
  assign n67771 = ~n67793;
  assign n67797 = ~n67794;
  assign n63868 = n67820 ^ n67821;
  assign n67765 = ~n67758;
  assign n67809 = ~n67828;
  assign n67835 = n67838 & n67839;
  assign n67814 = ~n67858;
  assign n67834 = n315 ^ n67863;
  assign n67872 = ~n67894;
  assign n67868 = n67904 ^ n67905;
  assign n67906 = n67904 & n67905;
  assign n67898 = ~n67904;
  assign n67741 = n322 ^ n67766;
  assign n67749 = ~n67792;
  assign n67780 = n67797 & n13411;
  assign n67791 = n63868 & n65502;
  assign n67781 = n67809 & n67810;
  assign n63891 = ~n63868;
  assign n67762 = n67833 ^ n67834;
  assign n67813 = ~n67835;
  assign n67836 = ~n67834;
  assign n67816 = n67867 ^ n67868;
  assign n67859 = n67872 & n67873;
  assign n67889 = n67898 & n67899;
  assign n67879 = ~n67906;
  assign n65746 = n67740 ^ n67741;
  assign n67681 = n67741 & n67740;
  assign n67770 = ~n67780;
  assign n67759 = n67781 ^ n67782;
  assign n67773 = ~n67791;
  assign n67779 = n67781 & n67796;
  assign n67784 = n63891 & n66594;
  assign n67783 = ~n67781;
  assign n67788 = n67813 & n67814;
  assign n67803 = n67762 & n65408;
  assign n67807 = ~n67762;
  assign n67760 = n67836 & n67837;
  assign n67840 = n67816 & n792;
  assign n67841 = ~n67859;
  assign n67843 = ~n67816;
  assign n67869 = n67879 & n67880;
  assign n67855 = ~n67889;
  assign n67154 = ~n65746;
  assign n67684 = ~n67681;
  assign n67718 = n67758 ^ n67759;
  assign n67754 = n67770 & n67771;
  assign n67764 = ~n67779;
  assign n67778 = n67783 & n67782;
  assign n67772 = ~n67784;
  assign n67763 = n67788 ^ n65408;
  assign n67752 = ~n67803;
  assign n67776 = ~n67788;
  assign n67800 = n67807 & n65454;
  assign n67811 = ~n67840;
  assign n67815 = n67841 & n67842;
  assign n67829 = n67843 & n314;
  assign n67854 = ~n67869;
  assign n67736 = n67718 & n321;
  assign n67737 = ~n67718;
  assign n67748 = ~n67754;
  assign n63828 = n67762 ^ n67763;
  assign n67753 = n67764 & n67765;
  assign n67701 = n67772 & n67773;
  assign n67743 = ~n67778;
  assign n67777 = ~n67800;
  assign n67785 = n67815 ^ n67816;
  assign n67812 = ~n67815;
  assign n67787 = ~n67829;
  assign n67827 = n67854 & n67855;
  assign n67694 = ~n67736;
  assign n67727 = n67737 & n13365;
  assign n67732 = n63828 & n66492;
  assign n67717 = n67748 & n67749;
  assign n67745 = n67701 & n67720;
  assign n63831 = ~n63828;
  assign n67742 = ~n67753;
  assign n67746 = ~n67701;
  assign n67768 = n67776 & n67777;
  assign n67761 = n314 ^ n67785;
  assign n67806 = n67811 & n67812;
  assign n67802 = n67827 ^ n67826;
  assign n67819 = n67827 & n67832;
  assign n67825 = ~n67827;
  assign n67698 = n67717 ^ n67718;
  assign n67716 = ~n67727;
  assign n67729 = n63831 & n65408;
  assign n67710 = ~n67732;
  assign n67715 = ~n67717;
  assign n67719 = n67742 & n67743;
  assign n67724 = ~n67745;
  assign n67734 = n67746 & n67747;
  assign n67700 = n67760 ^ n67761;
  assign n67751 = ~n67768;
  assign n67709 = n67761 & n67760;
  assign n67757 = n67801 ^ n67802;
  assign n67786 = ~n67806;
  assign n67804 = ~n67819;
  assign n67808 = n67825 & n67826;
  assign n67682 = n321 ^ n67698;
  assign n67705 = n67715 & n67716;
  assign n67702 = n67719 ^ n67720;
  assign n67711 = ~n67729;
  assign n67704 = ~n67734;
  assign n67723 = ~n67719;
  assign n67733 = n67700 & n65328;
  assign n67730 = ~n67700;
  assign n67744 = n67751 & n67752;
  assign n67767 = n67757 & n313;
  assign n67769 = ~n67757;
  assign n67756 = n67786 & n67787;
  assign n67795 = n67804 & n67805;
  assign n67775 = ~n67808;
  assign n65674 = n67681 ^ n67682;
  assign n67683 = ~n67682;
  assign n67670 = n67701 ^ n67702;
  assign n67693 = ~n67705;
  assign n67656 = n67710 & n67711;
  assign n67707 = n67723 & n67724;
  assign n67728 = n67730 & n65373;
  assign n67692 = ~n67733;
  assign n67713 = ~n67744;
  assign n67735 = n67756 ^ n67757;
  assign n67722 = ~n67767;
  assign n67755 = n67769 & n746;
  assign n67739 = ~n67756;
  assign n67774 = ~n67795;
  assign n67106 = ~n65674;
  assign n67637 = n67683 & n67684;
  assign n67679 = n67670 & n13319;
  assign n67669 = n67693 & n67694;
  assign n67675 = ~n67670;
  assign n67664 = ~n67656;
  assign n67703 = ~n67707;
  assign n67699 = n67713 ^ n65373;
  assign n67714 = ~n67728;
  assign n67712 = n313 ^ n67735;
  assign n67738 = ~n67755;
  assign n67750 = n67774 & n67775;
  assign n67650 = n67669 ^ n67670;
  assign n67634 = ~n67637;
  assign n67668 = n67675 & n320;
  assign n67665 = ~n67679;
  assign n67666 = ~n67669;
  assign n63772 = n67699 ^ n67700;
  assign n67680 = n67703 & n67704;
  assign n67648 = n67709 ^ n67712;
  assign n67706 = n67713 & n67714;
  assign n67708 = ~n67712;
  assign n67731 = n67738 & n67739;
  assign n67725 = n312 ^ n67750;
  assign n67638 = n320 ^ n67650;
  assign n67660 = n67665 & n67666;
  assign n67647 = ~n67668;
  assign n67657 = n67680 ^ n67678;
  assign n67687 = n67680 & n67688;
  assign n67676 = n63772 & n66440;
  assign n67677 = ~n67680;
  assign n63795 = ~n63772;
  assign n67690 = n67648 & n65240;
  assign n67695 = ~n67648;
  assign n67691 = ~n67706;
  assign n67685 = n67708 & n67709;
  assign n67697 = n67725 ^ n67726;
  assign n67721 = ~n67731;
  assign n65583 = n67637 ^ n67638;
  assign n67633 = ~n67638;
  assign n67623 = n67656 ^ n67657;
  assign n67646 = ~n67660;
  assign n67655 = ~n67676;
  assign n67671 = n67677 & n67678;
  assign n67672 = n63795 & n65328;
  assign n67663 = ~n67687;
  assign n67674 = ~n67690;
  assign n67667 = n67691 & n67692;
  assign n67689 = n67695 & n65268;
  assign n67696 = n67721 & n67722;
  assign n67038 = ~n65583;
  assign n67596 = n67633 & n67634;
  assign n67642 = n67623 & n335;
  assign n67622 = n67646 & n67647;
  assign n67643 = ~n67623;
  assign n67659 = n67663 & n67664;
  assign n67649 = n67667 ^ n65240;
  assign n67645 = ~n67671;
  assign n67654 = ~n67672;
  assign n67673 = ~n67667;
  assign n67652 = ~n67689;
  assign n67686 = n67696 ^ n67697;
  assign n67608 = n67622 ^ n67623;
  assign n67620 = ~n67622;
  assign n67605 = ~n67642;
  assign n67629 = n67643 & n13293;
  assign n63734 = n67648 ^ n67649;
  assign n67606 = n67654 & n67655;
  assign n67644 = ~n67659;
  assign n67662 = n67673 & n67674;
  assign n67612 = n67685 ^ n67686;
  assign n67597 = n335 ^ n67608;
  assign n67619 = ~n67629;
  assign n67630 = n63734 & n66357;
  assign n67627 = n67644 & n67645;
  assign n63756 = ~n63734;
  assign n67641 = n67606 & n67628;
  assign n67639 = ~n67606;
  assign n67651 = ~n67662;
  assign n67661 = n67612 & n65162;
  assign n67658 = ~n67612;
  assign n65538 = n67596 ^ n67597;
  assign n67548 = n67597 & n67596;
  assign n67611 = n67619 & n67620;
  assign n67607 = n67627 ^ n67628;
  assign n67624 = n63756 & n65268;
  assign n67616 = ~n67630;
  assign n67631 = n67639 & n67640;
  assign n67625 = ~n67627;
  assign n67626 = ~n67641;
  assign n67632 = n67651 & n67652;
  assign n67653 = n67658 & n65183;
  assign n67636 = ~n67661;
  assign n66987 = ~n65538;
  assign n67586 = n67606 ^ n67607;
  assign n67604 = ~n67611;
  assign n67617 = ~n67624;
  assign n67618 = n67625 & n67626;
  assign n67610 = ~n67631;
  assign n67613 = n67632 ^ n65162;
  assign n67635 = ~n67632;
  assign n67615 = ~n67653;
  assign n67598 = n67586 & n13253;
  assign n67599 = ~n67586;
  assign n67585 = n67604 & n67605;
  assign n63672 = n67612 ^ n67613;
  assign n67573 = n67616 & n67617;
  assign n67609 = ~n67618;
  assign n67621 = n67635 & n67636;
  assign n67567 = n67585 ^ n67586;
  assign n67576 = ~n67598;
  assign n67587 = n67599 & n334;
  assign n67577 = ~n67585;
  assign n67601 = n63672 & n66308;
  assign n67582 = ~n67573;
  assign n63728 = ~n63672;
  assign n67594 = n67609 & n67610;
  assign n67614 = ~n67621;
  assign n67549 = n334 ^ n67567;
  assign n67575 = n67576 & n67577;
  assign n67565 = ~n67587;
  assign n67574 = n67594 ^ n67595;
  assign n67593 = n63728 & n65183;
  assign n67580 = ~n67601;
  assign n67589 = n67594 & n67595;
  assign n67590 = ~n67594;
  assign n67603 = n67614 & n67615;
  assign n65421 = n67548 ^ n67549;
  assign n67550 = ~n67549;
  assign n67542 = n67573 ^ n67574;
  assign n67564 = ~n67575;
  assign n67581 = ~n67589;
  assign n67588 = n67590 & n67591;
  assign n67579 = ~n67593;
  assign n67600 = n67603 & n65125;
  assign n67602 = ~n67603;
  assign n66909 = ~n65421;
  assign n67505 = n67550 & n67548;
  assign n67541 = n67564 & n67565;
  assign n67557 = n67542 & n13222;
  assign n67556 = ~n67542;
  assign n67524 = n67579 & n67580;
  assign n67571 = n67581 & n67582;
  assign n67563 = ~n67588;
  assign n67583 = ~n67600;
  assign n67592 = n67602 & n65061;
  assign n67530 = n67541 ^ n67542;
  assign n67518 = ~n67505;
  assign n67553 = n67556 & n333;
  assign n67547 = ~n67557;
  assign n67546 = ~n67541;
  assign n67566 = n67524 & n67568;
  assign n67561 = ~n67524;
  assign n67562 = ~n67571;
  assign n67578 = n67583 & n67584;
  assign n67570 = ~n67592;
  assign n67506 = n333 ^ n67530;
  assign n67538 = n67546 & n67547;
  assign n67527 = ~n67553;
  assign n67560 = n67561 & n67545;
  assign n67544 = n67562 & n67563;
  assign n67540 = ~n67566;
  assign n67569 = ~n67578;
  assign n67572 = n67570 & n67583;
  assign n65325 = n67505 ^ n67506;
  assign n67476 = n67506 & n67518;
  assign n67526 = ~n67538;
  assign n67525 = n67544 ^ n67545;
  assign n67539 = ~n67544;
  assign n67529 = ~n67560;
  assign n67551 = n67569 & n67570;
  assign n67558 = ~n67572;
  assign n66827 = ~n65325;
  assign n67487 = ~n67476;
  assign n67510 = n67524 ^ n67525;
  assign n67509 = n67526 & n67527;
  assign n67536 = n67539 & n67540;
  assign n67533 = n67551 ^ n67552;
  assign n63655 = n67558 ^ n67559;
  assign n67554 = ~n67551;
  assign n67493 = n67509 ^ n67510;
  assign n67517 = n67510 & n332;
  assign n67511 = ~n67510;
  assign n67490 = ~n67509;
  assign n63613 = n64979 ^ n67533;
  assign n67528 = ~n67536;
  assign n67531 = n67533 & n65013;
  assign n67537 = n63655 & n65061;
  assign n63690 = ~n63655;
  assign n67543 = n67554 & n67555;
  assign n67477 = n332 ^ n67493;
  assign n67503 = n67511 & n13196;
  assign n67474 = ~n67517;
  assign n63642 = ~n63613;
  assign n67513 = n67528 & n67529;
  assign n67496 = ~n67531;
  assign n67523 = ~n67537;
  assign n67532 = n63690 & n66225;
  assign n67534 = ~n67543;
  assign n65232 = n67476 ^ n67477;
  assign n67422 = n67477 & n67487;
  assign n67489 = ~n67503;
  assign n67492 = n67513 ^ n67514;
  assign n67507 = n63642 & n66209;
  assign n67512 = n67513 & n67514;
  assign n67515 = ~n67513;
  assign n67522 = ~n67532;
  assign n67521 = n67534 & n67535;
  assign n66734 = ~n65232;
  assign n67488 = n67489 & n67490;
  assign n67495 = ~n67507;
  assign n67499 = ~n67512;
  assign n67504 = n67515 & n67516;
  assign n67498 = n67521 ^ n64906;
  assign n67491 = n67522 & n67523;
  assign n67519 = ~n67521;
  assign n67473 = ~n67488;
  assign n67457 = n67491 ^ n67492;
  assign n67448 = n67495 & n67496;
  assign n63548 = n67497 ^ n67498;
  assign n67482 = ~n67504;
  assign n67508 = n67519 & n67520;
  assign n67500 = ~n67491;
  assign n67456 = n67473 & n67474;
  assign n67469 = n67457 & n13171;
  assign n67480 = n67448 & n67459;
  assign n67472 = ~n67457;
  assign n67478 = n63548 & n66152;
  assign n67485 = ~n67448;
  assign n63591 = ~n63548;
  assign n67494 = n67499 & n67500;
  assign n67501 = ~n67508;
  assign n67443 = n67456 ^ n67457;
  assign n67454 = ~n67456;
  assign n67455 = ~n67469;
  assign n67468 = n67472 & n331;
  assign n67462 = ~n67478;
  assign n67471 = n63591 & n64906;
  assign n67465 = ~n67480;
  assign n67470 = n67485 & n67486;
  assign n67481 = ~n67494;
  assign n67479 = n67501 & n67502;
  assign n67425 = n331 ^ n67443;
  assign n67452 = n67454 & n67455;
  assign n67440 = ~n67468;
  assign n67451 = ~n67470;
  assign n67463 = ~n67471;
  assign n67467 = n67479 ^ n64851;
  assign n67458 = n67481 & n67482;
  assign n67483 = ~n67479;
  assign n65146 = n67422 ^ n67425;
  assign n67421 = ~n67425;
  assign n67439 = ~n67452;
  assign n67449 = n67458 ^ n67459;
  assign n67411 = n67462 & n67463;
  assign n63530 = n67466 ^ n67467;
  assign n67464 = ~n67458;
  assign n67475 = n67483 & n67484;
  assign n66653 = ~n65146;
  assign n67384 = n67421 & n67422;
  assign n67423 = n67439 & n67440;
  assign n67424 = n67448 ^ n67449;
  assign n67444 = n63530 & n66112;
  assign n67415 = ~n67411;
  assign n63556 = ~n63530;
  assign n67453 = n67464 & n67465;
  assign n67460 = ~n67475;
  assign n67391 = ~n67384;
  assign n67402 = n67423 ^ n67424;
  assign n67437 = n67424 & n13098;
  assign n67417 = ~n67423;
  assign n67427 = ~n67424;
  assign n67434 = ~n67444;
  assign n67441 = n63556 & n64851;
  assign n67450 = ~n67453;
  assign n67445 = n67460 & n67461;
  assign n67385 = n330 ^ n67402;
  assign n67419 = n67427 & n330;
  assign n67416 = ~n67437;
  assign n67433 = ~n67441;
  assign n67431 = n67445 ^ n64755;
  assign n67432 = n67450 & n67451;
  assign n67446 = ~n67445;
  assign n65071 = n67384 ^ n67385;
  assign n67340 = n67385 & n67391;
  assign n67403 = n67416 & n67417;
  assign n67396 = ~n67419;
  assign n63479 = n67430 ^ n67431;
  assign n67412 = n67432 ^ n67429;
  assign n67362 = n67433 & n67434;
  assign n67426 = n67432 & n67438;
  assign n67428 = ~n67432;
  assign n67442 = n67446 & n67447;
  assign n66581 = ~n65071;
  assign n67349 = ~n67340;
  assign n67395 = ~n67403;
  assign n67380 = n67411 ^ n67412;
  assign n67404 = n63479 & n64755;
  assign n67410 = n67362 & n67418;
  assign n63523 = ~n63479;
  assign n67413 = ~n67362;
  assign n67414 = ~n67426;
  assign n67420 = n67428 & n67429;
  assign n67435 = ~n67442;
  assign n67379 = n67395 & n67396;
  assign n67387 = n67380 & n329;
  assign n67386 = ~n67380;
  assign n67400 = n63523 & n66069;
  assign n67390 = ~n67404;
  assign n67377 = ~n67410;
  assign n67399 = n67413 & n67382;
  assign n67409 = n67414 & n67415;
  assign n67398 = ~n67420;
  assign n67405 = n67435 & n67436;
  assign n67364 = n67379 ^ n67380;
  assign n67370 = ~n67379;
  assign n67383 = n67386 & n13075;
  assign n67357 = ~n67387;
  assign n67361 = ~n67399;
  assign n67389 = ~n67400;
  assign n67388 = n67405 ^ n67406;
  assign n67397 = ~n67409;
  assign n67407 = ~n67405;
  assign n67341 = n329 ^ n67364;
  assign n67371 = ~n67383;
  assign n63447 = n64707 ^ n67388;
  assign n67309 = n67389 & n67390;
  assign n67392 = n67388 & n64745;
  assign n67381 = n67397 & n67398;
  assign n67401 = n67407 & n67408;
  assign n64992 = n67340 ^ n67341;
  assign n67300 = n67341 & n67349;
  assign n67366 = n67370 & n67371;
  assign n67369 = n63447 & n67378;
  assign n67363 = n67381 ^ n67382;
  assign n63484 = ~n63447;
  assign n67376 = ~n67381;
  assign n67359 = ~n67392;
  assign n67393 = ~n67401;
  assign n67299 = ~n67300;
  assign n67330 = n67362 ^ n67363;
  assign n67356 = ~n67366;
  assign n66089 = ~n67369;
  assign n67368 = n63484 & n66116;
  assign n67365 = n63484 & n66006;
  assign n67372 = n67376 & n67377;
  assign n67373 = n67393 & n67394;
  assign n67344 = n67330 & n328;
  assign n67342 = ~n67330;
  assign n67329 = n67356 & n67357;
  assign n67358 = ~n67365;
  assign n66118 = ~n67368;
  assign n67360 = ~n67372;
  assign n67353 = n67373 ^ n64689;
  assign n67374 = ~n67373;
  assign n67313 = n67329 ^ n67330;
  assign n67339 = n67342 & n13017;
  assign n67307 = ~n67344;
  assign n67324 = ~n67329;
  assign n63398 = n67352 ^ n67353;
  assign n67289 = n67358 & n67359;
  assign n67350 = n67360 & n67361;
  assign n67367 = n67374 & n67375;
  assign n67301 = n328 ^ n67313;
  assign n67323 = ~n67339;
  assign n67332 = n63398 & n67347;
  assign n67336 = n67289 & n67348;
  assign n67333 = n63398 & n64689;
  assign n67343 = n67350 & n67351;
  assign n67338 = ~n67289;
  assign n63442 = ~n63398;
  assign n67345 = ~n67350;
  assign n67354 = ~n67367;
  assign n67272 = n67300 ^ n67301;
  assign n67298 = ~n67301;
  assign n67318 = n67323 & n67324;
  assign n67325 = n63442 & n66064;
  assign n66034 = ~n67332;
  assign n67315 = ~n67333;
  assign n67287 = ~n67336;
  assign n67328 = n67338 & n67271;
  assign n67327 = n63442 & n65935;
  assign n67322 = ~n67343;
  assign n67331 = n67345 & n67346;
  assign n67337 = n67354 & n67355;
  assign n63131 = n67272 ^ n64198;
  assign n67165 = n67272 & n64200;
  assign n67278 = ~n67272;
  assign n67236 = n67298 & n67299;
  assign n67306 = ~n67318;
  assign n66059 = ~n67325;
  assign n67314 = ~n67327;
  assign n67321 = n67322 & n67309;
  assign n67268 = ~n67328;
  assign n67312 = ~n67331;
  assign n67320 = n67337 ^ n64634;
  assign n67334 = ~n67337;
  assign n67260 = n63131 & n66125;
  assign n63113 = ~n63131;
  assign n67269 = n67278 & n64200;
  assign n67247 = ~n67236;
  assign n67281 = n67306 & n67307;
  assign n67223 = n67314 & n67315;
  assign n63369 = n67319 ^ n67320;
  assign n67311 = ~n67321;
  assign n67308 = n67312 & n67322;
  assign n67326 = n67334 & n67335;
  assign n67234 = ~n67260;
  assign n67235 = ~n67269;
  assign n67263 = ~n67281;
  assign n67294 = n67223 & n67305;
  assign n67297 = n63369 & n65839;
  assign n67282 = n67308 ^ n67309;
  assign n67296 = n63369 & n67310;
  assign n67304 = ~n67223;
  assign n63384 = ~n63369;
  assign n67288 = n67311 & n67312;
  assign n67316 = ~n67326;
  assign n67219 = n67234 & n67235;
  assign n67266 = n67281 ^ n67282;
  assign n67270 = n67288 ^ n67289;
  assign n67283 = n67282 & n343;
  assign n67244 = ~n67294;
  assign n67285 = ~n67282;
  assign n66001 = ~n67296;
  assign n67280 = ~n67297;
  assign n67291 = n63384 & n65970;
  assign n67290 = n67304 & n67249;
  assign n67293 = n63384 & n64653;
  assign n67286 = ~n67288;
  assign n67295 = n67316 & n67317;
  assign n67190 = n67219 ^ n67220;
  assign n67221 = ~n67219;
  assign n67237 = n343 ^ n67266;
  assign n67214 = n67270 ^ n67271;
  assign n67239 = ~n67283;
  assign n67275 = n67285 & n12996;
  assign n67284 = n67286 & n67287;
  assign n67226 = ~n67290;
  assign n65974 = ~n67291;
  assign n67279 = ~n67293;
  assign n67277 = n67295 ^ n64596;
  assign n67302 = ~n67295;
  assign n64586 = n359 ^ n67190;
  assign n66907 = n67190 & n359;
  assign n67022 = n67221 & n67222;
  assign n67227 = n67236 ^ n67237;
  assign n67168 = n67237 & n67247;
  assign n67246 = n67214 & n342;
  assign n67251 = ~n67214;
  assign n67262 = ~n67275;
  assign n63321 = n67276 ^ n67277;
  assign n67174 = n67279 & n67280;
  assign n67267 = ~n67284;
  assign n67292 = n67302 & n67303;
  assign n65737 = ~n64586;
  assign n67218 = n67227 & n64106;
  assign n67212 = ~n67227;
  assign n67186 = ~n67246;
  assign n67241 = n67251 & n12940;
  assign n67256 = n63321 & n65797;
  assign n67253 = n67262 & n67263;
  assign n67259 = n67174 & n67264;
  assign n67254 = n63321 & n67265;
  assign n67248 = n67267 & n67268;
  assign n63340 = ~n63321;
  assign n67255 = ~n67174;
  assign n67273 = ~n67292;
  assign n67202 = n67212 & n64109;
  assign n67171 = ~n67218;
  assign n67216 = ~n67241;
  assign n67224 = n67248 ^ n67249;
  assign n67238 = ~n67253;
  assign n65940 = ~n67254;
  assign n67242 = n67255 & n67200;
  assign n67228 = ~n67256;
  assign n67252 = n63340 & n65938;
  assign n67198 = ~n67259;
  assign n67245 = n63340 & n64596;
  assign n67243 = ~n67248;
  assign n67261 = n67273 & n67274;
  assign n67187 = ~n67202;
  assign n67167 = n67223 ^ n67224;
  assign n67213 = n67238 & n67239;
  assign n67177 = ~n67242;
  assign n67240 = n67243 & n67244;
  assign n67229 = ~n67245;
  assign n65907 = ~n67252;
  assign n67233 = n67261 ^ n64559;
  assign n67257 = ~n67261;
  assign n67184 = n67187 & n67165;
  assign n67164 = n67187 & n67171;
  assign n67193 = n67167 & n341;
  assign n67191 = n67213 ^ n67214;
  assign n67201 = ~n67167;
  assign n67125 = n67228 & n67229;
  assign n67217 = ~n67213;
  assign n63282 = n67232 ^ n67233;
  assign n67225 = ~n67240;
  assign n67250 = n67257 & n67258;
  assign n63020 = n67164 ^ n67165;
  assign n67170 = ~n67184;
  assign n67169 = n342 ^ n67191;
  assign n67136 = ~n67193;
  assign n67188 = n67201 & n12900;
  assign n67210 = n63282 & n67215;
  assign n67207 = n63282 & n64559;
  assign n67205 = n67125 & n67145;
  assign n67211 = n67216 & n67217;
  assign n67203 = ~n67125;
  assign n67199 = n67225 & n67226;
  assign n63316 = ~n63282;
  assign n67230 = ~n67250;
  assign n67143 = n63020 & n64106;
  assign n63022 = ~n63020;
  assign n67117 = n67168 ^ n67169;
  assign n67142 = n67170 & n67171;
  assign n67119 = n67169 & n67168;
  assign n67172 = ~n67188;
  assign n67175 = n67199 ^ n67200;
  assign n67195 = n63316 & n65644;
  assign n67192 = n67203 & n67204;
  assign n67194 = n63316 & n65821;
  assign n67152 = ~n67205;
  assign n67182 = ~n67207;
  assign n65830 = ~n67210;
  assign n67185 = ~n67211;
  assign n67197 = ~n67199;
  assign n67206 = n67230 & n67231;
  assign n67134 = n63022 & n65997;
  assign n67118 = n67142 ^ n64051;
  assign n67111 = ~n67143;
  assign n67138 = n67117 & n64082;
  assign n67122 = ~n67142;
  assign n67137 = ~n67117;
  assign n67114 = n67174 ^ n67175;
  assign n67166 = n67185 & n67186;
  assign n67124 = ~n67192;
  assign n65867 = ~n67194;
  assign n67183 = ~n67195;
  assign n67189 = n67197 & n67198;
  assign n67179 = n67206 ^ n64527;
  assign n67208 = ~n67206;
  assign n62915 = n67117 ^ n67118;
  assign n67110 = ~n67134;
  assign n67131 = n67137 & n64051;
  assign n67121 = ~n67138;
  assign n67153 = n67114 & n340;
  assign n67141 = n67166 ^ n67167;
  assign n67150 = ~n67114;
  assign n67173 = ~n67166;
  assign n63245 = n67178 ^ n67179;
  assign n67060 = n67182 & n67183;
  assign n67176 = ~n67189;
  assign n67196 = n67208 & n67209;
  assign n67085 = n62915 & n64051;
  assign n62957 = ~n62915;
  assign n67098 = n67110 & n67111;
  assign n67112 = n67121 & n67122;
  assign n67097 = ~n67131;
  assign n67120 = n341 ^ n67141;
  assign n67140 = n67150 & n12857;
  assign n67076 = ~n67153;
  assign n67162 = n67060 & n67163;
  assign n67161 = n63245 & n65746;
  assign n67155 = n67172 & n67173;
  assign n67159 = n63245 & n65601;
  assign n67160 = ~n67060;
  assign n63268 = ~n63245;
  assign n67144 = n67176 & n67177;
  assign n67180 = ~n67196;
  assign n67070 = n62957 & n65966;
  assign n67056 = ~n67085;
  assign n67084 = n67098 & n67099;
  assign n67079 = ~n67098;
  assign n67096 = ~n67112;
  assign n67017 = n67119 ^ n67120;
  assign n67051 = n67120 & n67119;
  assign n67116 = ~n67140;
  assign n67126 = n67144 ^ n67145;
  assign n67148 = n63268 & n67154;
  assign n67135 = ~n67155;
  assign n67146 = n63268 & n64527;
  assign n67130 = ~n67159;
  assign n67147 = n67160 & n67089;
  assign n65791 = ~n67161;
  assign n67094 = ~n67162;
  assign n67151 = ~n67144;
  assign n67156 = n67180 & n67181;
  assign n67055 = ~n67070;
  assign n67073 = n67079 & n67080;
  assign n67047 = ~n67084;
  assign n67074 = n67017 & n64018;
  assign n67083 = n67096 & n67097;
  assign n67082 = ~n67017;
  assign n67058 = n67125 ^ n67126;
  assign n67113 = n67135 & n67136;
  assign n67129 = ~n67146;
  assign n67063 = ~n67147;
  assign n65745 = ~n67148;
  assign n67139 = n67151 & n67152;
  assign n67133 = n67156 ^ n64471;
  assign n67157 = ~n67156;
  assign n66949 = n67055 & n67056;
  assign n67050 = n67047 & n67022;
  assign n67033 = ~n67073;
  assign n67064 = ~n67074;
  assign n67067 = n67082 & n64041;
  assign n67054 = ~n67083;
  assign n67095 = n67058 & n12818;
  assign n67078 = n67113 ^ n67114;
  assign n67087 = ~n67058;
  assign n66995 = n67129 & n67130;
  assign n67115 = ~n67113;
  assign n63194 = n67132 ^ n67133;
  assign n67123 = ~n67139;
  assign n67149 = n67157 & n67158;
  assign n67011 = n66949 & n67000;
  assign n67009 = ~n66949;
  assign n67021 = n67033 & n67047;
  assign n67032 = ~n67050;
  assign n67016 = n67054 ^ n64041;
  assign n67059 = n67064 & n67054;
  assign n67036 = ~n67067;
  assign n67052 = n340 ^ n67078;
  assign n67081 = n67087 & n339;
  assign n67049 = ~n67095;
  assign n67107 = n67115 & n67116;
  assign n67104 = n63194 & n64471;
  assign n67102 = n63194 & n65674;
  assign n67105 = n66995 & n67026;
  assign n67088 = n67123 & n67124;
  assign n67108 = ~n66995;
  assign n63231 = ~n63194;
  assign n67127 = ~n67149;
  assign n67003 = n67009 & n67010;
  assign n66992 = ~n67011;
  assign n62837 = n67016 ^ n67017;
  assign n66994 = n67021 ^ n67022;
  assign n66999 = n67032 & n67033;
  assign n66961 = n67051 ^ n67052;
  assign n67035 = ~n67059;
  assign n66976 = n67052 & n67051;
  assign n67020 = ~n67081;
  assign n67061 = n67088 ^ n67089;
  assign n65662 = ~n67102;
  assign n67072 = ~n67104;
  assign n67028 = ~n67105;
  assign n67086 = n63231 & n65473;
  assign n67091 = n63231 & n67106;
  assign n67075 = ~n67107;
  assign n67090 = n67108 & n67109;
  assign n67093 = ~n67088;
  assign n67103 = n67127 & n67128;
  assign n66982 = n62837 & n65835;
  assign n66977 = n66994 & n358;
  assign n66950 = n66999 ^ n67000;
  assign n66983 = ~n66994;
  assign n66960 = ~n67003;
  assign n62853 = ~n62837;
  assign n66993 = ~n66999;
  assign n67013 = n66961 & n64005;
  assign n66990 = n67035 & n67036;
  assign n67014 = ~n66961;
  assign n66980 = n67060 ^ n67061;
  assign n67057 = n67075 & n67076;
  assign n67071 = ~n67086;
  assign n66998 = ~n67090;
  assign n65707 = ~n67091;
  assign n67077 = n67093 & n67094;
  assign n67069 = n67103 ^ n64408;
  assign n67100 = ~n67103;
  assign n66861 = n66949 ^ n66950;
  assign n66903 = ~n66977;
  assign n66939 = ~n66982;
  assign n66970 = n66983 & n4928;
  assign n66965 = n62853 & n64041;
  assign n66962 = n66990 ^ n63982;
  assign n66981 = n66992 & n66993;
  assign n66988 = ~n67013;
  assign n67001 = n67014 & n63982;
  assign n66989 = ~n66990;
  assign n67024 = n66980 & n338;
  assign n67034 = ~n66980;
  assign n67015 = n67057 ^ n67058;
  assign n67048 = ~n67057;
  assign n63129 = n67068 ^ n67069;
  assign n66919 = n67071 & n67072;
  assign n67062 = ~n67077;
  assign n67092 = n67100 & n67101;
  assign n66921 = n66861 & n4867;
  assign n66926 = ~n66861;
  assign n62769 = n66961 ^ n66962;
  assign n66940 = ~n66965;
  assign n66937 = ~n66970;
  assign n66959 = ~n66981;
  assign n66986 = n66988 & n66989;
  assign n66958 = ~n67001;
  assign n66978 = n339 ^ n67015;
  assign n66944 = ~n67024;
  assign n67012 = n67034 & n12767;
  assign n67037 = n67048 & n67049;
  assign n67044 = n66919 & n67053;
  assign n67039 = n63129 & n65583;
  assign n67046 = n63129 & n65389;
  assign n63166 = ~n63129;
  assign n67045 = ~n66919;
  assign n67025 = n67062 & n67063;
  assign n67065 = ~n67092;
  assign n66868 = ~n66921;
  assign n66918 = n66926 & n357;
  assign n66923 = n62769 & n63982;
  assign n66906 = n66937 & n66903;
  assign n66873 = n66939 & n66940;
  assign n62802 = ~n62769;
  assign n66933 = n66937 & n66907;
  assign n66924 = n66959 & n66960;
  assign n66878 = n66976 ^ n66978;
  assign n66957 = ~n66986;
  assign n66975 = ~n66978;
  assign n66985 = ~n67012;
  assign n66996 = n67025 ^ n67026;
  assign n67019 = ~n67037;
  assign n67023 = n63166 & n67038;
  assign n67030 = n63166 & n64457;
  assign n65626 = ~n67039;
  assign n66956 = ~n67044;
  assign n67029 = n67045 & n66948;
  assign n67005 = ~n67046;
  assign n67027 = ~n67025;
  assign n67040 = n67065 & n67066;
  assign n64534 = n66906 ^ n66907;
  assign n66836 = ~n66918;
  assign n66871 = ~n66923;
  assign n66874 = n66924 ^ n66925;
  assign n66913 = n66873 & n66925;
  assign n66908 = n62802 & n65799;
  assign n66902 = ~n66933;
  assign n66900 = ~n66873;
  assign n66877 = ~n66924;
  assign n66922 = n66957 & n66958;
  assign n66946 = n66878 & n63959;
  assign n66942 = ~n66878;
  assign n66904 = n66975 & n66976;
  assign n66912 = n66995 ^ n66996;
  assign n66979 = n67019 & n67020;
  assign n65591 = ~n67023;
  assign n67018 = n67027 & n67028;
  assign n66928 = ~n67029;
  assign n67004 = ~n67030;
  assign n67002 = n67040 ^ n67041;
  assign n67042 = ~n67040;
  assign n66794 = n66873 ^ n66874;
  assign n64556 = ~n64534;
  assign n66899 = n66900 & n66901;
  assign n66860 = n66902 & n66903;
  assign n66872 = ~n66908;
  assign n66876 = ~n66913;
  assign n66879 = n66922 ^ n63934;
  assign n66916 = ~n66922;
  assign n66936 = n66942 & n63934;
  assign n66858 = ~n66946;
  assign n66951 = n66912 & n12734;
  assign n66945 = n66979 ^ n66980;
  assign n66963 = ~n66912;
  assign n63091 = n64361 ^ n67002;
  assign n66881 = n67004 & n67005;
  assign n66984 = ~n66979;
  assign n66997 = ~n67018;
  assign n67006 = ~n67002;
  assign n67031 = n67042 & n67043;
  assign n66840 = n66794 & n4824;
  assign n66834 = n66860 ^ n66861;
  assign n66839 = ~n66794;
  assign n66763 = n66871 & n66872;
  assign n66866 = n66876 & n66877;
  assign n62698 = n66878 ^ n66879;
  assign n66869 = ~n66860;
  assign n66844 = ~n66899;
  assign n66917 = ~n66936;
  assign n66905 = n338 ^ n66945;
  assign n66915 = ~n66951;
  assign n66941 = n66963 & n337;
  assign n66971 = n66984 & n66985;
  assign n66969 = n66881 & n66838;
  assign n66968 = n63091 & n66987;
  assign n66972 = ~n66881;
  assign n63135 = ~n63091;
  assign n66947 = n66997 & n66998;
  assign n66991 = n67006 & n64361;
  assign n67007 = ~n67031;
  assign n66777 = n357 ^ n66834;
  assign n66824 = n66839 & n356;
  assign n66781 = ~n66840;
  assign n66841 = n66763 & n66852;
  assign n66842 = n62698 & n63959;
  assign n66847 = ~n66763;
  assign n66843 = ~n66866;
  assign n62732 = ~n62698;
  assign n66848 = n66868 & n66869;
  assign n66789 = n66904 ^ n66905;
  assign n66889 = n66916 & n66917;
  assign n66820 = n66905 & n66904;
  assign n66864 = ~n66941;
  assign n66920 = n66947 ^ n66948;
  assign n66952 = n63135 & n65381;
  assign n65495 = ~n66968;
  assign n66883 = ~n66969;
  assign n66943 = ~n66971;
  assign n66964 = n66972 & n66973;
  assign n66953 = n63135 & n65538;
  assign n66955 = ~n66947;
  assign n66935 = ~n66991;
  assign n66974 = n67007 & n67008;
  assign n65558 = n66777 ^ n64534;
  assign n66779 = ~n66777;
  assign n66757 = ~n66824;
  assign n66805 = ~n66841;
  assign n66798 = ~n66842;
  assign n66795 = n66843 & n66844;
  assign n66830 = n62732 & n65701;
  assign n66825 = n66847 & n66796;
  assign n66835 = ~n66848;
  assign n66862 = n66789 & n63935;
  assign n66857 = ~n66889;
  assign n66867 = ~n66789;
  assign n66832 = n66919 ^ n66920;
  assign n66911 = n66943 & n66944;
  assign n66934 = ~n66952;
  assign n65550 = ~n66953;
  assign n66938 = n66955 & n66956;
  assign n66846 = ~n66964;
  assign n66930 = n66974 ^ n64340;
  assign n66966 = ~n66974;
  assign n65556 = ~n65558;
  assign n66699 = n66779 & n64556;
  assign n66764 = n66795 ^ n66796;
  assign n66768 = ~n66825;
  assign n66806 = ~n66795;
  assign n66799 = ~n66830;
  assign n66793 = n66835 & n66836;
  assign n66826 = n66857 & n66858;
  assign n66821 = ~n66862;
  assign n66853 = n66867 & n63899;
  assign n66875 = n66832 & n336;
  assign n66888 = ~n66832;
  assign n66870 = n66911 ^ n66912;
  assign n63047 = n66929 ^ n66930;
  assign n66809 = n66934 & n66935;
  assign n66914 = ~n66911;
  assign n66927 = ~n66938;
  assign n66954 = n66966 & n66967;
  assign n66697 = n66763 ^ n66764;
  assign n66748 = n66793 ^ n66794;
  assign n66678 = n66798 & n66799;
  assign n66792 = n66805 & n66806;
  assign n66782 = ~n66793;
  assign n66790 = n66826 ^ n63899;
  assign n66788 = ~n66853;
  assign n66822 = ~n66826;
  assign n66833 = n337 ^ n66870;
  assign n66785 = ~n66875;
  assign n66865 = n66888 & n12647;
  assign n66894 = n63047 & n65282;
  assign n66892 = n63047 & n66909;
  assign n66893 = n66809 & n66910;
  assign n66897 = n66914 & n66915;
  assign n66898 = ~n66809;
  assign n63065 = ~n63047;
  assign n66880 = n66927 & n66928;
  assign n66931 = ~n66954;
  assign n66718 = n66697 & n355;
  assign n66713 = n356 ^ n66748;
  assign n66729 = ~n66697;
  assign n66760 = n66678 & n66731;
  assign n66771 = n66781 & n66782;
  assign n66761 = ~n66678;
  assign n62644 = n66789 ^ n66790;
  assign n66767 = ~n66792;
  assign n66811 = n66821 & n66822;
  assign n66701 = n66820 ^ n66833;
  assign n66819 = ~n66833;
  assign n66829 = ~n66865;
  assign n66837 = n66880 ^ n66881;
  assign n65465 = ~n66892;
  assign n66802 = ~n66893;
  assign n66850 = ~n66894;
  assign n66885 = n63065 & n65421;
  assign n66863 = ~n66897;
  assign n66887 = n66898 & n66766;
  assign n66884 = n63065 & n64340;
  assign n66882 = ~n66880;
  assign n66895 = n66931 & n66932;
  assign n64461 = n66699 ^ n66713;
  assign n66640 = ~n66718;
  assign n66700 = n66729 & n4762;
  assign n66698 = ~n66713;
  assign n66721 = ~n66760;
  assign n66747 = n66761 & n66762;
  assign n66746 = n62644 & n63899;
  assign n66730 = n66767 & n66768;
  assign n66756 = ~n66771;
  assign n62656 = ~n62644;
  assign n66780 = n66701 & n63868;
  assign n66787 = ~n66811;
  assign n66791 = ~n66701;
  assign n66752 = n66819 & n66820;
  assign n66750 = n66837 ^ n66838;
  assign n66831 = n66863 & n66864;
  assign n66859 = n66882 & n66883;
  assign n66849 = ~n66884;
  assign n65420 = ~n66885;
  assign n66759 = ~n66887;
  assign n66851 = n66895 ^ n66896;
  assign n66890 = ~n66895;
  assign n65470 = ~n64461;
  assign n66615 = n66698 & n66699;
  assign n66686 = ~n66700;
  assign n66679 = n66730 ^ n66731;
  assign n66714 = ~n66746;
  assign n66685 = ~n66747;
  assign n66722 = ~n66730;
  assign n66735 = n62656 & n65619;
  assign n66696 = n66756 & n66757;
  assign n66704 = ~n66780;
  assign n66751 = n66787 & n66788;
  assign n66776 = n66791 & n63891;
  assign n66800 = n66750 & n12617;
  assign n66797 = ~n66750;
  assign n66778 = n66831 ^ n66832;
  assign n66725 = n66849 & n66850;
  assign n62972 = n64296 ^ n66851;
  assign n66828 = ~n66831;
  assign n66845 = ~n66859;
  assign n66854 = n66851 & n64320;
  assign n66886 = n66890 & n66891;
  assign n66601 = n66678 ^ n66679;
  assign n66668 = n66696 ^ n66697;
  assign n66707 = n66721 & n66722;
  assign n66687 = ~n66696;
  assign n66715 = ~n66735;
  assign n66702 = n66751 ^ n63868;
  assign n66744 = ~n66751;
  assign n66745 = ~n66776;
  assign n66753 = n336 ^ n66778;
  assign n66783 = n66797 & n351;
  assign n66755 = ~n66800;
  assign n66813 = n66725 & n66823;
  assign n66814 = n62972 & n66827;
  assign n66818 = n66828 & n66829;
  assign n66815 = ~n66725;
  assign n63023 = ~n62972;
  assign n66808 = n66845 & n66846;
  assign n66770 = ~n66854;
  assign n66855 = ~n66886;
  assign n66649 = n66601 & n4727;
  assign n66633 = ~n66601;
  assign n66616 = n355 ^ n66668;
  assign n66676 = n66686 & n66687;
  assign n62588 = n66701 ^ n66702;
  assign n66684 = ~n66707;
  assign n66606 = n66714 & n66715;
  assign n66736 = n66744 & n66745;
  assign n66629 = n66752 ^ n66753;
  assign n66666 = n66753 & n66752;
  assign n66710 = ~n66783;
  assign n66765 = n66808 ^ n66809;
  assign n66804 = n63023 & n65207;
  assign n66717 = ~n66813;
  assign n65330 = ~n66814;
  assign n66803 = n66815 & n66681;
  assign n66810 = n63023 & n65325;
  assign n66784 = ~n66818;
  assign n66801 = ~n66808;
  assign n66812 = n66855 & n66856;
  assign n64417 = n66615 ^ n66616;
  assign n66631 = n66633 & n354;
  assign n66604 = ~n66649;
  assign n66517 = n66616 & n66615;
  assign n66639 = ~n66676;
  assign n66664 = n62588 & n65502;
  assign n66647 = n66684 & n66685;
  assign n66669 = n66606 & n66688;
  assign n62603 = ~n62588;
  assign n66663 = ~n66606;
  assign n66711 = n66629 & n63828;
  assign n66703 = ~n66736;
  assign n66712 = ~n66629;
  assign n66673 = n66765 ^ n66766;
  assign n66749 = n66784 & n66785;
  assign n66786 = n66801 & n66802;
  assign n66683 = ~n66803;
  assign n66769 = ~n66804;
  assign n65369 = ~n66810;
  assign n66773 = n66812 ^ n64253;
  assign n66816 = ~n66812;
  assign n65393 = ~n64417;
  assign n66554 = ~n66631;
  assign n66600 = n66639 & n66640;
  assign n66607 = n66647 ^ n66648;
  assign n66652 = n66663 & n66648;
  assign n66644 = ~n66647;
  assign n66659 = n62603 & n63868;
  assign n66620 = ~n66664;
  assign n66643 = ~n66669;
  assign n66667 = n66703 & n66704;
  assign n66675 = ~n66711;
  assign n66693 = n66712 & n63831;
  assign n66728 = n66673 & n350;
  assign n66706 = n66749 ^ n66750;
  assign n66719 = ~n66673;
  assign n66754 = ~n66749;
  assign n66602 = n66769 & n66770;
  assign n62897 = n66772 ^ n66773;
  assign n66758 = ~n66786;
  assign n66807 = n66816 & n66817;
  assign n66552 = n66600 ^ n66601;
  assign n66528 = n66606 ^ n66607;
  assign n66605 = ~n66600;
  assign n66627 = n66643 & n66644;
  assign n66597 = ~n66652;
  assign n66619 = ~n66659;
  assign n66630 = n66667 ^ n63828;
  assign n66625 = ~n66693;
  assign n66674 = ~n66667;
  assign n66677 = n351 ^ n66706;
  assign n66705 = n66719 & n12503;
  assign n66618 = ~n66728;
  assign n66738 = n62897 & n65232;
  assign n66741 = n62897 & n64287;
  assign n66740 = n66602 & n66637;
  assign n66739 = n66754 & n66755;
  assign n66724 = n66758 & n66759;
  assign n66742 = ~n66602;
  assign n62954 = ~n62897;
  assign n66774 = ~n66807;
  assign n66518 = n354 ^ n66552;
  assign n66557 = n66528 & n353;
  assign n66556 = ~n66528;
  assign n66595 = n66604 & n66605;
  assign n66519 = n66619 & n66620;
  assign n66596 = ~n66627;
  assign n62539 = n66629 ^ n66630;
  assign n66662 = n66674 & n66675;
  assign n66550 = n66666 ^ n66677;
  assign n66665 = ~n66677;
  assign n66671 = ~n66705;
  assign n66680 = n66724 ^ n66725;
  assign n66726 = n62954 & n66734;
  assign n65245 = ~n66738;
  assign n66727 = n62954 & n65084;
  assign n66709 = ~n66739;
  assign n66646 = ~n66740;
  assign n66689 = ~n66741;
  assign n66723 = n66742 & n66743;
  assign n66716 = ~n66724;
  assign n66737 = n66774 & n66775;
  assign n64378 = n66517 ^ n66518;
  assign n66531 = ~n66518;
  assign n66545 = n66556 & n4683;
  assign n66487 = ~n66557;
  assign n66553 = ~n66595;
  assign n66558 = n66596 & n66597;
  assign n66590 = n66519 & n66559;
  assign n66587 = n62539 & n65408;
  assign n66593 = ~n66519;
  assign n62568 = ~n62539;
  assign n66621 = n66550 & n63795;
  assign n66628 = ~n66550;
  assign n66624 = ~n66662;
  assign n66584 = n66665 & n66666;
  assign n66583 = n66680 ^ n66681;
  assign n66672 = n66709 & n66710;
  assign n66708 = n66716 & n66717;
  assign n66599 = ~n66723;
  assign n65297 = ~n66726;
  assign n66690 = ~n66727;
  assign n66692 = n66737 ^ n64212;
  assign n66732 = ~n66737;
  assign n65280 = ~n64378;
  assign n66453 = n66531 & n66517;
  assign n66515 = ~n66545;
  assign n66527 = n66553 & n66554;
  assign n66520 = n66558 ^ n66559;
  assign n66548 = ~n66587;
  assign n66560 = ~n66590;
  assign n66578 = n62568 & n63831;
  assign n66561 = ~n66558;
  assign n66573 = n66593 & n66594;
  assign n66543 = ~n66621;
  assign n66586 = n66624 & n66625;
  assign n66612 = n66628 & n63772;
  assign n66642 = n66583 & n349;
  assign n66634 = ~n66583;
  assign n66622 = n66672 ^ n66673;
  assign n66529 = n66689 & n66690;
  assign n62820 = n66691 ^ n66692;
  assign n66670 = ~n66672;
  assign n66682 = ~n66708;
  assign n66720 = n66732 & n66733;
  assign n66450 = ~n66453;
  assign n66446 = n66519 ^ n66520;
  assign n66483 = n66527 ^ n66528;
  assign n66516 = ~n66527;
  assign n66541 = n66560 & n66561;
  assign n66526 = ~n66573;
  assign n66549 = ~n66578;
  assign n66551 = n66586 ^ n63772;
  assign n66588 = ~n66586;
  assign n66589 = ~n66612;
  assign n66585 = n350 ^ n66622;
  assign n66626 = n66634 & n12444;
  assign n66538 = ~n66642;
  assign n66654 = n62820 & n64212;
  assign n66650 = n66670 & n66671;
  assign n66656 = n62820 & n65146;
  assign n66655 = n66529 & n66564;
  assign n66636 = n66682 & n66683;
  assign n62881 = ~n62820;
  assign n66657 = ~n66529;
  assign n66694 = ~n66720;
  assign n66454 = n353 ^ n66483;
  assign n66482 = n66446 & n4635;
  assign n66477 = ~n66446;
  assign n66513 = n66515 & n66516;
  assign n66525 = ~n66541;
  assign n66457 = n66548 & n66549;
  assign n62495 = n66550 ^ n66551;
  assign n66467 = n66584 ^ n66585;
  assign n66574 = n66588 & n66589;
  assign n66505 = n66585 & n66584;
  assign n66592 = ~n66626;
  assign n66603 = n66636 ^ n66637;
  assign n66617 = ~n66650;
  assign n66641 = n62881 & n66653;
  assign n66608 = ~n66654;
  assign n66566 = ~n66655;
  assign n65151 = ~n66656;
  assign n66632 = n66657 & n66658;
  assign n66635 = n62881 & n65024;
  assign n66645 = ~n66636;
  assign n66651 = n66694 & n66695;
  assign n64345 = n66453 ^ n66454;
  assign n66449 = ~n66454;
  assign n66462 = n66477 & n352;
  assign n66443 = ~n66482;
  assign n66486 = ~n66513;
  assign n66511 = n66457 & n66521;
  assign n66491 = n66525 & n66526;
  assign n66512 = n62495 & n63795;
  assign n66514 = ~n66457;
  assign n62529 = ~n62495;
  assign n66539 = n66467 & n63734;
  assign n66542 = ~n66574;
  assign n66546 = ~n66467;
  assign n66508 = n66602 ^ n66603;
  assign n66582 = n66617 & n66618;
  assign n66523 = ~n66632;
  assign n66609 = ~n66635;
  assign n65205 = ~n66641;
  assign n66623 = n66645 & n66646;
  assign n66611 = n66651 ^ n64166;
  assign n66660 = ~n66651;
  assign n65213 = ~n64345;
  assign n66387 = n66449 & n66450;
  assign n66423 = ~n66462;
  assign n66445 = n66486 & n66487;
  assign n66458 = n66491 ^ n66492;
  assign n66488 = ~n66511;
  assign n66495 = n62529 & n65328;
  assign n66474 = ~n66512;
  assign n66489 = ~n66491;
  assign n66494 = n66514 & n66492;
  assign n66503 = ~n66539;
  assign n66504 = n66542 & n66543;
  assign n66536 = n66546 & n63756;
  assign n66562 = n66508 & n12352;
  assign n66540 = n66582 ^ n66583;
  assign n66555 = ~n66508;
  assign n66447 = n66608 & n66609;
  assign n62749 = n66610 ^ n66611;
  assign n66591 = ~n66582;
  assign n66598 = ~n66623;
  assign n66638 = n66660 & n66661;
  assign n66390 = ~n66387;
  assign n66416 = n66445 ^ n66446;
  assign n66377 = n66457 ^ n66458;
  assign n66444 = ~n66445;
  assign n66475 = n66488 & n66489;
  assign n66452 = ~n66494;
  assign n66473 = ~n66495;
  assign n66468 = n66504 ^ n63734;
  assign n66470 = ~n66536;
  assign n66502 = ~n66504;
  assign n66506 = n349 ^ n66540;
  assign n66544 = n66555 & n348;
  assign n66510 = ~n66562;
  assign n66575 = n66591 & n66592;
  assign n66572 = n62749 & n65071;
  assign n66577 = n66447 & n66481;
  assign n66576 = n62749 & n64942;
  assign n66563 = n66598 & n66599;
  assign n66570 = ~n66447;
  assign n62751 = ~n62749;
  assign n66613 = ~n66638;
  assign n66388 = n352 ^ n66416;
  assign n66412 = n66377 & n367;
  assign n66421 = ~n66377;
  assign n66442 = n66443 & n66444;
  assign n62458 = n66467 ^ n66468;
  assign n66391 = n66473 & n66474;
  assign n66451 = ~n66475;
  assign n66496 = n66502 & n66503;
  assign n66395 = n66505 ^ n66506;
  assign n66435 = n66506 & n66505;
  assign n66464 = ~n66544;
  assign n66530 = n66563 ^ n66564;
  assign n66569 = n66570 & n66571;
  assign n66568 = n62751 & n64168;
  assign n65109 = ~n66572;
  assign n66537 = ~n66575;
  assign n66534 = ~n66576;
  assign n66485 = ~n66577;
  assign n66567 = n62751 & n66581;
  assign n66565 = ~n66563;
  assign n66579 = n66613 & n66614;
  assign n64307 = n66387 ^ n66388;
  assign n66389 = ~n66388;
  assign n66355 = ~n66412;
  assign n66398 = n66421 & n4592;
  assign n66422 = ~n66442;
  assign n66419 = n66451 & n66452;
  assign n66432 = n66391 & n66420;
  assign n66431 = n62458 & n65268;
  assign n66439 = ~n66391;
  assign n62481 = ~n62458;
  assign n66472 = n66395 & n63672;
  assign n66465 = ~n66395;
  assign n66469 = ~n66496;
  assign n66438 = n66529 ^ n66530;
  assign n66507 = n66537 & n66538;
  assign n66547 = n66565 & n66566;
  assign n65074 = ~n66567;
  assign n66535 = ~n66568;
  assign n66456 = ~n66569;
  assign n62754 = n66579 ^ n66580;
  assign n65110 = ~n64307;
  assign n66325 = n66389 & n66390;
  assign n66383 = ~n66398;
  assign n66392 = n66419 ^ n66420;
  assign n66376 = n66422 & n66423;
  assign n66414 = ~n66419;
  assign n66399 = ~n66431;
  assign n66425 = n62481 & n63756;
  assign n66413 = ~n66432;
  assign n66424 = n66439 & n66440;
  assign n66461 = n66465 & n63728;
  assign n66428 = n66469 & n66470;
  assign n66434 = ~n66472;
  assign n66479 = n66438 & n12313;
  assign n66466 = n66507 ^ n66508;
  assign n66490 = ~n66438;
  assign n66509 = ~n66507;
  assign n66380 = n66534 & n66535;
  assign n66522 = ~n66547;
  assign n66533 = n62754 & n64875;
  assign n66532 = ~n62754;
  assign n66346 = n66376 ^ n66377;
  assign n66324 = n66391 ^ n66392;
  assign n66384 = ~n66376;
  assign n66397 = n66413 & n66414;
  assign n66379 = ~n66424;
  assign n66400 = ~n66425;
  assign n66396 = n66428 ^ n63672;
  assign n66433 = ~n66428;
  assign n66407 = ~n66461;
  assign n66436 = n348 ^ n66466;
  assign n66430 = ~n66479;
  assign n66476 = n66490 & n347;
  assign n66497 = n66509 & n66510;
  assign n66493 = n66380 & n66410;
  assign n66480 = n66522 & n66523;
  assign n66498 = ~n66380;
  assign n66524 = n66532 & n64171;
  assign n66500 = ~n66533;
  assign n66326 = n367 ^ n66346;
  assign n66347 = n66324 & n4556;
  assign n66350 = ~n66324;
  assign n66365 = n66383 & n66384;
  assign n62425 = n66395 ^ n66396;
  assign n66378 = ~n66397;
  assign n66317 = n66399 & n66400;
  assign n66426 = n66433 & n66434;
  assign n66341 = n66435 ^ n66436;
  assign n66441 = ~n66436;
  assign n66405 = ~n66476;
  assign n66448 = n66480 ^ n66481;
  assign n66418 = ~n66493;
  assign n66463 = ~n66497;
  assign n66478 = n66498 & n66499;
  assign n66484 = ~n66480;
  assign n66501 = ~n66524;
  assign n64259 = n66325 ^ n66326;
  assign n66269 = n66326 & n66325;
  assign n66328 = ~n66347;
  assign n66335 = n66350 & n366;
  assign n66354 = ~n66365;
  assign n66356 = n66378 & n66379;
  assign n66367 = n66317 & n66382;
  assign n66366 = n62425 & n65183;
  assign n62443 = ~n62425;
  assign n66364 = ~n66317;
  assign n66394 = n66341 & n63655;
  assign n66406 = ~n66426;
  assign n66403 = ~n66341;
  assign n66362 = n66441 & n66435;
  assign n66373 = n66447 ^ n66448;
  assign n66437 = n66463 & n66464;
  assign n66386 = ~n66478;
  assign n66471 = n66484 & n66485;
  assign n66459 = n66500 & n66501;
  assign n65025 = ~n64259;
  assign n66297 = ~n66335;
  assign n66323 = n66354 & n66355;
  assign n66318 = n66356 ^ n66357;
  assign n66352 = ~n66356;
  assign n66359 = n66364 & n66357;
  assign n66333 = ~n66366;
  assign n66351 = ~n66367;
  assign n66358 = n62443 & n63728;
  assign n66337 = ~n66394;
  assign n66393 = n66403 & n63690;
  assign n66368 = n66406 & n66407;
  assign n66415 = n66373 & n12199;
  assign n66408 = n66437 ^ n66438;
  assign n66411 = ~n66373;
  assign n66322 = n66459 ^ n66460;
  assign n66429 = ~n66437;
  assign n66455 = ~n66471;
  assign n66275 = n66317 ^ n66318;
  assign n66294 = n66323 ^ n66324;
  assign n66327 = ~n66323;
  assign n66332 = n66351 & n66352;
  assign n66334 = ~n66358;
  assign n66330 = ~n66359;
  assign n66342 = n66368 ^ n63655;
  assign n66370 = ~n66393;
  assign n66369 = ~n66368;
  assign n66363 = n347 ^ n66408;
  assign n66401 = n66411 & n346;
  assign n66375 = ~n66415;
  assign n66427 = n66429 & n66430;
  assign n66409 = n66455 & n66456;
  assign n66270 = n366 ^ n66294;
  assign n66295 = n66275 & n365;
  assign n66293 = ~n66275;
  assign n66306 = n66327 & n66328;
  assign n66329 = ~n66332;
  assign n66319 = n66333 & n66334;
  assign n62389 = n66341 ^ n66342;
  assign n66284 = n66362 ^ n66363;
  assign n66361 = n66369 & n66370;
  assign n66371 = ~n66363;
  assign n66340 = ~n66401;
  assign n66381 = n66409 ^ n66410;
  assign n66404 = ~n66427;
  assign n66417 = ~n66409;
  assign n64939 = n66269 ^ n66270;
  assign n66276 = ~n66270;
  assign n66282 = n66293 & n4506;
  assign n66244 = ~n66295;
  assign n66296 = ~n66306;
  assign n66309 = n66319 & n66320;
  assign n66303 = n62389 & n65061;
  assign n66266 = n66329 & n66330;
  assign n66307 = ~n66319;
  assign n62383 = ~n62389;
  assign n66343 = n66284 & n63613;
  assign n66345 = ~n66284;
  assign n66336 = ~n66361;
  assign n66304 = n66371 & n66362;
  assign n66314 = n66380 ^ n66381;
  assign n66372 = n66404 & n66405;
  assign n66402 = n66417 & n66418;
  assign n66222 = n66276 & n66269;
  assign n66267 = ~n66282;
  assign n66274 = n66296 & n66297;
  assign n66287 = ~n66303;
  assign n66292 = ~n66266;
  assign n66298 = n66307 & n66308;
  assign n66280 = ~n66309;
  assign n66299 = n62383 & n63655;
  assign n66302 = n66336 & n66337;
  assign n66279 = ~n66343;
  assign n66331 = n66345 & n63642;
  assign n66353 = n66314 & n12147;
  assign n66338 = n66372 ^ n66373;
  assign n66348 = ~n66314;
  assign n66374 = ~n66372;
  assign n66385 = ~n66402;
  assign n66247 = n66274 ^ n66275;
  assign n66268 = ~n66274;
  assign n66291 = n66292 & n66280;
  assign n66273 = ~n66298;
  assign n66288 = ~n66299;
  assign n66285 = n66302 ^ n63613;
  assign n66316 = ~n66331;
  assign n66315 = ~n66302;
  assign n66305 = n346 ^ n66338;
  assign n66344 = n66348 & n345;
  assign n66312 = ~n66353;
  assign n66360 = n66374 & n66375;
  assign n66349 = n66385 & n66386;
  assign n66223 = n365 ^ n66247;
  assign n66253 = n66267 & n66268;
  assign n66265 = n66273 & n66280;
  assign n62332 = n66284 ^ n66285;
  assign n66249 = n66287 & n66288;
  assign n66272 = ~n66291;
  assign n66238 = n66304 ^ n66305;
  assign n66300 = n66315 & n66316;
  assign n66310 = ~n66305;
  assign n66290 = ~n66344;
  assign n66321 = n344 ^ n66349;
  assign n66339 = ~n66360;
  assign n66200 = n66222 ^ n66223;
  assign n66176 = n66223 & n66222;
  assign n66243 = ~n66253;
  assign n66219 = n66265 ^ n66266;
  assign n66254 = n66249 & n66271;
  assign n66248 = n66272 & n66273;
  assign n66255 = n62332 & n65013;
  assign n66264 = ~n66249;
  assign n62359 = ~n62332;
  assign n66283 = n66238 & n63591;
  assign n66278 = ~n66300;
  assign n66286 = ~n66238;
  assign n66259 = n66310 & n66304;
  assign n66263 = n66321 ^ n66322;
  assign n66313 = n66339 & n66340;
  assign n62048 = n66200 ^ n63131;
  assign n66201 = n66200 & n63113;
  assign n66197 = ~n66200;
  assign n66183 = ~n66176;
  assign n66218 = n66243 & n66244;
  assign n66224 = n66248 ^ n66249;
  assign n66233 = n66219 & n4471;
  assign n66230 = ~n66219;
  assign n66251 = n62359 & n63613;
  assign n66245 = ~n66248;
  assign n66246 = ~n66254;
  assign n66241 = ~n66255;
  assign n66250 = n66264 & n66225;
  assign n66256 = n66278 & n66279;
  assign n66232 = ~n66283;
  assign n66277 = n66286 & n63548;
  assign n66281 = n66313 ^ n66314;
  assign n66311 = ~n66313;
  assign n66180 = ~n62048;
  assign n66086 = n66197 & n63113;
  assign n66150 = ~n66201;
  assign n66196 = n66218 ^ n66219;
  assign n66174 = n66224 ^ n66225;
  assign n66226 = ~n66218;
  assign n66228 = n66230 & n364;
  assign n66227 = ~n66233;
  assign n66234 = n66245 & n66246;
  assign n66221 = ~n66250;
  assign n66242 = ~n66251;
  assign n66239 = n66256 ^ n63548;
  assign n66257 = ~n66256;
  assign n66258 = ~n66277;
  assign n66260 = n345 ^ n66281;
  assign n66301 = n66311 & n66312;
  assign n66163 = n66180 & n64200;
  assign n66177 = n364 ^ n66196;
  assign n66202 = n66174 & n363;
  assign n66203 = ~n66174;
  assign n66217 = n66226 & n66227;
  assign n66195 = ~n66228;
  assign n66220 = ~n66234;
  assign n62297 = n66238 ^ n66239;
  assign n66171 = n66241 & n66242;
  assign n66252 = n66257 & n66258;
  assign n66190 = n66259 ^ n66260;
  assign n66261 = ~n66260;
  assign n66289 = ~n66301;
  assign n66149 = ~n66163;
  assign n66161 = n66176 ^ n66177;
  assign n66131 = n66177 & n66183;
  assign n66147 = ~n66202;
  assign n66187 = n66203 & n4427;
  assign n66194 = ~n66217;
  assign n66211 = n66171 & n66193;
  assign n66192 = n66220 & n66221;
  assign n66210 = n62297 & n63591;
  assign n66208 = ~n66171;
  assign n62323 = ~n62297;
  assign n66235 = n66190 & n63556;
  assign n66240 = ~n66190;
  assign n66231 = ~n66252;
  assign n66236 = n66261 & n66259;
  assign n66262 = n66289 & n66290;
  assign n66130 = n66149 & n66150;
  assign n66148 = n66161 & n63022;
  assign n66154 = ~n66161;
  assign n66134 = ~n66131;
  assign n66182 = ~n66187;
  assign n66172 = n66192 ^ n66193;
  assign n66173 = n66194 & n66195;
  assign n66207 = n66208 & n66209;
  assign n66206 = n62323 & n64906;
  assign n66198 = ~n66192;
  assign n66189 = ~n66210;
  assign n66199 = ~n66211;
  assign n66212 = n66231 & n66232;
  assign n66186 = ~n66235;
  assign n66229 = n66240 & n63530;
  assign n66237 = n66262 ^ n66263;
  assign n66093 = n66130 ^ n66125;
  assign n66124 = ~n66130;
  assign n66133 = ~n66148;
  assign n66136 = n66154 & n63020;
  assign n66120 = n66171 ^ n66172;
  assign n66153 = n66173 ^ n66174;
  assign n66181 = ~n66173;
  assign n66184 = n66198 & n66199;
  assign n66188 = ~n66206;
  assign n66179 = ~n66207;
  assign n66191 = n66212 ^ n63530;
  assign n66215 = ~n66212;
  assign n66216 = ~n66229;
  assign n66167 = n66236 ^ n66237;
  assign n63941 = n391 ^ n66093;
  assign n66094 = ~n66093;
  assign n65928 = n66124 & n66125;
  assign n66121 = n66133 & n66086;
  assign n66109 = ~n66136;
  assign n66132 = n363 ^ n66153;
  assign n66145 = n66120 & n4376;
  assign n66157 = ~n66120;
  assign n66162 = n66181 & n66182;
  assign n66178 = ~n66184;
  assign n66122 = n66188 & n66189;
  assign n62258 = n66190 ^ n66191;
  assign n66204 = n66215 & n66216;
  assign n66213 = n66167 & n63523;
  assign n66214 = ~n66167;
  assign n65635 = ~n63941;
  assign n65813 = n66094 & n391;
  assign n66108 = ~n66121;
  assign n66055 = n66131 ^ n66132;
  assign n66114 = n66133 & n66109;
  assign n66072 = n66132 & n66134;
  assign n66128 = ~n66145;
  assign n66139 = n66157 & n362;
  assign n66146 = ~n66162;
  assign n66165 = n66122 & n66175;
  assign n66151 = n66178 & n66179;
  assign n66164 = n62258 & n63556;
  assign n62286 = ~n62258;
  assign n66170 = ~n66122;
  assign n66185 = ~n66204;
  assign n66169 = ~n66213;
  assign n66205 = n66214 & n63479;
  assign n66092 = n66055 & n62915;
  assign n66079 = n66108 & n66109;
  assign n66103 = ~n66055;
  assign n66087 = ~n66114;
  assign n66078 = ~n66072;
  assign n66102 = ~n66139;
  assign n66119 = n66146 & n66147;
  assign n66123 = n66151 ^ n66152;
  assign n66159 = n62286 & n64851;
  assign n66155 = ~n66151;
  assign n66144 = ~n66164;
  assign n66156 = ~n66165;
  assign n66158 = n66170 & n66152;
  assign n66166 = n66185 & n66186;
  assign n66138 = ~n66205;
  assign n66056 = n66079 ^ n62915;
  assign n61962 = n66086 ^ n66087;
  assign n66041 = ~n66092;
  assign n66071 = ~n66079;
  assign n66090 = n66103 & n62957;
  assign n66100 = n66119 ^ n66120;
  assign n66039 = n66122 ^ n66123;
  assign n66129 = ~n66119;
  assign n66142 = n66155 & n66156;
  assign n66127 = ~n66158;
  assign n66143 = ~n66159;
  assign n66141 = n66166 ^ n66167;
  assign n66168 = ~n66166;
  assign n61852 = n66055 ^ n66056;
  assign n66061 = n61962 & n64106;
  assign n61956 = ~n61962;
  assign n66070 = ~n66090;
  assign n66073 = n362 ^ n66100;
  assign n66099 = n66039 & n361;
  assign n66104 = ~n66039;
  assign n66110 = n66128 & n66129;
  assign n62203 = n63479 ^ n66141;
  assign n66126 = ~n66142;
  assign n66066 = n66143 & n66144;
  assign n66140 = ~n66141;
  assign n66160 = n66168 & n66169;
  assign n66025 = n61852 & n64051;
  assign n61889 = ~n61852;
  assign n66051 = n61956 & n63020;
  assign n66032 = ~n66061;
  assign n66065 = n66070 & n66071;
  assign n65979 = n66072 ^ n66073;
  assign n66012 = n66073 & n66078;
  assign n66050 = ~n66099;
  assign n66082 = n66104 & n4334;
  assign n66101 = ~n66110;
  assign n66095 = n66126 & n66127;
  assign n66113 = n66066 & n66096;
  assign n66111 = ~n66066;
  assign n62250 = ~n62203;
  assign n66135 = n66140 & n63479;
  assign n66137 = ~n66160;
  assign n65991 = ~n66025;
  assign n66011 = n61889 & n62915;
  assign n66042 = n65979 & n62837;
  assign n66031 = ~n66051;
  assign n66045 = ~n65979;
  assign n66040 = ~n66065;
  assign n66024 = ~n66012;
  assign n66077 = ~n66082;
  assign n66067 = n66095 ^ n66096;
  assign n66068 = n66101 & n66102;
  assign n66105 = n66111 & n66112;
  assign n66098 = ~n66113;
  assign n66097 = ~n66095;
  assign n66106 = n62250 & n64793;
  assign n66084 = ~n66135;
  assign n66115 = n66137 & n66138;
  assign n65990 = ~n66011;
  assign n66015 = n66031 & n66032;
  assign n66014 = n66040 & n66041;
  assign n66010 = ~n66042;
  assign n66027 = n66045 & n62853;
  assign n66022 = n66066 ^ n66067;
  assign n66038 = n361 ^ n66068;
  assign n66076 = ~n66068;
  assign n66081 = n66097 & n66098;
  assign n66075 = ~n66105;
  assign n66083 = ~n66106;
  assign n66091 = n66115 ^ n66116;
  assign n66117 = ~n66115;
  assign n65876 = n65990 & n65991;
  assign n65980 = n66014 ^ n62837;
  assign n66002 = n66015 & n66016;
  assign n65996 = ~n66015;
  assign n65978 = ~n66027;
  assign n66009 = ~n66014;
  assign n66013 = n66038 ^ n66039;
  assign n66048 = n66022 & n4295;
  assign n66037 = ~n66022;
  assign n66060 = n66076 & n66077;
  assign n66074 = ~n66081;
  assign n66044 = n66083 & n66084;
  assign n62181 = n63447 ^ n66091;
  assign n66085 = ~n66091;
  assign n66107 = n66117 & n66118;
  assign n65964 = n65876 & n65915;
  assign n65965 = ~n65876;
  assign n61779 = n65979 ^ n65980;
  assign n65995 = n65996 & n65997;
  assign n65972 = ~n66002;
  assign n66004 = n66009 & n66010;
  assign n65920 = n66012 ^ n66013;
  assign n65946 = n66013 & n66024;
  assign n66029 = n66037 & n360;
  assign n66018 = ~n66048;
  assign n66049 = ~n66060;
  assign n66057 = n66044 & n66069;
  assign n66043 = n66074 & n66075;
  assign n66062 = ~n66044;
  assign n62211 = ~n62181;
  assign n66080 = n66085 & n63447;
  assign n66088 = ~n66107;
  assign n65916 = ~n65964;
  assign n65949 = n61779 & n64041;
  assign n65959 = n65965 & n65966;
  assign n61811 = ~n61779;
  assign n65967 = n65972 & n65928;
  assign n65956 = ~n65995;
  assign n65977 = ~n66004;
  assign n65987 = ~n66029;
  assign n66019 = n66043 ^ n66044;
  assign n66021 = n66049 & n66050;
  assign n66046 = ~n66057;
  assign n66052 = n62211 & n64745;
  assign n66047 = ~n66043;
  assign n66053 = n66062 & n66020;
  assign n66036 = ~n66080;
  assign n66063 = n66088 & n66089;
  assign n65922 = ~n65949;
  assign n65882 = ~n65959;
  assign n65941 = n61811 & n62853;
  assign n65955 = ~n65967;
  assign n65963 = n65956 & n65972;
  assign n65948 = n65977 & n65978;
  assign n65952 = n66019 ^ n66020;
  assign n65985 = n66021 ^ n66022;
  assign n66017 = ~n66021;
  assign n66028 = n66046 & n66047;
  assign n66035 = ~n66052;
  assign n66008 = ~n66053;
  assign n66030 = n66063 ^ n66064;
  assign n66058 = ~n66063;
  assign n65923 = ~n65941;
  assign n65921 = n65948 ^ n62769;
  assign n65914 = n65955 & n65956;
  assign n65929 = ~n65963;
  assign n65950 = n65948 & n62802;
  assign n65962 = ~n65948;
  assign n65947 = n360 ^ n65985;
  assign n65981 = n65952 & n375;
  assign n65984 = ~n65952;
  assign n65998 = n66017 & n66018;
  assign n66007 = ~n66028;
  assign n62108 = n63398 ^ n66030;
  assign n65983 = n66035 & n66036;
  assign n66026 = ~n66030;
  assign n66054 = n66058 & n66059;
  assign n65877 = n65914 ^ n65915;
  assign n61695 = n65920 ^ n65921;
  assign n65807 = n65922 & n65923;
  assign n65905 = n65928 ^ n65929;
  assign n65917 = ~n65914;
  assign n65817 = n65946 ^ n65947;
  assign n65932 = ~n65950;
  assign n65936 = n65962 & n62769;
  assign n65945 = ~n65947;
  assign n65927 = ~n65981;
  assign n65968 = n65984 & n4257;
  assign n65986 = ~n65998;
  assign n65982 = n66007 & n66008;
  assign n66003 = n65983 & n65954;
  assign n66005 = ~n65983;
  assign n62173 = ~n62108;
  assign n66023 = n66026 & n63398;
  assign n66033 = ~n66054;
  assign n65793 = n65876 ^ n65877;
  assign n65878 = n61695 & n63982;
  assign n65880 = n65807 & n65892;
  assign n65875 = ~n65807;
  assign n61713 = ~n61695;
  assign n65893 = n65905 & n16646;
  assign n65898 = n65916 & n65917;
  assign n65896 = ~n65905;
  assign n65919 = n65932 & n65920;
  assign n65910 = n65817 & n62698;
  assign n65895 = ~n65936;
  assign n65911 = ~n65817;
  assign n65883 = n65945 & n65946;
  assign n65957 = ~n65968;
  assign n65953 = n65982 ^ n65983;
  assign n65951 = n65986 & n65987;
  assign n65989 = ~n65982;
  assign n65988 = ~n66003;
  assign n65993 = n62173 & n64689;
  assign n65992 = n66005 & n66006;
  assign n65976 = ~n66023;
  assign n65999 = n66033 & n66034;
  assign n65840 = n65793 & n16551;
  assign n65841 = ~n65793;
  assign n65865 = n65875 & n65835;
  assign n65869 = n61713 & n62769;
  assign n65846 = ~n65878;
  assign n65843 = ~n65880;
  assign n65861 = ~n65893;
  assign n65879 = n65896 & n390;
  assign n65881 = ~n65898;
  assign n65820 = ~n65910;
  assign n65901 = n65911 & n62732;
  assign n65894 = ~n65919;
  assign n65887 = ~n65883;
  assign n65913 = n65951 ^ n65952;
  assign n65874 = n65953 ^ n65954;
  assign n65958 = ~n65951;
  assign n65969 = n65988 & n65989;
  assign n65961 = ~n65992;
  assign n65975 = ~n65993;
  assign n65971 = n65999 ^ n63369;
  assign n66000 = ~n65999;
  assign n65785 = ~n65840;
  assign n65827 = n65841 & n389;
  assign n65857 = n65861 & n65813;
  assign n65810 = ~n65865;
  assign n65845 = ~n65869;
  assign n65826 = ~n65879;
  assign n65834 = n65881 & n65882;
  assign n65860 = n65894 & n65895;
  assign n65859 = ~n65901;
  assign n65884 = n375 ^ n65913;
  assign n65912 = n65874 & n4218;
  assign n65918 = ~n65874;
  assign n65942 = n65957 & n65958;
  assign n65960 = ~n65969;
  assign n62100 = n65970 ^ n65971;
  assign n65888 = n65975 & n65976;
  assign n65994 = n66000 & n66001;
  assign n65753 = ~n65827;
  assign n65808 = n65834 ^ n65835;
  assign n65730 = n65845 & n65846;
  assign n65825 = ~n65857;
  assign n65818 = n65860 ^ n62698;
  assign n65847 = n65861 & n65826;
  assign n65844 = ~n65834;
  assign n65858 = ~n65860;
  assign n65740 = n65883 ^ n65884;
  assign n65886 = ~n65884;
  assign n65871 = ~n65912;
  assign n65904 = n65918 & n374;
  assign n65926 = ~n65942;
  assign n65944 = n62100 & n63384;
  assign n65943 = n65888 & n65909;
  assign n65908 = n65960 & n65961;
  assign n65934 = ~n65888;
  assign n62125 = ~n62100;
  assign n65973 = ~n65994;
  assign n65712 = n65807 ^ n65808;
  assign n61611 = n65817 ^ n65818;
  assign n65800 = n65730 & n65771;
  assign n65798 = ~n65730;
  assign n65792 = n65825 & n65826;
  assign n65824 = n65843 & n65844;
  assign n65814 = ~n65847;
  assign n65836 = n65858 & n65859;
  assign n65852 = n65740 & n62644;
  assign n65848 = ~n65740;
  assign n65811 = n65886 & n65887;
  assign n65854 = ~n65904;
  assign n65889 = n65908 ^ n65909;
  assign n65873 = n65926 & n65927;
  assign n65931 = n65934 & n65935;
  assign n65925 = ~n65908;
  assign n65930 = n62125 & n64653;
  assign n65924 = ~n65943;
  assign n65902 = ~n65944;
  assign n65937 = n65973 & n65974;
  assign n65769 = n65712 & n388;
  assign n65748 = n65792 ^ n65793;
  assign n65767 = ~n65712;
  assign n65781 = n61611 & n63959;
  assign n65794 = n65798 & n65799;
  assign n65763 = ~n65800;
  assign n61633 = ~n61611;
  assign n63887 = n65813 ^ n65814;
  assign n65786 = ~n65792;
  assign n65809 = ~n65824;
  assign n65819 = ~n65836;
  assign n65828 = n65848 & n62656;
  assign n65739 = ~n65852;
  assign n65842 = n65873 ^ n65874;
  assign n65802 = n65888 ^ n65889;
  assign n65872 = ~n65873;
  assign n65899 = n65924 & n65925;
  assign n65903 = ~n65930;
  assign n65891 = ~n65931;
  assign n65900 = n65937 ^ n65938;
  assign n65939 = ~n65937;
  assign n65714 = n389 ^ n65748;
  assign n65749 = n65767 & n16413;
  assign n65670 = ~n65769;
  assign n65765 = n61633 & n62698;
  assign n65743 = ~n65781;
  assign n65780 = n65785 & n65786;
  assign n65733 = ~n65794;
  assign n65719 = ~n63887;
  assign n65770 = n65809 & n65810;
  assign n65777 = n65819 & n65820;
  assign n65783 = ~n65828;
  assign n65812 = n374 ^ n65842;
  assign n65837 = n65802 & n4169;
  assign n65851 = ~n65802;
  assign n65870 = n65871 & n65872;
  assign n65890 = ~n65899;
  assign n62029 = n63321 ^ n65900;
  assign n65815 = n65902 & n65903;
  assign n65897 = n65900 & n63340;
  assign n65933 = n65939 & n65940;
  assign n63854 = n65714 ^ n63887;
  assign n65632 = n65714 & n65719;
  assign n65709 = ~n65749;
  assign n65742 = ~n65765;
  assign n65731 = n65770 ^ n65771;
  assign n65741 = n65777 ^ n62644;
  assign n65752 = ~n65780;
  assign n65764 = ~n65770;
  assign n65782 = ~n65777;
  assign n65654 = n65811 ^ n65812;
  assign n65728 = n65812 & n65811;
  assign n65803 = ~n65837;
  assign n65831 = n65851 & n373;
  assign n65853 = ~n65870;
  assign n65864 = n65815 & n65885;
  assign n65838 = n65890 & n65891;
  assign n62078 = ~n62029;
  assign n65868 = ~n65815;
  assign n65833 = ~n65897;
  assign n65906 = ~n65933;
  assign n65453 = ~n63854;
  assign n65637 = n65730 ^ n65731;
  assign n61528 = n65740 ^ n65741;
  assign n65647 = n65742 & n65743;
  assign n65711 = n65752 & n65753;
  assign n65750 = n65763 & n65764;
  assign n65772 = n65654 & n62603;
  assign n65773 = n65782 & n65783;
  assign n65766 = ~n65654;
  assign n65723 = ~n65728;
  assign n65759 = ~n65831;
  assign n65816 = n65838 ^ n65839;
  assign n65801 = n65853 & n65854;
  assign n65850 = ~n65864;
  assign n65849 = ~n65838;
  assign n65855 = n62078 & n64596;
  assign n65862 = n65868 & n65839;
  assign n65863 = n65906 & n65907;
  assign n65692 = n65637 & n16311;
  assign n65667 = n65711 ^ n65712;
  assign n65702 = n65647 & n65681;
  assign n65679 = ~n65637;
  assign n65698 = n61528 & n63899;
  assign n65700 = ~n65647;
  assign n61546 = ~n61528;
  assign n65710 = ~n65711;
  assign n65732 = ~n65750;
  assign n65754 = n65766 & n62588;
  assign n65660 = ~n65772;
  assign n65738 = ~n65773;
  assign n65762 = n65801 ^ n65802;
  assign n65725 = n65815 ^ n65816;
  assign n65804 = ~n65801;
  assign n65823 = n65849 & n65850;
  assign n65832 = ~n65855;
  assign n65806 = ~n65862;
  assign n65822 = n65863 ^ n63282;
  assign n65866 = ~n65863;
  assign n65633 = n388 ^ n65667;
  assign n65666 = n65679 & n387;
  assign n65628 = ~n65692;
  assign n65676 = n61546 & n62644;
  assign n65656 = ~n65698;
  assign n65677 = n65700 & n65701;
  assign n65663 = ~n65702;
  assign n65699 = n65709 & n65710;
  assign n65680 = n65732 & n65733;
  assign n65705 = n65738 & n65739;
  assign n65704 = ~n65754;
  assign n65729 = n373 ^ n65762;
  assign n65768 = n65725 & n372;
  assign n65776 = ~n65725;
  assign n65795 = n65803 & n65804;
  assign n61986 = n65821 ^ n65822;
  assign n65805 = ~n65823;
  assign n65720 = n65832 & n65833;
  assign n65856 = n65866 & n65867;
  assign n63815 = n65632 ^ n65633;
  assign n65634 = ~n65633;
  assign n65588 = ~n65666;
  assign n65657 = ~n65676;
  assign n65631 = ~n65677;
  assign n65648 = n65680 ^ n65681;
  assign n65669 = ~n65699;
  assign n65655 = n65705 ^ n62588;
  assign n65664 = ~n65680;
  assign n65703 = ~n65705;
  assign n65575 = n65728 ^ n65729;
  assign n65722 = ~n65729;
  assign n65691 = ~n65768;
  assign n65757 = n65776 & n4120;
  assign n65758 = ~n65795;
  assign n65774 = n65805 & n65806;
  assign n65788 = n61986 & n63282;
  assign n65787 = n65720 & n65775;
  assign n62021 = ~n61986;
  assign n65796 = ~n65720;
  assign n65829 = ~n65856;
  assign n65372 = ~n63815;
  assign n65553 = n65634 & n65632;
  assign n65542 = n65647 ^ n65648;
  assign n61451 = n65654 ^ n65655;
  assign n65551 = n65656 & n65657;
  assign n65658 = n65663 & n65664;
  assign n65636 = n65669 & n65670;
  assign n65685 = n65703 & n65704;
  assign n65678 = n65575 & n62539;
  assign n65684 = ~n65575;
  assign n65650 = n65722 & n65723;
  assign n65734 = ~n65757;
  assign n65724 = n65758 & n65759;
  assign n65721 = n65774 ^ n65775;
  assign n65761 = ~n65774;
  assign n65760 = ~n65787;
  assign n65756 = ~n65788;
  assign n65779 = n62021 & n64559;
  assign n65778 = n65796 & n65797;
  assign n65789 = n65829 & n65830;
  assign n65605 = n65542 & n16246;
  assign n65620 = n61451 & n62603;
  assign n65617 = n61451 & n65635;
  assign n65614 = n65551 & n65586;
  assign n65606 = ~n65542;
  assign n65580 = n65636 ^ n65637;
  assign n61499 = ~n61451;
  assign n65618 = ~n65551;
  assign n65629 = ~n65636;
  assign n65630 = ~n65658;
  assign n65616 = ~n65678;
  assign n65668 = n65684 & n62568;
  assign n65659 = ~n65685;
  assign n65653 = n65720 ^ n65721;
  assign n65693 = n65724 ^ n65725;
  assign n65735 = ~n65724;
  assign n65751 = n65760 & n65761;
  assign n65727 = ~n65778;
  assign n65755 = ~n65779;
  assign n65747 = n65789 ^ n63245;
  assign n65790 = ~n65789;
  assign n65554 = n387 ^ n65580;
  assign n65547 = ~n65605;
  assign n65589 = n65606 & n386;
  assign n65599 = n61499 & n63868;
  assign n65579 = ~n65614;
  assign n63938 = ~n65617;
  assign n65602 = n65618 & n65619;
  assign n65603 = n61499 & n63941;
  assign n65574 = ~n65620;
  assign n65613 = n65628 & n65629;
  assign n65585 = n65630 & n65631;
  assign n65612 = n65659 & n65660;
  assign n65572 = ~n65668;
  assign n65651 = n372 ^ n65693;
  assign n65686 = n65653 & n4067;
  assign n65689 = ~n65653;
  assign n65717 = n65734 & n65735;
  assign n61906 = n65746 ^ n65747;
  assign n65726 = ~n65751;
  assign n65688 = n65755 & n65756;
  assign n65784 = n65790 & n65791;
  assign n63800 = n65553 ^ n65554;
  assign n65461 = n65554 & n65553;
  assign n65552 = n65585 ^ n65586;
  assign n65505 = ~n65589;
  assign n65573 = ~n65599;
  assign n65546 = ~n65602;
  assign n63962 = ~n65603;
  assign n65576 = n65612 ^ n62539;
  assign n65587 = ~n65613;
  assign n65578 = ~n65585;
  assign n65615 = ~n65612;
  assign n65487 = n65650 ^ n65651;
  assign n65563 = n65651 & n65650;
  assign n65646 = ~n65686;
  assign n65671 = n65689 & n371;
  assign n65690 = ~n65717;
  assign n65687 = n65726 & n65727;
  assign n65716 = n61906 & n64527;
  assign n65715 = n65688 & n65736;
  assign n65713 = n61906 & n65737;
  assign n65718 = ~n65688;
  assign n61939 = ~n61906;
  assign n65744 = ~n65784;
  assign n65276 = ~n63800;
  assign n65469 = ~n65461;
  assign n65458 = n65551 ^ n65552;
  assign n65459 = n65573 & n65574;
  assign n61371 = n65575 ^ n65576;
  assign n65577 = n65578 & n65579;
  assign n65541 = n65587 & n65588;
  assign n65597 = n65487 & n62529;
  assign n65595 = n65615 & n65616;
  assign n65607 = ~n65487;
  assign n65609 = ~n65671;
  assign n65643 = n65687 ^ n65688;
  assign n65652 = n65690 & n65691;
  assign n65682 = ~n65687;
  assign n64610 = ~n65713;
  assign n65683 = ~n65715;
  assign n65696 = n61939 & n64586;
  assign n65673 = ~n65716;
  assign n65694 = n61939 & n63268;
  assign n65695 = n65718 & n65644;
  assign n65708 = n65744 & n65745;
  assign n65508 = n65458 & n16138;
  assign n65499 = ~n65458;
  assign n65503 = n65541 ^ n65542;
  assign n65527 = n61371 & n63831;
  assign n65532 = n65459 & n65555;
  assign n61405 = ~n61371;
  assign n65533 = ~n65459;
  assign n65548 = ~n65541;
  assign n65545 = ~n65577;
  assign n65571 = ~n65595;
  assign n65535 = ~n65597;
  assign n65581 = n65607 & n62495;
  assign n65560 = n65643 ^ n65644;
  assign n65604 = n65652 ^ n65653;
  assign n65645 = ~n65652;
  assign n65665 = n65682 & n65683;
  assign n65672 = ~n65694;
  assign n65642 = ~n65695;
  assign n64591 = ~n65696;
  assign n65675 = n65708 ^ n63194;
  assign n65706 = ~n65708;
  assign n65486 = n65499 & n385;
  assign n65462 = n386 ^ n65503;
  assign n65466 = ~n65508;
  assign n65490 = ~n65527;
  assign n65517 = n61405 & n62568;
  assign n65507 = ~n65532;
  assign n65516 = n65533 & n65502;
  assign n65501 = n65545 & n65546;
  assign n65536 = n65547 & n65548;
  assign n65528 = n65571 & n65572;
  assign n65492 = ~n65581;
  assign n65564 = n371 ^ n65604;
  assign n65596 = n65560 & n370;
  assign n65598 = ~n65560;
  assign n65624 = n65645 & n65646;
  assign n65641 = ~n65665;
  assign n65566 = n65672 & n65673;
  assign n61831 = n65674 ^ n65675;
  assign n65697 = n65706 & n65707;
  assign n63735 = n65461 ^ n65462;
  assign n65406 = ~n65486;
  assign n65468 = ~n65462;
  assign n65460 = n65501 ^ n65502;
  assign n65456 = ~n65516;
  assign n65489 = ~n65517;
  assign n65488 = n65528 ^ n62495;
  assign n65506 = ~n65501;
  assign n65504 = ~n65536;
  assign n65534 = ~n65528;
  assign n65403 = n65563 ^ n65564;
  assign n65565 = ~n65564;
  assign n65523 = ~n65596;
  assign n65582 = n65598 & n4032;
  assign n65608 = ~n65624;
  assign n65600 = n65641 & n65642;
  assign n65627 = n65566 & n65649;
  assign n65638 = n61831 & n64471;
  assign n65640 = ~n65566;
  assign n61873 = ~n61831;
  assign n65661 = ~n65697;
  assign n65197 = ~n63735;
  assign n65375 = n65459 ^ n65460;
  assign n65376 = n65468 & n65469;
  assign n61289 = n65487 ^ n65488;
  assign n65363 = n65489 & n65490;
  assign n65457 = n65504 & n65505;
  assign n65485 = n65506 & n65507;
  assign n65518 = n65534 & n65535;
  assign n65525 = n65403 & n62481;
  assign n65524 = ~n65403;
  assign n65478 = n65565 & n65563;
  assign n65561 = ~n65582;
  assign n65567 = n65600 ^ n65601;
  assign n65559 = n65608 & n65609;
  assign n65611 = ~n65627;
  assign n65622 = n61873 & n63194;
  assign n65610 = ~n65600;
  assign n65592 = ~n65638;
  assign n65623 = n65640 & n65601;
  assign n65639 = n65661 & n65662;
  assign n65413 = n65375 & n384;
  assign n65412 = ~n65375;
  assign n65390 = ~n65376;
  assign n65440 = n61289 & n65453;
  assign n65441 = n61289 & n62495;
  assign n65439 = n65363 & n65454;
  assign n65411 = n65457 ^ n65458;
  assign n65446 = ~n65363;
  assign n61341 = ~n61289;
  assign n65455 = ~n65485;
  assign n65467 = ~n65457;
  assign n65491 = ~n65518;
  assign n65498 = n65524 & n62458;
  assign n65397 = ~n65525;
  assign n65477 = ~n65478;
  assign n65520 = n65559 ^ n65560;
  assign n65475 = n65566 ^ n65567;
  assign n65562 = ~n65559;
  assign n65594 = n65610 & n65611;
  assign n65593 = ~n65622;
  assign n65570 = ~n65623;
  assign n65584 = n65639 ^ n63129;
  assign n65625 = ~n65639;
  assign n65377 = n385 ^ n65411;
  assign n65398 = n65412 & n16072;
  assign n65319 = ~n65413;
  assign n65410 = ~n65439;
  assign n63852 = ~n65440;
  assign n65400 = ~n65441;
  assign n65423 = n65446 & n65408;
  assign n65424 = n61341 & n63795;
  assign n65425 = n61341 & n63854;
  assign n65407 = n65455 & n65456;
  assign n65449 = n65466 & n65467;
  assign n65445 = n65491 & n65492;
  assign n65443 = ~n65498;
  assign n65479 = n370 ^ n65520;
  assign n65521 = n65475 & n369;
  assign n65519 = ~n65475;
  assign n65557 = n65561 & n65562;
  assign n61781 = n65583 ^ n65584;
  assign n65513 = n65592 & n65593;
  assign n65569 = ~n65594;
  assign n65621 = n65625 & n65626;
  assign n63697 = n65376 ^ n65377;
  assign n65289 = n65377 & n65390;
  assign n65371 = ~n65398;
  assign n65364 = n65407 ^ n65408;
  assign n65379 = ~n65423;
  assign n65401 = ~n65424;
  assign n63871 = ~n65425;
  assign n65409 = ~n65407;
  assign n65404 = n65445 ^ n62458;
  assign n65405 = ~n65449;
  assign n65444 = ~n65445;
  assign n65314 = n65478 ^ n65479;
  assign n65476 = ~n65479;
  assign n65511 = n65519 & n3990;
  assign n65435 = ~n65521;
  assign n65522 = ~n65557;
  assign n65544 = n61781 & n65558;
  assign n65543 = n61781 & n64457;
  assign n65539 = n65513 & n65568;
  assign n65512 = n65569 & n65570;
  assign n65540 = ~n65513;
  assign n61762 = ~n61781;
  assign n65590 = ~n65621;
  assign n65124 = ~n63697;
  assign n65284 = n65363 ^ n65364;
  assign n65287 = n65400 & n65401;
  assign n61233 = n65403 ^ n65404;
  assign n65374 = n65405 & n65406;
  assign n65402 = n65409 & n65410;
  assign n65437 = n65443 & n65444;
  assign n65436 = n65314 & n62443;
  assign n65432 = ~n65314;
  assign n65384 = n65476 & n65477;
  assign n65484 = ~n65511;
  assign n65472 = n65512 ^ n65513;
  assign n65474 = n65522 & n65523;
  assign n65515 = ~n65539;
  assign n65529 = n65540 & n65473;
  assign n65510 = ~n65543;
  assign n64525 = ~n65544;
  assign n65514 = ~n65512;
  assign n65530 = n61762 & n65556;
  assign n65531 = n61762 & n63166;
  assign n65537 = n65590 & n65591;
  assign n65323 = n65284 & n399;
  assign n65324 = ~n65284;
  assign n65360 = n61233 & n62481;
  assign n65359 = n61233 & n65372;
  assign n65361 = n65287 & n65373;
  assign n65320 = n65374 ^ n65375;
  assign n61268 = ~n61233;
  assign n65353 = ~n65287;
  assign n65370 = ~n65374;
  assign n65378 = ~n65402;
  assign n65414 = n65432 & n62425;
  assign n65317 = ~n65436;
  assign n65396 = ~n65437;
  assign n65399 = ~n65384;
  assign n65387 = n65472 ^ n65473;
  assign n65426 = n65474 ^ n65475;
  assign n65483 = ~n65474;
  assign n65500 = n65514 & n65515;
  assign n65481 = ~n65529;
  assign n64498 = ~n65530;
  assign n65509 = ~n65531;
  assign n65496 = n65537 ^ n65538;
  assign n65549 = ~n65537;
  assign n65290 = n384 ^ n65320;
  assign n65238 = ~n65323;
  assign n65310 = n65324 & n15958;
  assign n65347 = n65353 & n65328;
  assign n65345 = n61268 & n63756;
  assign n63818 = ~n65359;
  assign n65346 = n61268 & n63815;
  assign n65312 = ~n65360;
  assign n65334 = ~n65361;
  assign n65362 = n65370 & n65371;
  assign n65327 = n65378 & n65379;
  assign n65354 = n65396 & n65397;
  assign n65358 = ~n65414;
  assign n65385 = n369 ^ n65426;
  assign n65433 = n65387 & n368;
  assign n65427 = ~n65387;
  assign n65471 = n65483 & n65484;
  assign n64520 = n64498 & n64525;
  assign n61660 = n63091 ^ n65496;
  assign n65480 = ~n65500;
  assign n65429 = n65509 & n65510;
  assign n65497 = ~n65496;
  assign n65526 = n65549 & n65550;
  assign n63658 = n65289 ^ n65290;
  assign n65286 = ~n65310;
  assign n65291 = ~n65290;
  assign n65288 = n65327 ^ n65328;
  assign n65311 = ~n65345;
  assign n63836 = ~n65346;
  assign n65293 = ~n65347;
  assign n65315 = n65354 ^ n62425;
  assign n65333 = ~n65327;
  assign n65318 = ~n65362;
  assign n65357 = ~n65354;
  assign n65225 = n65384 ^ n65385;
  assign n65304 = n65385 & n65399;
  assign n65417 = n65427 & n3965;
  assign n65350 = ~n65433;
  assign n65434 = ~n65471;
  assign n65428 = n65480 & n65481;
  assign n65450 = n65429 & n65482;
  assign n65463 = n61660 & n64461;
  assign n61742 = ~n61660;
  assign n65451 = ~n65429;
  assign n65493 = n65497 & n63091;
  assign n65494 = ~n65526;
  assign n65014 = ~n63658;
  assign n65192 = n65287 ^ n65288;
  assign n65201 = n65291 & n65289;
  assign n65193 = n65311 & n65312;
  assign n61156 = n65314 ^ n65315;
  assign n65283 = n65318 & n65319;
  assign n65313 = n65333 & n65334;
  assign n65336 = n65357 & n65358;
  assign n65337 = n65225 & n62383;
  assign n65348 = ~n65225;
  assign n65309 = ~n65304;
  assign n65392 = ~n65417;
  assign n65388 = n65428 ^ n65429;
  assign n65386 = n65434 & n65435;
  assign n65431 = ~n65450;
  assign n65448 = n65451 & n65389;
  assign n65438 = n61742 & n64361;
  assign n64455 = ~n65463;
  assign n65442 = n61742 & n65470;
  assign n65430 = ~n65428;
  assign n65416 = ~n65493;
  assign n65452 = n65494 & n65495;
  assign n65230 = n65192 & n398;
  assign n65235 = ~n65192;
  assign n65218 = ~n65201;
  assign n65269 = n61156 & n62443;
  assign n65236 = n65283 ^ n65284;
  assign n65270 = n61156 & n63800;
  assign n65272 = n65193 & n65240;
  assign n61173 = ~n61156;
  assign n65267 = ~n65193;
  assign n65292 = ~n65313;
  assign n65285 = ~n65283;
  assign n65316 = ~n65336;
  assign n65228 = ~n65337;
  assign n65335 = n65348 & n62389;
  assign n65338 = n65386 ^ n65387;
  assign n65299 = n65388 ^ n65389;
  assign n65391 = ~n65386;
  assign n65418 = n65430 & n65431;
  assign n65415 = ~n65438;
  assign n64486 = ~n65442;
  assign n65395 = ~n65448;
  assign n65422 = n65452 ^ n63047;
  assign n65464 = ~n65452;
  assign n65156 = ~n65230;
  assign n65229 = n65235 & n15897;
  assign n65202 = n399 ^ n65236;
  assign n65255 = n65267 & n65268;
  assign n65221 = ~n65269;
  assign n63775 = ~n65270;
  assign n65262 = n61173 & n63728;
  assign n65247 = ~n65272;
  assign n65257 = n61173 & n65276;
  assign n65263 = n65285 & n65286;
  assign n65239 = n65292 & n65293;
  assign n65266 = n65316 & n65317;
  assign n65274 = ~n65335;
  assign n65305 = n368 ^ n65338;
  assign n65339 = n65299 & n383;
  assign n65344 = ~n65299;
  assign n65365 = n65391 & n65392;
  assign n65343 = n65415 & n65416;
  assign n65394 = ~n65418;
  assign n61575 = n65421 ^ n65422;
  assign n65447 = n65464 & n65465;
  assign n63616 = n65201 ^ n65202;
  assign n65118 = n65202 & n65218;
  assign n65190 = ~n65229;
  assign n65194 = n65239 ^ n65240;
  assign n65199 = ~n65255;
  assign n63797 = ~n65257;
  assign n65222 = ~n65262;
  assign n65237 = ~n65263;
  assign n65226 = n65266 ^ n62389;
  assign n65246 = ~n65239;
  assign n65140 = n65304 ^ n65305;
  assign n65275 = ~n65266;
  assign n65308 = ~n65305;
  assign n65261 = ~n65339;
  assign n65321 = n65344 & n3911;
  assign n65349 = ~n65365;
  assign n65382 = n65343 & n65307;
  assign n65366 = n61575 & n65393;
  assign n65367 = n61575 & n63065;
  assign n65342 = n65394 & n65395;
  assign n65380 = ~n65343;
  assign n61662 = ~n61575;
  assign n65419 = ~n65447;
  assign n64918 = ~n63616;
  assign n65115 = n65193 ^ n65194;
  assign n65104 = ~n65118;
  assign n65116 = n65221 & n65222;
  assign n61084 = n65225 ^ n65226;
  assign n65191 = n65237 & n65238;
  assign n65223 = n65246 & n65247;
  assign n65254 = n65140 & n62359;
  assign n65256 = n65274 & n65275;
  assign n65248 = ~n65140;
  assign n65211 = n65308 & n65309;
  assign n65303 = ~n65321;
  assign n65306 = n65342 ^ n65343;
  assign n65298 = n65349 & n65350;
  assign n64427 = ~n65366;
  assign n65331 = ~n65367;
  assign n65351 = n61662 & n64340;
  assign n65356 = n61662 & n64417;
  assign n65355 = n65380 & n65381;
  assign n65340 = ~n65382;
  assign n65341 = ~n65342;
  assign n65383 = n65419 & n65420;
  assign n65160 = n65115 & n15813;
  assign n65152 = ~n65115;
  assign n65157 = n65191 ^ n65192;
  assign n65184 = n61084 & n65197;
  assign n65185 = n61084 & n62383;
  assign n65187 = n65116 & n65162;
  assign n65182 = ~n65116;
  assign n61123 = ~n61084;
  assign n65198 = ~n65223;
  assign n65189 = ~n65191;
  assign n65234 = n65248 & n62332;
  assign n65143 = ~n65254;
  assign n65227 = ~n65256;
  assign n65224 = ~n65211;
  assign n65253 = n65298 ^ n65299;
  assign n65210 = n65306 ^ n65307;
  assign n65302 = ~n65298;
  assign n65322 = n65340 & n65341;
  assign n65332 = ~n65351;
  assign n65301 = ~n65355;
  assign n64438 = ~n65356;
  assign n65326 = n65383 ^ n62972;
  assign n65368 = ~n65383;
  assign n65139 = n65152 & n397;
  assign n65119 = n398 ^ n65157;
  assign n65121 = ~n65160;
  assign n65165 = n61123 & n63735;
  assign n65172 = n61123 & n63655;
  assign n65173 = n65182 & n65183;
  assign n63738 = ~n65184;
  assign n65145 = ~n65185;
  assign n65153 = ~n65187;
  assign n65178 = n65189 & n65190;
  assign n65161 = n65198 & n65199;
  assign n65181 = n65227 & n65228;
  assign n65180 = ~n65234;
  assign n65212 = n383 ^ n65253;
  assign n65252 = n65210 & n3849;
  assign n65249 = ~n65210;
  assign n65277 = n65302 & n65303;
  assign n65300 = ~n65322;
  assign n61491 = n65325 ^ n65326;
  assign n65251 = n65331 & n65332;
  assign n65352 = n65368 & n65369;
  assign n63578 = n65118 ^ n65119;
  assign n65103 = ~n65119;
  assign n65058 = ~n65139;
  assign n65117 = n65161 ^ n65162;
  assign n63761 = ~n65165;
  assign n65144 = ~n65172;
  assign n65113 = ~n65173;
  assign n65154 = ~n65161;
  assign n65155 = ~n65178;
  assign n65141 = n65181 ^ n62332;
  assign n65052 = n65211 ^ n65212;
  assign n65179 = ~n65181;
  assign n65133 = n65212 & n65224;
  assign n65241 = n65249 & n382;
  assign n65217 = ~n65252;
  assign n65260 = ~n65277;
  assign n65279 = n61491 & n64378;
  assign n65250 = n65300 & n65301;
  assign n65294 = n65251 & n65215;
  assign n65295 = n61491 & n62972;
  assign n65281 = ~n65251;
  assign n61581 = ~n61491;
  assign n65329 = ~n65352;
  assign n64864 = ~n63578;
  assign n65036 = n65103 & n65104;
  assign n65033 = n65116 ^ n65117;
  assign n61048 = n65140 ^ n65141;
  assign n65028 = n65144 & n65145;
  assign n65137 = n65153 & n65154;
  assign n65114 = n65155 & n65156;
  assign n65166 = n65179 & n65180;
  assign n65138 = ~n65133;
  assign n65164 = ~n65241;
  assign n65214 = n65250 ^ n65251;
  assign n65209 = n65260 & n65261;
  assign n64389 = ~n65279;
  assign n65258 = ~n65250;
  assign n65273 = n61581 & n65280;
  assign n65265 = n65281 & n65282;
  assign n65271 = n61581 & n64320;
  assign n65259 = ~n65294;
  assign n65242 = ~n65295;
  assign n65278 = n65329 & n65330;
  assign n65075 = n65033 & n15732;
  assign n65059 = ~n65033;
  assign n65102 = n61048 & n62359;
  assign n65069 = n65114 ^ n65115;
  assign n65100 = n61048 & n65124;
  assign n65093 = n65028 & n65125;
  assign n61075 = ~n61048;
  assign n65092 = ~n65028;
  assign n65120 = ~n65114;
  assign n65112 = ~n65137;
  assign n65142 = ~n65166;
  assign n65167 = n65209 ^ n65210;
  assign n65132 = n65214 ^ n65215;
  assign n65216 = ~n65209;
  assign n65231 = n65258 & n65259;
  assign n65220 = ~n65265;
  assign n65243 = ~n65271;
  assign n64403 = ~n65273;
  assign n65233 = n65278 ^ n62897;
  assign n65296 = ~n65278;
  assign n65054 = n65059 & n396;
  assign n65037 = n397 ^ n65069;
  assign n65034 = ~n65075;
  assign n65086 = n65092 & n65061;
  assign n65067 = ~n65093;
  assign n65090 = n61075 & n63613;
  assign n63704 = ~n65100;
  assign n65085 = n61075 & n63697;
  assign n65056 = ~n65102;
  assign n65060 = n65112 & n65113;
  assign n65091 = n65120 & n65121;
  assign n65101 = n65142 & n65143;
  assign n65134 = n382 ^ n65167;
  assign n65170 = n65132 & n3787;
  assign n65171 = ~n65132;
  assign n65196 = n65216 & n65217;
  assign n65219 = ~n65231;
  assign n61410 = n65232 ^ n65233;
  assign n65169 = n65242 & n65243;
  assign n65264 = n65296 & n65297;
  assign n63554 = n65036 ^ n65037;
  assign n64952 = n65037 & n65036;
  assign n64984 = ~n65054;
  assign n65029 = n65060 ^ n65061;
  assign n63718 = ~n65085;
  assign n65031 = ~n65086;
  assign n65055 = ~n65090;
  assign n65057 = ~n65091;
  assign n65068 = ~n65060;
  assign n65053 = n65101 ^ n62297;
  assign n65094 = n65101 & n62323;
  assign n65099 = ~n65101;
  assign n64958 = n65133 ^ n65134;
  assign n65048 = n65134 & n65138;
  assign n65126 = ~n65170;
  assign n65149 = n65171 & n381;
  assign n65163 = ~n65196;
  assign n65208 = n61410 & n64287;
  assign n65200 = n61410 & n65213;
  assign n65203 = n65169 & n65136;
  assign n65168 = n65219 & n65220;
  assign n65206 = ~n65169;
  assign n61470 = ~n61410;
  assign n65244 = ~n65264;
  assign n64790 = ~n63554;
  assign n64950 = n65028 ^ n65029;
  assign n60991 = n65052 ^ n65053;
  assign n64954 = n65055 & n65056;
  assign n65032 = n65057 & n65058;
  assign n65050 = n65067 & n65068;
  assign n65066 = ~n65094;
  assign n65078 = n65099 & n62297;
  assign n65079 = n64958 & n62286;
  assign n65087 = ~n64958;
  assign n65081 = ~n65149;
  assign n65131 = n65163 & n65164;
  assign n65135 = n65168 ^ n65169;
  assign n65174 = ~n65168;
  assign n65177 = n61470 & n62897;
  assign n64358 = ~n65200;
  assign n65175 = ~n65203;
  assign n65176 = n65206 & n65207;
  assign n65159 = ~n65208;
  assign n65188 = n61470 & n64345;
  assign n65195 = n65244 & n65245;
  assign n64977 = n64950 & n395;
  assign n64988 = ~n64950;
  assign n65019 = n60991 & n63591;
  assign n65010 = n64954 & n64979;
  assign n64991 = n65032 ^ n65033;
  assign n65015 = n60991 & n63658;
  assign n65012 = ~n64954;
  assign n61017 = ~n60991;
  assign n65030 = ~n65050;
  assign n65035 = ~n65032;
  assign n65051 = n65066 & n65052;
  assign n65022 = ~n65078;
  assign n64990 = ~n65079;
  assign n65062 = n65087 & n62258;
  assign n65088 = n65131 ^ n65132;
  assign n65041 = n65135 ^ n65136;
  assign n65127 = ~n65131;
  assign n65148 = n65174 & n65175;
  assign n65130 = ~n65176;
  assign n65158 = ~n65177;
  assign n64348 = ~n65188;
  assign n65147 = n65195 ^ n62820;
  assign n65204 = ~n65195;
  assign n64913 = ~n64977;
  assign n64972 = n64988 & n15662;
  assign n64953 = n396 ^ n64991;
  assign n64981 = ~n65010;
  assign n65002 = n65012 & n65013;
  assign n64996 = n61017 & n65014;
  assign n65003 = n61017 & n62297;
  assign n63679 = ~n65015;
  assign n64975 = ~n65019;
  assign n64978 = n65030 & n65031;
  assign n65011 = n65034 & n65035;
  assign n65021 = ~n65051;
  assign n64946 = ~n65062;
  assign n65049 = n381 ^ n65088;
  assign n65089 = n65041 & n3736;
  assign n65082 = ~n65041;
  assign n65111 = n65126 & n65127;
  assign n61336 = n65146 ^ n65147;
  assign n65129 = ~n65148;
  assign n65044 = n65158 & n65159;
  assign n65186 = n65204 & n65205;
  assign n63494 = n64952 ^ n64953;
  assign n64883 = n64953 & n64952;
  assign n64957 = ~n64972;
  assign n64955 = n64978 ^ n64979;
  assign n63661 = ~n64996;
  assign n64948 = ~n65002;
  assign n64976 = ~n65003;
  assign n64983 = ~n65011;
  assign n64980 = ~n64978;
  assign n64995 = n65021 & n65022;
  assign n64885 = n65048 ^ n65049;
  assign n64966 = n65049 & n65048;
  assign n65070 = n65082 & n380;
  assign n65043 = ~n65089;
  assign n65080 = ~n65111;
  assign n65123 = n65044 & n65128;
  assign n65083 = n65129 & n65130;
  assign n65105 = n61336 & n64307;
  assign n65107 = n61336 & n64212;
  assign n65122 = ~n65044;
  assign n61415 = ~n61336;
  assign n65150 = ~n65186;
  assign n64739 = ~n63494;
  assign n64899 = ~n64883;
  assign n64869 = n64954 ^ n64955;
  assign n64880 = n64975 & n64976;
  assign n64973 = n64980 & n64981;
  assign n64949 = n64983 & n64984;
  assign n64959 = n64995 ^ n62258;
  assign n64989 = ~n64995;
  assign n64998 = n64885 & n62203;
  assign n64997 = ~n64885;
  assign n64969 = ~n64966;
  assign n65001 = ~n65070;
  assign n65040 = n65080 & n65081;
  assign n65045 = n65083 ^ n65084;
  assign n65076 = ~n65083;
  assign n64318 = ~n65105;
  assign n65064 = ~n65107;
  assign n65097 = n61415 & n62820;
  assign n65095 = n61415 & n65110;
  assign n65098 = n65122 & n65084;
  assign n65077 = ~n65123;
  assign n65106 = n65150 & n65151;
  assign n64916 = n64869 & n15572;
  assign n64917 = ~n64869;
  assign n64936 = n64880 & n64944;
  assign n64911 = n64949 ^ n64950;
  assign n60937 = n64958 ^ n64959;
  assign n64934 = ~n64880;
  assign n64947 = ~n64973;
  assign n64956 = ~n64949;
  assign n64974 = n64989 & n64990;
  assign n64982 = n64997 & n62250;
  assign n64873 = ~n64998;
  assign n64999 = n65040 ^ n65041;
  assign n64965 = n65044 ^ n65045;
  assign n65042 = ~n65040;
  assign n65063 = n65076 & n65077;
  assign n64298 = ~n65095;
  assign n65065 = ~n65097;
  assign n65047 = ~n65098;
  assign n65072 = n65106 ^ n62749;
  assign n65108 = ~n65106;
  assign n64884 = n395 ^ n64911;
  assign n64870 = ~n64916;
  assign n64904 = n64917 & n394;
  assign n64907 = n60937 & n63616;
  assign n64923 = n60937 & n62258;
  assign n64929 = n64934 & n64906;
  assign n60980 = ~n60937;
  assign n64915 = ~n64936;
  assign n64905 = n64947 & n64948;
  assign n64938 = n64956 & n64957;
  assign n64945 = ~n64974;
  assign n64920 = ~n64982;
  assign n64967 = n380 ^ n64999;
  assign n65005 = n64965 & n379;
  assign n65004 = ~n64965;
  assign n65027 = n65042 & n65043;
  assign n65046 = ~n65063;
  assign n64962 = n65064 & n65065;
  assign n61264 = n65071 ^ n65072;
  assign n65096 = n65108 & n65109;
  assign n63457 = n64883 ^ n64884;
  assign n64815 = n64884 & n64899;
  assign n64854 = ~n64904;
  assign n64881 = n64905 ^ n64906;
  assign n63619 = ~n64907;
  assign n64901 = n60980 & n63556;
  assign n64900 = n60980 & n64918;
  assign n64876 = ~n64923;
  assign n64879 = ~n64929;
  assign n64914 = ~n64905;
  assign n64912 = ~n64938;
  assign n64908 = n64945 & n64946;
  assign n64810 = n64966 ^ n64967;
  assign n64968 = ~n64967;
  assign n64987 = n65004 & n3634;
  assign n64931 = ~n65005;
  assign n65000 = ~n65027;
  assign n65039 = n61264 & n64168;
  assign n65026 = n64962 & n65009;
  assign n65038 = n61264 & n64259;
  assign n65008 = n65046 & n65047;
  assign n65023 = ~n64962;
  assign n61322 = ~n61264;
  assign n65073 = ~n65096;
  assign n64696 = ~n63457;
  assign n64831 = ~n64815;
  assign n64820 = n64880 ^ n64881;
  assign n63636 = ~n64900;
  assign n64877 = ~n64901;
  assign n64886 = n64908 ^ n62203;
  assign n64868 = n64912 & n64913;
  assign n64902 = n64914 & n64915;
  assign n64919 = ~n64908;
  assign n64835 = ~n64810;
  assign n64897 = n64968 & n64969;
  assign n64971 = ~n64987;
  assign n64964 = n65000 & n65001;
  assign n64963 = n65008 ^ n65009;
  assign n65016 = n65023 & n65024;
  assign n65017 = n61322 & n65025;
  assign n65018 = n61322 & n62751;
  assign n65007 = ~n65026;
  assign n65006 = ~n65008;
  assign n64281 = ~n65038;
  assign n64986 = ~n65039;
  assign n65020 = n65073 & n65074;
  assign n64849 = n64820 & n393;
  assign n64846 = ~n64820;
  assign n64852 = n64868 ^ n64869;
  assign n64821 = n64876 & n64877;
  assign n60902 = n64885 ^ n64886;
  assign n64871 = ~n64868;
  assign n64878 = ~n64902;
  assign n64903 = n64919 & n64920;
  assign n64888 = ~n64897;
  assign n64896 = n64962 ^ n64963;
  assign n64924 = n64964 ^ n64965;
  assign n64970 = ~n64964;
  assign n64994 = n65006 & n65007;
  assign n64961 = ~n65016;
  assign n64257 = ~n65017;
  assign n64985 = ~n65018;
  assign n64993 = n65020 ^ n62754;
  assign n64836 = n64846 & n15529;
  assign n64788 = ~n64849;
  assign n64816 = n394 ^ n64852;
  assign n64848 = n60902 & n64864;
  assign n64847 = n60902 & n63479;
  assign n64844 = n64821 & n64865;
  assign n64850 = ~n64821;
  assign n60888 = ~n60902;
  assign n64867 = n64870 & n64871;
  assign n64856 = n64878 & n64879;
  assign n64872 = ~n64903;
  assign n64898 = n379 ^ n64924;
  assign n64925 = n64896 & n3578;
  assign n64926 = ~n64896;
  assign n64940 = n64970 & n64971;
  assign n64893 = n64985 & n64986;
  assign n61293 = n64992 ^ n64993;
  assign n64960 = ~n64994;
  assign n63406 = n64815 ^ n64816;
  assign n64760 = n64816 & n64831;
  assign n64817 = ~n64836;
  assign n64823 = ~n64844;
  assign n64808 = ~n64847;
  assign n63595 = ~n64848;
  assign n64840 = n64850 & n64851;
  assign n64838 = n60888 & n62203;
  assign n64837 = n60888 & n63578;
  assign n64822 = n64856 ^ n64851;
  assign n64824 = ~n64856;
  assign n64853 = ~n64867;
  assign n64845 = n64872 & n64873;
  assign n64748 = n64897 ^ n64898;
  assign n64887 = ~n64898;
  assign n64890 = ~n64925;
  assign n64921 = n64926 & n378;
  assign n64242 = n64939 ^ n61293;
  assign n64930 = ~n64940;
  assign n64927 = n64960 & n64961;
  assign n64951 = n61293 & n62754;
  assign n64943 = n64893 & n64928;
  assign n62824 = ~n61293;
  assign n64941 = ~n64893;
  assign n64654 = ~n63406;
  assign n64770 = n64821 ^ n64822;
  assign n64814 = n64823 & n64824;
  assign n63580 = ~n64837;
  assign n64809 = ~n64838;
  assign n64804 = ~n64840;
  assign n64811 = n64845 ^ n62181;
  assign n64819 = n64853 & n64854;
  assign n64841 = n64845 & n62211;
  assign n64858 = n64748 & n62108;
  assign n64855 = ~n64845;
  assign n64857 = ~n64748;
  assign n64829 = n64887 & n64888;
  assign n64861 = ~n64921;
  assign n64894 = n64927 ^ n64928;
  assign n64895 = n64930 & n64931;
  assign n64935 = n64941 & n64942;
  assign n64933 = ~n64943;
  assign n64910 = ~n64951;
  assign n64937 = n62824 & n64171;
  assign n64932 = ~n64927;
  assign n64791 = n64770 & n392;
  assign n64789 = ~n64770;
  assign n64781 = n64808 & n64809;
  assign n60780 = n64810 ^ n64811;
  assign n64803 = ~n64814;
  assign n64794 = n64819 ^ n64820;
  assign n64818 = ~n64819;
  assign n64834 = ~n64841;
  assign n64839 = n64855 & n62181;
  assign n64842 = n64857 & n62173;
  assign n64751 = ~n64858;
  assign n64826 = n64893 ^ n64894;
  assign n64862 = n64895 ^ n64896;
  assign n64889 = ~n64895;
  assign n64922 = n64932 & n64933;
  assign n64892 = ~n64935;
  assign n64909 = ~n64937;
  assign n64785 = n64789 & n15486;
  assign n64743 = ~n64791;
  assign n64761 = n393 ^ n64794;
  assign n64780 = n64803 & n64804;
  assign n64796 = n64781 & n64755;
  assign n64795 = n60780 & n63554;
  assign n64797 = n60780 & n62181;
  assign n60851 = ~n60780;
  assign n64792 = ~n64781;
  assign n64807 = n64817 & n64818;
  assign n64812 = n64834 & n64835;
  assign n64802 = ~n64839;
  assign n64772 = ~n64842;
  assign n64830 = n378 ^ n64862;
  assign n64859 = n64826 & n3502;
  assign n64863 = ~n64826;
  assign n64882 = n64889 & n64890;
  assign n64874 = n64909 & n64910;
  assign n64891 = ~n64922;
  assign n63374 = n64760 ^ n64761;
  assign n64754 = n64780 ^ n64781;
  assign n64766 = ~n64761;
  assign n64762 = ~n64785;
  assign n64783 = n60851 & n63447;
  assign n64782 = n60851 & n64790;
  assign n64784 = n64792 & n64793;
  assign n63535 = ~n64795;
  assign n64778 = ~n64796;
  assign n64768 = ~n64797;
  assign n64779 = ~n64780;
  assign n64787 = ~n64807;
  assign n64801 = ~n64812;
  assign n64710 = n64829 ^ n64830;
  assign n64774 = n64830 & n64829;
  assign n64828 = ~n64859;
  assign n64843 = n64863 & n377;
  assign n64833 = n64874 ^ n64875;
  assign n64860 = ~n64882;
  assign n64866 = n64891 & n64892;
  assign n64717 = n64754 ^ n64755;
  assign n64616 = ~n63374;
  assign n64715 = n64766 & n64760;
  assign n64764 = n64778 & n64779;
  assign n63558 = ~n64782;
  assign n64767 = ~n64783;
  assign n64757 = ~n64784;
  assign n64769 = n64787 & n64788;
  assign n64773 = n64801 & n64802;
  assign n64806 = n64710 & n62100;
  assign n64805 = ~n64710;
  assign n64800 = ~n64843;
  assign n64825 = n64860 & n64861;
  assign n64832 = n376 ^ n64866;
  assign n64737 = n64717 & n15473;
  assign n64725 = ~n64717;
  assign n64756 = ~n64764;
  assign n64727 = n64767 & n64768;
  assign n64741 = n64769 ^ n64770;
  assign n64749 = n64773 ^ n62108;
  assign n64763 = ~n64769;
  assign n64771 = ~n64773;
  assign n64786 = n64805 & n62125;
  assign n64702 = ~n64806;
  assign n64798 = n64825 ^ n64826;
  assign n64777 = n64832 ^ n64833;
  assign n64827 = ~n64825;
  assign n64724 = n64725 & n407;
  assign n64712 = ~n64737;
  assign n64723 = n392 ^ n64741;
  assign n60730 = n64748 ^ n64749;
  assign n64726 = n64756 & n64757;
  assign n64746 = n64727 & n64707;
  assign n64744 = ~n64727;
  assign n64759 = n64762 & n64763;
  assign n64765 = n64771 & n64772;
  assign n64736 = ~n64786;
  assign n64775 = n377 ^ n64798;
  assign n64813 = n64827 & n64828;
  assign n63322 = n64715 ^ n64723;
  assign n64699 = ~n64724;
  assign n64706 = n64726 ^ n64727;
  assign n64714 = ~n64723;
  assign n64728 = n60730 & n64739;
  assign n64729 = n60730 & n63398;
  assign n64730 = ~n64726;
  assign n60748 = ~n60730;
  assign n64738 = n64744 & n64745;
  assign n64731 = ~n64746;
  assign n64742 = ~n64759;
  assign n64750 = ~n64765;
  assign n64665 = n64774 ^ n64775;
  assign n64752 = n64775 & n64774;
  assign n64799 = ~n64813;
  assign n64673 = n64706 ^ n64707;
  assign n64579 = ~n63322;
  assign n64681 = n64714 & n64715;
  assign n63515 = ~n64728;
  assign n64708 = ~n64729;
  assign n64718 = n64730 & n64731;
  assign n64719 = n60748 & n62108;
  assign n64721 = n60748 & n63494;
  assign n64705 = ~n64738;
  assign n64716 = n64742 & n64743;
  assign n64732 = n64750 & n64751;
  assign n64758 = n64665 & n62029;
  assign n64747 = ~n64665;
  assign n64776 = n64799 & n64800;
  assign n64685 = n64673 & n15399;
  assign n64687 = ~n64673;
  assign n64700 = n64716 ^ n64717;
  assign n64704 = ~n64718;
  assign n64709 = ~n64719;
  assign n63497 = ~n64721;
  assign n64711 = n64732 ^ n62100;
  assign n64713 = ~n64716;
  assign n64735 = ~n64732;
  assign n64740 = n64747 & n62078;
  assign n64669 = ~n64758;
  assign n64753 = n64776 ^ n64777;
  assign n64675 = ~n64685;
  assign n64679 = n64687 & n406;
  assign n64682 = n407 ^ n64700;
  assign n64688 = n64704 & n64705;
  assign n64662 = n64708 & n64709;
  assign n60649 = n64710 ^ n64711;
  assign n64703 = n64712 & n64713;
  assign n64720 = n64735 & n64736;
  assign n64693 = ~n64740;
  assign n64627 = n64752 ^ n64753;
  assign n64661 = ~n64679;
  assign n63288 = n64681 ^ n64682;
  assign n64635 = n64682 & n64681;
  assign n64663 = n64688 ^ n64689;
  assign n64690 = n60649 & n64696;
  assign n64695 = n64688 & n64697;
  assign n64694 = n60649 & n63384;
  assign n60698 = ~n60649;
  assign n64677 = ~n64662;
  assign n64691 = ~n64688;
  assign n64698 = ~n64703;
  assign n64701 = ~n64720;
  assign n64733 = n64627 & n61986;
  assign n64734 = ~n64627;
  assign n64640 = n64662 ^ n64663;
  assign n64516 = ~n63288;
  assign n63473 = ~n64690;
  assign n64683 = n64691 & n64689;
  assign n64684 = n60698 & n62100;
  assign n64678 = n60698 & n63457;
  assign n64671 = ~n64694;
  assign n64676 = ~n64695;
  assign n64672 = n64698 & n64699;
  assign n64686 = n64701 & n64702;
  assign n64632 = ~n64733;
  assign n64722 = n64734 & n62021;
  assign n64646 = n64640 & n405;
  assign n64655 = ~n64640;
  assign n64657 = n64672 ^ n64673;
  assign n64664 = n64676 & n64677;
  assign n63449 = ~n64678;
  assign n64659 = ~n64683;
  assign n64670 = ~n64684;
  assign n64674 = ~n64672;
  assign n64666 = n64686 ^ n62029;
  assign n64692 = ~n64686;
  assign n64651 = ~n64722;
  assign n64614 = ~n64646;
  assign n64641 = n64655 & n15354;
  assign n64636 = n406 ^ n64657;
  assign n64658 = ~n64664;
  assign n60570 = n64665 ^ n64666;
  assign n64618 = n64670 & n64671;
  assign n64667 = n64674 & n64675;
  assign n64680 = n64692 & n64693;
  assign n63239 = n64635 ^ n64636;
  assign n64630 = ~n64641;
  assign n64597 = n64636 & n64635;
  assign n64648 = n64618 & n64634;
  assign n64633 = n64658 & n64659;
  assign n64656 = n60570 & n63406;
  assign n64647 = n60570 & n63340;
  assign n64652 = ~n64618;
  assign n60641 = ~n60570;
  assign n64660 = ~n64667;
  assign n64668 = ~n64680;
  assign n64504 = ~n63239;
  assign n64619 = n64633 ^ n64634;
  assign n64625 = ~n64647;
  assign n64637 = ~n64648;
  assign n64643 = n60641 & n62029;
  assign n64645 = n64652 & n64653;
  assign n64642 = n60641 & n64654;
  assign n63429 = ~n64656;
  assign n64638 = ~n64633;
  assign n64639 = n64660 & n64661;
  assign n64649 = n64668 & n64669;
  assign n64593 = n64618 ^ n64619;
  assign n64626 = n64637 & n64638;
  assign n64617 = n64639 ^ n64640;
  assign n63409 = ~n64642;
  assign n64624 = ~n64643;
  assign n64622 = ~n64645;
  assign n64629 = ~n64639;
  assign n64628 = n64649 ^ n61986;
  assign n64650 = ~n64649;
  assign n64599 = n64593 & n15327;
  assign n64594 = ~n64593;
  assign n64598 = n405 ^ n64617;
  assign n64576 = n64624 & n64625;
  assign n64621 = ~n64626;
  assign n60488 = n64627 ^ n64628;
  assign n64623 = n64629 & n64630;
  assign n64644 = n64650 & n64651;
  assign n64584 = n64594 & n404;
  assign n63215 = n64597 ^ n64598;
  assign n64582 = ~n64599;
  assign n64602 = ~n64598;
  assign n64607 = n60488 & n63282;
  assign n64612 = n64576 & n64620;
  assign n64611 = n60488 & n63374;
  assign n64595 = n64621 & n64622;
  assign n64608 = ~n64576;
  assign n64613 = ~n64623;
  assign n60546 = ~n60488;
  assign n64631 = ~n64644;
  assign n64442 = ~n63215;
  assign n64564 = ~n64584;
  assign n64577 = n64595 ^ n64596;
  assign n64549 = n64602 & n64597;
  assign n64600 = ~n64595;
  assign n64589 = ~n64607;
  assign n64603 = n64608 & n64596;
  assign n63388 = ~n64611;
  assign n64601 = ~n64612;
  assign n64606 = n60546 & n61986;
  assign n64592 = n64613 & n64614;
  assign n64604 = n60546 & n64616;
  assign n64615 = n64631 & n64632;
  assign n64545 = n64576 ^ n64577;
  assign n64573 = n64592 ^ n64593;
  assign n64585 = n64600 & n64601;
  assign n64583 = ~n64592;
  assign n64575 = ~n64603;
  assign n63363 = ~n64604;
  assign n64588 = ~n64606;
  assign n64587 = n64615 ^ n61906;
  assign n64609 = ~n64615;
  assign n64560 = n64545 & n403;
  assign n64557 = ~n64545;
  assign n64550 = n404 ^ n64573;
  assign n64580 = n64582 & n64583;
  assign n64574 = ~n64585;
  assign n60401 = n64586 ^ n64587;
  assign n64542 = n64588 & n64589;
  assign n64605 = n64609 & n64610;
  assign n63148 = n64549 ^ n64550;
  assign n64551 = n64557 & n15296;
  assign n64506 = n64550 & n64549;
  assign n64519 = ~n64560;
  assign n64558 = n64574 & n64575;
  assign n64568 = n64542 & n64578;
  assign n64567 = n60401 & n64579;
  assign n64569 = n60401 & n61939;
  assign n64563 = ~n64580;
  assign n64572 = ~n64542;
  assign n60491 = ~n60401;
  assign n64590 = ~n64605;
  assign n64399 = ~n63148;
  assign n64535 = ~n64551;
  assign n64512 = ~n64506;
  assign n64543 = n64558 ^ n64559;
  assign n64544 = n64563 & n64564;
  assign n64554 = ~n64558;
  assign n63325 = ~n64567;
  assign n64555 = ~n64568;
  assign n64552 = ~n64569;
  assign n64565 = n60491 & n63322;
  assign n64566 = n64572 & n64559;
  assign n64561 = n60491 & n63268;
  assign n64581 = n64590 & n64591;
  assign n64493 = n64542 ^ n64543;
  assign n64528 = n64544 ^ n64545;
  assign n64546 = n64554 & n64555;
  assign n64536 = ~n64544;
  assign n64553 = ~n64561;
  assign n63347 = ~n64565;
  assign n64538 = ~n64566;
  assign n64571 = n64581 & n61831;
  assign n64570 = ~n64581;
  assign n64515 = n64493 & n402;
  assign n64507 = n403 ^ n64528;
  assign n64517 = ~n64493;
  assign n64532 = n64535 & n64536;
  assign n64537 = ~n64546;
  assign n64499 = n64552 & n64553;
  assign n64562 = n64570 & n61873;
  assign n64548 = ~n64571;
  assign n63098 = n64506 ^ n64507;
  assign n64463 = n64507 & n64512;
  assign n64480 = ~n64515;
  assign n64513 = n64517 & n15251;
  assign n64518 = ~n64532;
  assign n64526 = n64537 & n64538;
  assign n64530 = n64499 & n64539;
  assign n64531 = ~n64499;
  assign n64547 = n64548 & n64556;
  assign n64541 = ~n64562;
  assign n64371 = ~n63098;
  assign n64451 = ~n64463;
  assign n64501 = ~n64513;
  assign n64492 = n64518 & n64519;
  assign n64500 = n64526 ^ n64527;
  assign n64523 = ~n64530;
  assign n64529 = n64531 & n64527;
  assign n64522 = ~n64526;
  assign n64540 = ~n64547;
  assign n64533 = n64541 & n64548;
  assign n64483 = n64492 ^ n64493;
  assign n64453 = n64499 ^ n64500;
  assign n64502 = ~n64492;
  assign n64509 = n64522 & n64523;
  assign n64495 = ~n64529;
  assign n60316 = n64533 ^ n64534;
  assign n64521 = n64540 & n64541;
  assign n64464 = n402 ^ n64483;
  assign n64481 = n64453 & n401;
  assign n64482 = ~n64453;
  assign n64489 = n64501 & n64502;
  assign n64494 = ~n64509;
  assign n64510 = n60316 & n64516;
  assign n60196 = n64520 ^ n64521;
  assign n64511 = n60316 & n63194;
  assign n60384 = ~n60316;
  assign n64524 = ~n64521;
  assign n63037 = n64463 ^ n64464;
  assign n64450 = ~n64464;
  assign n64441 = ~n64481;
  assign n64474 = n64482 & n15210;
  assign n64479 = ~n64489;
  assign n64475 = n64494 & n64495;
  assign n64496 = n60196 & n64504;
  assign n64503 = n60196 & n63166;
  assign n63308 = ~n64510;
  assign n64508 = n60384 & n61873;
  assign n64505 = n60384 & n63288;
  assign n64490 = ~n64511;
  assign n60343 = ~n60196;
  assign n64514 = n64524 & n64525;
  assign n64321 = ~n63037;
  assign n64414 = n64450 & n64451;
  assign n64459 = ~n64474;
  assign n64468 = n64475 ^ n64471;
  assign n64452 = n64479 & n64480;
  assign n64466 = ~n64475;
  assign n63262 = ~n64496;
  assign n64487 = n60343 & n61762;
  assign n64488 = n60343 & n63239;
  assign n64478 = ~n64503;
  assign n63284 = ~n64505;
  assign n64491 = ~n64508;
  assign n64497 = ~n64514;
  assign n64446 = n64452 ^ n64453;
  assign n64458 = ~n64452;
  assign n64477 = ~n64487;
  assign n63242 = ~n64488;
  assign n64467 = n64490 & n64491;
  assign n64484 = n64497 & n64498;
  assign n64425 = n401 ^ n64446;
  assign n64449 = n64458 & n64459;
  assign n64416 = n64467 ^ n64468;
  assign n64472 = n64467 & n64476;
  assign n64422 = n64477 & n64478;
  assign n64462 = n64484 ^ n61660;
  assign n64470 = ~n64467;
  assign n64485 = ~n64484;
  assign n62979 = n64414 ^ n64425;
  assign n64413 = ~n64425;
  assign n64434 = n64416 & n400;
  assign n64439 = ~n64416;
  assign n64440 = ~n64449;
  assign n60098 = n64461 ^ n64462;
  assign n64460 = n64422 & n64408;
  assign n64469 = n64470 & n64471;
  assign n64465 = ~n64472;
  assign n64456 = ~n64422;
  assign n64473 = n64485 & n64486;
  assign n64288 = ~n62979;
  assign n64380 = n64413 & n64414;
  assign n64397 = ~n64434;
  assign n64430 = n64439 & n15157;
  assign n64415 = n64440 & n64441;
  assign n64445 = n60098 & n63091;
  assign n64435 = n60098 & n63215;
  assign n60178 = ~n60098;
  assign n64448 = n64456 & n64457;
  assign n64420 = ~n64460;
  assign n64447 = n64465 & n64466;
  assign n64444 = ~n64469;
  assign n64454 = ~n64473;
  assign n64390 = ~n64380;
  assign n64395 = n64415 ^ n64416;
  assign n64428 = ~n64415;
  assign n64429 = ~n64430;
  assign n63217 = ~n64435;
  assign n64431 = n60178 & n64442;
  assign n64432 = n60178 & n61660;
  assign n64423 = ~n64445;
  assign n64443 = ~n64447;
  assign n64405 = ~n64448;
  assign n64436 = n64454 & n64455;
  assign n64381 = n400 ^ n64395;
  assign n64411 = n64428 & n64429;
  assign n63200 = ~n64431;
  assign n64424 = ~n64432;
  assign n64418 = n64436 ^ n61575;
  assign n64421 = n64443 & n64444;
  assign n64437 = ~n64436;
  assign n62900 = n64380 ^ n64381;
  assign n64334 = n64381 & n64390;
  assign n64396 = ~n64411;
  assign n60021 = n64417 ^ n64418;
  assign n64407 = n64421 ^ n64422;
  assign n64385 = n64423 & n64424;
  assign n64419 = ~n64421;
  assign n64433 = n64437 & n64438;
  assign n64246 = ~n62900;
  assign n64386 = n64396 & n64397;
  assign n64387 = n64407 ^ n64408;
  assign n64409 = n60021 & n63148;
  assign n64401 = n60021 & n61575;
  assign n64400 = n64385 & n64410;
  assign n64398 = ~n64385;
  assign n60135 = ~n60021;
  assign n64412 = n64419 & n64420;
  assign n64426 = ~n64433;
  assign n64363 = n64386 ^ n64387;
  assign n64374 = n64387 & n15109;
  assign n64369 = ~n64386;
  assign n64377 = ~n64387;
  assign n64391 = n64398 & n64361;
  assign n64392 = n60135 & n64399;
  assign n64382 = ~n64400;
  assign n64375 = ~n64401;
  assign n64393 = n60135 & n63065;
  assign n63151 = ~n64409;
  assign n64404 = ~n64412;
  assign n64406 = n64426 & n64427;
  assign n64335 = n415 ^ n64363;
  assign n64368 = ~n64374;
  assign n64372 = n64377 & n415;
  assign n64356 = ~n64391;
  assign n63170 = ~n64392;
  assign n64376 = ~n64393;
  assign n64384 = n64404 & n64405;
  assign n64379 = n64406 ^ n61491;
  assign n64402 = ~n64406;
  assign n64206 = n64334 ^ n64335;
  assign n64336 = ~n64335;
  assign n64362 = n64368 & n64369;
  assign n64350 = ~n64372;
  assign n64326 = n64375 & n64376;
  assign n59969 = n64378 ^ n64379;
  assign n64360 = n64384 ^ n64385;
  assign n64383 = ~n64384;
  assign n64394 = n64402 & n64403;
  assign n64291 = n64336 & n64334;
  assign n64331 = n64360 ^ n64361;
  assign n64349 = ~n64362;
  assign n64359 = n59969 & n62972;
  assign n64365 = n64326 & n64370;
  assign n64366 = n59969 & n64371;
  assign n64364 = ~n64326;
  assign n60043 = ~n59969;
  assign n64373 = n64382 & n64383;
  assign n64388 = ~n64394;
  assign n64330 = n64349 & n64350;
  assign n64338 = n64331 & n414;
  assign n64337 = ~n64331;
  assign n64351 = n60043 & n61491;
  assign n64354 = n60043 & n63098;
  assign n64344 = ~n64359;
  assign n64353 = n64364 & n64340;
  assign n64341 = ~n64365;
  assign n63126 = ~n64366;
  assign n64355 = ~n64373;
  assign n64367 = n64388 & n64389;
  assign n64309 = n64330 ^ n64331;
  assign n64332 = n64337 & n15067;
  assign n64304 = ~n64338;
  assign n64328 = ~n64330;
  assign n64343 = ~n64351;
  assign n64324 = ~n64353;
  assign n63095 = ~n64354;
  assign n64339 = n64355 & n64356;
  assign n64346 = n64367 ^ n61410;
  assign n64357 = ~n64367;
  assign n64292 = n414 ^ n64309;
  assign n64329 = ~n64332;
  assign n64327 = n64339 ^ n64340;
  assign n64282 = n64343 & n64344;
  assign n59885 = n64345 ^ n64346;
  assign n64342 = ~n64339;
  assign n64352 = n64357 & n64358;
  assign n64268 = n64291 ^ n64292;
  assign n64244 = n64292 & n64291;
  assign n64277 = n64326 ^ n64327;
  assign n64314 = n64328 & n64329;
  assign n64316 = n59885 & n63037;
  assign n64322 = n59885 & n61470;
  assign n64315 = n64282 & n64296;
  assign n64319 = ~n64282;
  assign n59958 = ~n59885;
  assign n64333 = n64341 & n64342;
  assign n64347 = ~n64352;
  assign n61006 = n64268 ^ n62048;
  assign n64267 = n64268 & n62048;
  assign n64266 = ~n64268;
  assign n64235 = ~n64244;
  assign n64305 = n64277 & n413;
  assign n64303 = ~n64314;
  assign n64306 = ~n64277;
  assign n64312 = n59958 & n62897;
  assign n64299 = ~n64315;
  assign n63032 = ~n64316;
  assign n64310 = n64319 & n64320;
  assign n64311 = n59958 & n64321;
  assign n64301 = ~n64322;
  assign n64323 = ~n64333;
  assign n64325 = n64347 & n64348;
  assign n64248 = n61006 & n63113;
  assign n61004 = ~n61006;
  assign n64159 = n64266 & n62048;
  assign n64225 = ~n64267;
  assign n64276 = n64303 & n64304;
  assign n64262 = ~n64305;
  assign n64294 = n64306 & n15056;
  assign n64285 = ~n64310;
  assign n63071 = ~n64311;
  assign n64302 = ~n64312;
  assign n64295 = n64323 & n64324;
  assign n64308 = n64325 ^ n61336;
  assign n64317 = ~n64325;
  assign n64224 = ~n64248;
  assign n64251 = n64276 ^ n64277;
  assign n64275 = ~n64276;
  assign n64274 = ~n64294;
  assign n64283 = n64295 ^ n64296;
  assign n64239 = n64301 & n64302;
  assign n59806 = n64307 ^ n64308;
  assign n64300 = ~n64295;
  assign n64313 = n64317 & n64318;
  assign n64197 = n64224 & n64225;
  assign n64245 = n413 ^ n64251;
  assign n64272 = n64274 & n64275;
  assign n64233 = n64282 ^ n64283;
  assign n64289 = n64239 & n64253;
  assign n64290 = n59806 & n62979;
  assign n64278 = n59806 & n62820;
  assign n59866 = ~n59806;
  assign n64286 = ~n64239;
  assign n64293 = n64299 & n64300;
  assign n64297 = ~n64313;
  assign n64179 = n64197 ^ n64198;
  assign n64199 = ~n64197;
  assign n64221 = n64244 ^ n64245;
  assign n64234 = ~n64245;
  assign n64258 = n64233 & n14988;
  assign n64263 = ~n64233;
  assign n64261 = ~n64272;
  assign n64254 = ~n64278;
  assign n64269 = n64286 & n64287;
  assign n64273 = n59866 & n64288;
  assign n64270 = n59866 & n61415;
  assign n64264 = ~n64289;
  assign n63006 = ~n64290;
  assign n64284 = ~n64293;
  assign n64279 = n64297 & n64298;
  assign n62434 = n423 ^ n64179;
  assign n64003 = n64179 & n423;
  assign n64064 = n64199 & n64200;
  assign n64205 = n64221 & n61956;
  assign n64214 = ~n64221;
  assign n64195 = n64234 & n64235;
  assign n64237 = ~n64258;
  assign n64232 = n64261 & n64262;
  assign n64249 = n64263 & n412;
  assign n64229 = ~n64269;
  assign n64255 = ~n64270;
  assign n62976 = ~n64273;
  assign n64260 = n64279 ^ n61264;
  assign n64252 = n64284 & n64285;
  assign n64280 = ~n64279;
  assign n62467 = ~n62434;
  assign n64176 = ~n64205;
  assign n64201 = n64214 & n61962;
  assign n64194 = ~n64195;
  assign n64207 = n64232 ^ n64233;
  assign n64210 = ~n64249;
  assign n64238 = ~n64232;
  assign n64240 = n64252 ^ n64253;
  assign n64182 = n64254 & n64255;
  assign n59733 = n64259 ^ n64260;
  assign n64265 = ~n64252;
  assign n64271 = n64280 & n64281;
  assign n64190 = ~n64201;
  assign n64196 = n412 ^ n64207;
  assign n64222 = n64237 & n64238;
  assign n64187 = n64239 ^ n64240;
  assign n64231 = n59733 & n64246;
  assign n64243 = n64182 & n64247;
  assign n64236 = n59733 & n62751;
  assign n59783 = ~n59733;
  assign n64230 = ~n64182;
  assign n64250 = n64264 & n64265;
  assign n64256 = ~n64271;
  assign n64178 = n64190 & n64159;
  assign n64180 = n64190 & n64176;
  assign n64122 = n64195 ^ n64196;
  assign n64193 = ~n64196;
  assign n64213 = n64187 & n14942;
  assign n64218 = ~n64187;
  assign n64209 = ~n64222;
  assign n64223 = n64230 & n64212;
  assign n62946 = ~n64231;
  assign n64226 = n59783 & n61322;
  assign n64220 = ~n64236;
  assign n64227 = n59783 & n62900;
  assign n64216 = ~n64243;
  assign n64228 = ~n64250;
  assign n64241 = n64256 & n64257;
  assign n64169 = n64122 & n61852;
  assign n64175 = ~n64178;
  assign n64160 = ~n64180;
  assign n64162 = ~n64122;
  assign n64143 = n64193 & n64194;
  assign n64186 = n64209 & n64210;
  assign n64188 = ~n64213;
  assign n64203 = n64218 & n411;
  assign n64192 = ~n64223;
  assign n64219 = ~n64226;
  assign n62903 = ~n64227;
  assign n64211 = n64228 & n64229;
  assign n59709 = n64241 ^ n64242;
  assign n60904 = n64159 ^ n64160;
  assign n64161 = n64162 & n61889;
  assign n64148 = ~n64169;
  assign n64156 = n64175 & n64176;
  assign n64155 = ~n64143;
  assign n64163 = n64186 ^ n64187;
  assign n64189 = ~n64186;
  assign n64174 = ~n64203;
  assign n62868 = n64206 ^ n59709;
  assign n64183 = n64211 ^ n64212;
  assign n64151 = n64219 & n64220;
  assign n64215 = n59709 & n62754;
  assign n64217 = ~n64211;
  assign n64208 = ~n59709;
  assign n64140 = n60904 & n63020;
  assign n60899 = ~n60904;
  assign n64142 = ~n64156;
  assign n64135 = ~n64161;
  assign n64144 = n411 ^ n64163;
  assign n64147 = n64182 ^ n64183;
  assign n64181 = n64188 & n64189;
  assign n64154 = ~n64151;
  assign n64204 = n64208 & n62824;
  assign n64184 = ~n64215;
  assign n64202 = n64216 & n64217;
  assign n64125 = ~n64140;
  assign n64121 = n64142 ^ n61889;
  assign n64138 = n60899 & n61956;
  assign n64093 = n64143 ^ n64144;
  assign n64139 = n64148 & n64142;
  assign n64110 = n64144 & n64155;
  assign n64164 = n64147 & n410;
  assign n64173 = ~n64181;
  assign n64172 = ~n64147;
  assign n64191 = ~n64202;
  assign n64185 = ~n64204;
  assign n60817 = n64121 ^ n64122;
  assign n64131 = n64093 & n61779;
  assign n64124 = ~n64138;
  assign n64134 = ~n64139;
  assign n64127 = ~n64093;
  assign n64119 = ~n64110;
  assign n64133 = ~n64164;
  assign n64157 = n64172 & n14910;
  assign n64146 = n64173 & n64174;
  assign n64170 = n64184 & n64185;
  assign n64165 = n64191 & n64192;
  assign n64102 = n60817 & n62915;
  assign n60847 = ~n60817;
  assign n64108 = n64124 & n64125;
  assign n64126 = n64127 & n61811;
  assign n64118 = ~n64131;
  assign n64116 = n64134 & n64135;
  assign n64130 = n64146 ^ n64147;
  assign n64149 = ~n64157;
  assign n64150 = ~n64146;
  assign n64152 = n64165 ^ n64166;
  assign n64099 = n64170 ^ n64171;
  assign n64177 = n64165 & n64166;
  assign n64167 = ~n64165;
  assign n64085 = ~n64102;
  assign n64101 = n60847 & n61889;
  assign n64107 = n64108 & n64109;
  assign n64094 = n64116 ^ n61779;
  assign n64105 = ~n64108;
  assign n64117 = ~n64116;
  assign n64096 = ~n64126;
  assign n64111 = n410 ^ n64130;
  assign n64141 = n64149 & n64150;
  assign n64115 = n64151 ^ n64152;
  assign n64158 = n64167 & n64168;
  assign n64153 = ~n64177;
  assign n60750 = n64093 ^ n64094;
  assign n64084 = ~n64101;
  assign n64100 = n64105 & n64106;
  assign n64088 = ~n64107;
  assign n64055 = n64110 ^ n64111;
  assign n64103 = n64117 & n64118;
  assign n64075 = n64111 & n64119;
  assign n64128 = n64115 & n14879;
  assign n64132 = ~n64141;
  assign n64129 = ~n64115;
  assign n64145 = n64153 & n64154;
  assign n64137 = ~n64158;
  assign n64079 = n60750 & n62853;
  assign n64042 = n64084 & n64085;
  assign n60782 = ~n60750;
  assign n64086 = n64088 & n64064;
  assign n64089 = n64055 & n61713;
  assign n64074 = ~n64100;
  assign n64095 = ~n64103;
  assign n64092 = ~n64055;
  assign n64113 = ~n64128;
  assign n64123 = n64129 & n409;
  assign n64114 = n64132 & n64133;
  assign n64136 = ~n64145;
  assign n64059 = ~n64079;
  assign n64068 = n64042 & n64082;
  assign n64067 = n60782 & n61811;
  assign n64070 = ~n64042;
  assign n64073 = ~n64086;
  assign n64083 = n64074 & n64088;
  assign n64061 = ~n64089;
  assign n64087 = n64092 & n61695;
  assign n64078 = n64095 & n64096;
  assign n64097 = n64114 ^ n64115;
  assign n64112 = ~n64114;
  assign n64091 = ~n64123;
  assign n64120 = n64136 & n64137;
  assign n64058 = ~n64067;
  assign n64062 = ~n64068;
  assign n64066 = n64070 & n64051;
  assign n64050 = n64073 & n64074;
  assign n64056 = n64078 ^ n61695;
  assign n64065 = ~n64083;
  assign n64072 = ~n64087;
  assign n64071 = ~n64078;
  assign n64076 = n409 ^ n64097;
  assign n64104 = n64112 & n64113;
  assign n64098 = n408 ^ n64120;
  assign n64043 = n64050 ^ n64051;
  assign n60656 = n64055 ^ n64056;
  assign n63999 = n64058 & n64059;
  assign n64047 = n64064 ^ n64065;
  assign n64034 = ~n64066;
  assign n64063 = ~n64050;
  assign n64069 = n64071 & n64072;
  assign n64015 = n64075 ^ n64076;
  assign n64077 = ~n64076;
  assign n64081 = n64098 ^ n64099;
  assign n64090 = ~n64104;
  assign n63990 = n64042 ^ n64043;
  assign n64039 = n63999 & n64018;
  assign n64036 = n60656 & n61713;
  assign n64046 = n64047 & n7609;
  assign n60667 = ~n60656;
  assign n64040 = ~n63999;
  assign n64045 = ~n64047;
  assign n64048 = n64062 & n64063;
  assign n64052 = n64015 & n61633;
  assign n64060 = ~n64069;
  assign n64057 = ~n64015;
  assign n64053 = n64077 & n64075;
  assign n64080 = n64090 & n64091;
  assign n64013 = n63990 & n421;
  assign n64021 = ~n63990;
  assign n64019 = ~n64036;
  assign n64026 = n60667 & n62769;
  assign n64011 = ~n64039;
  assign n64029 = n64040 & n64041;
  assign n64035 = n64045 & n422;
  assign n64025 = ~n64046;
  assign n64033 = ~n64048;
  assign n64023 = ~n64052;
  assign n64049 = n64057 & n61611;
  assign n64032 = n64060 & n64061;
  assign n64054 = n64080 ^ n64081;
  assign n63972 = ~n64013;
  assign n64007 = n64021 & n7523;
  assign n64020 = ~n64026;
  assign n63995 = ~n64029;
  assign n64024 = n64025 & n64003;
  assign n64016 = n64032 ^ n61611;
  assign n64017 = n64033 & n64034;
  assign n64010 = ~n64035;
  assign n64037 = ~n64032;
  assign n64038 = ~n64049;
  assign n64044 = n64053 ^ n64054;
  assign n63985 = ~n64007;
  assign n60556 = n64015 ^ n64016;
  assign n64000 = n64017 ^ n64018;
  assign n63964 = n64019 & n64020;
  assign n64009 = ~n64024;
  assign n64014 = n64025 & n64010;
  assign n64012 = ~n64017;
  assign n64027 = n64037 & n64038;
  assign n64031 = n64044 & n61546;
  assign n64030 = ~n64044;
  assign n63946 = n63999 ^ n64000;
  assign n63997 = n63964 & n64005;
  assign n63998 = n60556 & n61633;
  assign n63996 = ~n63964;
  assign n60590 = ~n60556;
  assign n63989 = n64009 & n64010;
  assign n64006 = n64011 & n64012;
  assign n64004 = ~n64014;
  assign n64022 = ~n64027;
  assign n64028 = n64030 & n61528;
  assign n63977 = ~n64031;
  assign n63983 = n63946 & n7437;
  assign n63973 = ~n63946;
  assign n63968 = n63989 ^ n63990;
  assign n63988 = n63996 & n63982;
  assign n63979 = ~n63997;
  assign n63993 = n60590 & n62698;
  assign n63974 = ~n63998;
  assign n63980 = n64003 ^ n64004;
  assign n63986 = ~n63989;
  assign n63994 = ~n64006;
  assign n63991 = n64022 & n64023;
  assign n64002 = ~n64028;
  assign n63955 = n421 ^ n63968;
  assign n63970 = n63973 & n420;
  assign n63676 = n63980 ^ n62467;
  assign n63947 = ~n63983;
  assign n63954 = n63980 & n62467;
  assign n63984 = n63985 & n63986;
  assign n63957 = ~n63988;
  assign n63975 = ~n63993;
  assign n63981 = n63994 & n63995;
  assign n64001 = ~n63991;
  assign n64008 = n64002 & n63977;
  assign n62375 = n63954 ^ n63955;
  assign n63949 = ~n63955;
  assign n63927 = ~n63970;
  assign n62410 = ~n63676;
  assign n63950 = ~n63954;
  assign n63919 = n63974 & n63975;
  assign n63965 = n63981 ^ n63982;
  assign n63971 = ~n63984;
  assign n63978 = ~n63981;
  assign n63987 = n64001 & n64002;
  assign n63992 = ~n64008;
  assign n63649 = ~n62375;
  assign n63912 = n63949 & n63950;
  assign n63911 = n63964 ^ n63965;
  assign n63963 = n63919 & n63934;
  assign n63945 = n63971 & n63972;
  assign n63958 = ~n63919;
  assign n63969 = n63978 & n63979;
  assign n63976 = ~n63987;
  assign n60452 = n63991 ^ n63992;
  assign n63932 = n63911 & n419;
  assign n63930 = n63945 ^ n63946;
  assign n63936 = ~n63911;
  assign n63953 = n63958 & n63959;
  assign n63940 = ~n63963;
  assign n63948 = ~n63945;
  assign n63956 = ~n63969;
  assign n63967 = n60452 & n61546;
  assign n63960 = n63976 & n63977;
  assign n60516 = ~n60452;
  assign n63913 = n420 ^ n63930;
  assign n63894 = ~n63932;
  assign n63931 = n63936 & n7333;
  assign n63943 = n63947 & n63948;
  assign n63922 = ~n63953;
  assign n63933 = n63956 & n63957;
  assign n63942 = n63960 ^ n61451;
  assign n63952 = ~n63967;
  assign n63966 = n60516 & n62644;
  assign n63961 = ~n63960;
  assign n62353 = n63912 ^ n63913;
  assign n63878 = n63913 & n63912;
  assign n63914 = ~n63931;
  assign n63920 = n63933 ^ n63934;
  assign n60370 = n63941 ^ n63942;
  assign n63926 = ~n63943;
  assign n63939 = ~n63933;
  assign n63944 = n63961 & n63962;
  assign n63951 = ~n63966;
  assign n63608 = ~n62353;
  assign n63882 = ~n63878;
  assign n63877 = n63919 ^ n63920;
  assign n63916 = n60370 & n61451;
  assign n63910 = n63926 & n63927;
  assign n60432 = ~n60370;
  assign n63928 = n63939 & n63940;
  assign n63937 = ~n63944;
  assign n63880 = n63951 & n63952;
  assign n63902 = n63877 & n7273;
  assign n63897 = ~n63877;
  assign n63892 = n63910 ^ n63911;
  assign n63904 = ~n63916;
  assign n63908 = n60432 & n62603;
  assign n63915 = ~n63910;
  assign n63921 = ~n63928;
  assign n63929 = n63880 & n63935;
  assign n63923 = n63937 & n63938;
  assign n63925 = ~n63880;
  assign n63879 = n419 ^ n63892;
  assign n63895 = n63897 & n418;
  assign n63874 = ~n63902;
  assign n63903 = ~n63908;
  assign n63907 = n63914 & n63915;
  assign n63898 = n63921 & n63922;
  assign n63918 = n63923 & n61371;
  assign n63924 = n63925 & n63899;
  assign n63906 = ~n63929;
  assign n63917 = ~n63923;
  assign n62305 = n63878 ^ n63879;
  assign n63842 = n63879 & n63882;
  assign n63857 = ~n63895;
  assign n63881 = n63898 ^ n63899;
  assign n63847 = n63903 & n63904;
  assign n63893 = ~n63907;
  assign n63905 = ~n63898;
  assign n63909 = n63917 & n61405;
  assign n63901 = ~n63918;
  assign n63885 = ~n63924;
  assign n63561 = ~n62305;
  assign n63844 = ~n63842;
  assign n63841 = n63880 ^ n63881;
  assign n63886 = n63847 & n63891;
  assign n63876 = n63893 & n63894;
  assign n63883 = ~n63847;
  assign n63896 = n63905 & n63906;
  assign n63900 = n63901 & n63887;
  assign n63890 = ~n63909;
  assign n63862 = n63841 & n417;
  assign n63861 = ~n63841;
  assign n63855 = n63876 ^ n63877;
  assign n63873 = n63883 & n63868;
  assign n63863 = ~n63886;
  assign n63875 = ~n63876;
  assign n63884 = ~n63896;
  assign n63889 = ~n63900;
  assign n63888 = n63890 & n63901;
  assign n63843 = n418 ^ n63855;
  assign n63858 = n63861 & n7227;
  assign n63823 = ~n63862;
  assign n63846 = ~n63873;
  assign n63872 = n63874 & n63875;
  assign n63867 = n63884 & n63885;
  assign n60290 = n63887 ^ n63888;
  assign n63869 = n63889 & n63890;
  assign n62282 = n63842 ^ n63843;
  assign n63801 = n63843 & n63844;
  assign n63839 = ~n63858;
  assign n63848 = n63867 ^ n63868;
  assign n63853 = n63869 ^ n61289;
  assign n63856 = ~n63872;
  assign n63865 = n60290 & n61405;
  assign n60325 = ~n60290;
  assign n63864 = ~n63867;
  assign n63870 = ~n63869;
  assign n63524 = ~n62282;
  assign n63804 = n63847 ^ n63848;
  assign n60184 = n63853 ^ n63854;
  assign n63840 = n63856 & n63857;
  assign n63859 = n63863 & n63864;
  assign n63860 = n60325 & n62568;
  assign n63849 = ~n63865;
  assign n63866 = n63870 & n63871;
  assign n63832 = n63804 & n416;
  assign n63837 = n60184 & n61289;
  assign n63819 = n63840 ^ n63841;
  assign n63829 = ~n63804;
  assign n60243 = ~n60184;
  assign n63838 = ~n63840;
  assign n63845 = ~n63859;
  assign n63850 = ~n63860;
  assign n63851 = ~n63866;
  assign n63802 = n417 ^ n63819;
  assign n63820 = n63829 & n7122;
  assign n63781 = ~n63832;
  assign n63824 = n60243 & n62495;
  assign n63811 = ~n63837;
  assign n63834 = n63838 & n63839;
  assign n63827 = n63845 & n63846;
  assign n63808 = n63849 & n63850;
  assign n63833 = n63851 & n63852;
  assign n62222 = n63801 ^ n63802;
  assign n63807 = ~n63802;
  assign n63806 = ~n63820;
  assign n63812 = ~n63824;
  assign n63809 = n63827 ^ n63828;
  assign n63816 = n63833 ^ n61233;
  assign n63822 = ~n63834;
  assign n63825 = n63808 & n63828;
  assign n63814 = ~n63827;
  assign n63830 = ~n63808;
  assign n63835 = ~n63833;
  assign n63483 = ~n62222;
  assign n63763 = n63807 & n63801;
  assign n63798 = n63808 ^ n63809;
  assign n63751 = n63811 & n63812;
  assign n60093 = n63815 ^ n63816;
  assign n63803 = n63822 & n63823;
  assign n63813 = ~n63825;
  assign n63821 = n63830 & n63831;
  assign n63826 = n63835 & n63836;
  assign n63786 = n63798 & n7117;
  assign n63769 = ~n63763;
  assign n63791 = n60093 & n61233;
  assign n63783 = n63803 ^ n63804;
  assign n63785 = ~n63798;
  assign n63790 = n63751 & n63772;
  assign n60142 = ~n60093;
  assign n63794 = ~n63751;
  assign n63805 = ~n63803;
  assign n63810 = n63813 & n63814;
  assign n63793 = ~n63821;
  assign n63817 = ~n63826;
  assign n63764 = n416 ^ n63783;
  assign n63782 = n63785 & n431;
  assign n63767 = ~n63786;
  assign n63784 = n60142 & n62481;
  assign n63776 = ~n63790;
  assign n63779 = ~n63791;
  assign n63788 = n63794 & n63795;
  assign n63789 = n63805 & n63806;
  assign n63792 = ~n63810;
  assign n63799 = n63817 & n63818;
  assign n62182 = n63763 ^ n63764;
  assign n63721 = n63764 & n63769;
  assign n63744 = ~n63782;
  assign n63778 = ~n63784;
  assign n63754 = ~n63788;
  assign n63780 = ~n63789;
  assign n63771 = n63792 & n63793;
  assign n63770 = n63799 ^ n63800;
  assign n63796 = ~n63799;
  assign n63440 = ~n62182;
  assign n63765 = n63767 & n63744;
  assign n60032 = n61156 ^ n63770;
  assign n63752 = n63771 ^ n63772;
  assign n63711 = n63778 & n63779;
  assign n63747 = n63780 & n63781;
  assign n63773 = n63770 & n61156;
  assign n63777 = ~n63771;
  assign n63787 = n63796 & n63797;
  assign n63724 = n63751 ^ n63752;
  assign n63757 = n60032 & n62443;
  assign n63758 = n63711 & n63734;
  assign n63748 = ~n63765;
  assign n63755 = ~n63711;
  assign n60051 = ~n60032;
  assign n63746 = ~n63773;
  assign n63766 = ~n63747;
  assign n63768 = n63776 & n63777;
  assign n63774 = ~n63787;
  assign n63722 = n63747 ^ n63748;
  assign n63742 = n63724 & n7047;
  assign n63741 = ~n63724;
  assign n63750 = n63755 & n63756;
  assign n63745 = ~n63757;
  assign n63739 = ~n63758;
  assign n63759 = n63766 & n63767;
  assign n63753 = ~n63768;
  assign n63762 = n63774 & n63775;
  assign n62138 = n63721 ^ n63722;
  assign n63732 = n63741 & n430;
  assign n63725 = ~n63742;
  assign n63730 = ~n63722;
  assign n63696 = n63745 & n63746;
  assign n63720 = ~n63750;
  assign n63733 = n63753 & n63754;
  assign n63743 = ~n63759;
  assign n63736 = n63762 ^ n61084;
  assign n63760 = ~n63762;
  assign n63400 = ~n62138;
  assign n63688 = n63730 & n63721;
  assign n63708 = ~n63732;
  assign n63729 = n63696 & n63672;
  assign n63712 = n63733 ^ n63734;
  assign n63727 = ~n63696;
  assign n59922 = n63735 ^ n63736;
  assign n63723 = n63743 & n63744;
  assign n63740 = ~n63733;
  assign n63749 = n63760 & n63761;
  assign n63693 = ~n63688;
  assign n63685 = n63711 ^ n63712;
  assign n63706 = n63723 ^ n63724;
  assign n63713 = n63727 & n63728;
  assign n63701 = ~n63729;
  assign n63714 = n59922 & n61084;
  assign n59961 = ~n59922;
  assign n63726 = ~n63723;
  assign n63731 = n63739 & n63740;
  assign n63737 = ~n63749;
  assign n63689 = n430 ^ n63706;
  assign n63705 = n63685 & n7015;
  assign n63694 = ~n63685;
  assign n63682 = ~n63713;
  assign n63700 = ~n63714;
  assign n63710 = n59961 & n62383;
  assign n63716 = n63725 & n63726;
  assign n63719 = ~n63731;
  assign n63715 = n63737 & n63738;
  assign n62089 = n63688 ^ n63689;
  assign n63643 = n63689 & n63693;
  assign n63691 = n63694 & n429;
  assign n63686 = ~n63705;
  assign n63699 = ~n63710;
  assign n63698 = n63715 ^ n61048;
  assign n63707 = ~n63716;
  assign n63695 = n63719 & n63720;
  assign n63717 = ~n63715;
  assign n63341 = ~n62089;
  assign n63666 = ~n63691;
  assign n63671 = n63695 ^ n63696;
  assign n59827 = n63697 ^ n63698;
  assign n63640 = n63699 & n63700;
  assign n63684 = n63707 & n63708;
  assign n63702 = ~n63695;
  assign n63709 = n63717 & n63718;
  assign n63646 = n63671 ^ n63672;
  assign n63664 = n63684 ^ n63685;
  assign n63674 = n59827 & n61048;
  assign n63675 = n59827 & n62410;
  assign n63673 = n63640 & n63690;
  assign n59876 = ~n59827;
  assign n63680 = ~n63640;
  assign n63687 = ~n63684;
  assign n63692 = n63701 & n63702;
  assign n63703 = ~n63709;
  assign n63644 = n429 ^ n63664;
  assign n63652 = n63646 & n6946;
  assign n63653 = ~n63646;
  assign n63663 = ~n63673;
  assign n63657 = ~n63674;
  assign n62414 = ~n63675;
  assign n63668 = n59876 & n62359;
  assign n63669 = n59876 & n63676;
  assign n63667 = n63680 & n63655;
  assign n63683 = n63686 & n63687;
  assign n63681 = ~n63692;
  assign n63677 = n63703 & n63704;
  assign n62034 = n63643 ^ n63644;
  assign n63606 = n63644 & n63643;
  assign n63647 = ~n63652;
  assign n63650 = n63653 & n428;
  assign n63638 = ~n63667;
  assign n63656 = ~n63668;
  assign n62429 = ~n63669;
  assign n63659 = n63677 ^ n60991;
  assign n63654 = n63681 & n63682;
  assign n63665 = ~n63683;
  assign n63678 = ~n63677;
  assign n63315 = ~n62034;
  assign n63624 = ~n63650;
  assign n63641 = n63654 ^ n63655;
  assign n63601 = n63656 & n63657;
  assign n59752 = n63658 ^ n63659;
  assign n63645 = n63665 & n63666;
  assign n63662 = ~n63654;
  assign n63670 = n63678 & n63679;
  assign n63605 = n63640 ^ n63641;
  assign n63632 = n63601 & n63642;
  assign n63625 = n63645 ^ n63646;
  assign n63633 = n59752 & n62297;
  assign n63631 = n59752 & n63649;
  assign n63639 = ~n63601;
  assign n59773 = ~n59752;
  assign n63648 = ~n63645;
  assign n63651 = n63662 & n63663;
  assign n63660 = ~n63670;
  assign n63620 = n63605 & n427;
  assign n63607 = n428 ^ n63625;
  assign n63611 = ~n63605;
  assign n62396 = ~n63631;
  assign n63615 = ~n63632;
  assign n63627 = n59773 & n62375;
  assign n63621 = ~n63633;
  assign n63629 = n59773 & n61017;
  assign n63626 = n63639 & n63613;
  assign n63630 = n63647 & n63648;
  assign n63637 = ~n63651;
  assign n63634 = n63660 & n63661;
  assign n61975 = n63606 ^ n63607;
  assign n63565 = n63607 & n63606;
  assign n63610 = n63611 & n6920;
  assign n63571 = ~n63620;
  assign n63600 = ~n63626;
  assign n62374 = ~n63627;
  assign n63622 = ~n63629;
  assign n63623 = ~n63630;
  assign n63617 = n63634 ^ n60937;
  assign n63612 = n63637 & n63638;
  assign n63635 = ~n63634;
  assign n63271 = ~n61975;
  assign n63567 = ~n63565;
  assign n63597 = ~n63610;
  assign n63602 = n63612 ^ n63613;
  assign n59642 = n63616 ^ n63617;
  assign n63582 = n63621 & n63622;
  assign n63604 = n63623 & n63624;
  assign n63614 = ~n63612;
  assign n63628 = n63635 & n63636;
  assign n63564 = n63601 ^ n63602;
  assign n63592 = n63582 & n63548;
  assign n63596 = n59642 & n62258;
  assign n63584 = n63604 ^ n63605;
  assign n63603 = n59642 & n63608;
  assign n63590 = ~n63582;
  assign n59711 = ~n59642;
  assign n63609 = n63614 & n63615;
  assign n63598 = ~n63604;
  assign n63618 = ~n63628;
  assign n63572 = n63564 & n426;
  assign n63566 = n427 ^ n63584;
  assign n63583 = ~n63564;
  assign n63586 = n63590 & n63591;
  assign n63574 = ~n63592;
  assign n63575 = ~n63596;
  assign n63585 = n63597 & n63598;
  assign n63587 = n59711 & n62353;
  assign n62355 = ~n63603;
  assign n63589 = n59711 & n60937;
  assign n63599 = ~n63609;
  assign n63593 = n63618 & n63619;
  assign n61915 = n63565 ^ n63566;
  assign n63519 = n63566 & n63567;
  assign n63541 = ~n63572;
  assign n63568 = n63583 & n6878;
  assign n63570 = ~n63585;
  assign n63550 = ~n63586;
  assign n62338 = ~n63587;
  assign n63576 = ~n63589;
  assign n63577 = n63593 ^ n60902;
  assign n63581 = n63599 & n63600;
  assign n63594 = ~n63593;
  assign n63219 = ~n61915;
  assign n63560 = ~n63568;
  assign n63563 = n63570 & n63571;
  assign n63516 = n63575 & n63576;
  assign n59614 = n63577 ^ n63578;
  assign n63547 = n63581 ^ n63582;
  assign n63573 = ~n63581;
  assign n63588 = n63594 & n63595;
  assign n63508 = n63547 ^ n63548;
  assign n63527 = n63563 ^ n63564;
  assign n63552 = n63516 & n63530;
  assign n63551 = n59614 & n60888;
  assign n63562 = n59614 & n62305;
  assign n63559 = ~n63563;
  assign n63555 = ~n63516;
  assign n59621 = ~n59614;
  assign n63569 = n63573 & n63574;
  assign n63579 = ~n63588;
  assign n63520 = n426 ^ n63527;
  assign n63537 = n63508 & n6844;
  assign n63528 = ~n63508;
  assign n63538 = ~n63551;
  assign n63532 = ~n63552;
  assign n63542 = n63555 & n63556;
  assign n63544 = n59621 & n62203;
  assign n63546 = n63559 & n63560;
  assign n63543 = n59621 & n63561;
  assign n62303 = ~n63562;
  assign n63549 = ~n63569;
  assign n63553 = n63579 & n63580;
  assign n61880 = n63519 ^ n63520;
  assign n63474 = n63520 & n63519;
  assign n63525 = n63528 & n425;
  assign n63510 = ~n63537;
  assign n63522 = ~n63542;
  assign n62316 = ~n63543;
  assign n63539 = ~n63544;
  assign n63540 = ~n63546;
  assign n63529 = n63549 & n63550;
  assign n63536 = n63553 ^ n63554;
  assign n63557 = ~n63553;
  assign n63184 = ~n61880;
  assign n63501 = ~n63525;
  assign n63517 = n63529 ^ n63530;
  assign n59587 = n63536 ^ n60851;
  assign n63489 = n63538 & n63539;
  assign n63507 = n63540 & n63541;
  assign n63533 = n63536 & n60780;
  assign n63531 = ~n63529;
  assign n63545 = n63557 & n63558;
  assign n63498 = n63507 ^ n63508;
  assign n63477 = n63516 ^ n63517;
  assign n63512 = n63489 & n63523;
  assign n63511 = n59587 & n63524;
  assign n63509 = ~n63507;
  assign n63518 = ~n63489;
  assign n59529 = ~n59587;
  assign n63526 = n63531 & n63532;
  assign n63491 = ~n63533;
  assign n63534 = ~n63545;
  assign n63475 = n425 ^ n63498;
  assign n63487 = n63477 & n6815;
  assign n63499 = ~n63477;
  assign n63502 = n63509 & n63510;
  assign n62267 = ~n63511;
  assign n63493 = ~n63512;
  assign n63504 = n59529 & n62181;
  assign n63505 = n59529 & n62282;
  assign n63503 = n63518 & n63479;
  assign n63521 = ~n63526;
  assign n63513 = n63534 & n63535;
  assign n61764 = n63474 ^ n63475;
  assign n63482 = ~n63475;
  assign n63481 = ~n63487;
  assign n63485 = n63499 & n424;
  assign n63500 = ~n63502;
  assign n63466 = ~n63503;
  assign n63490 = ~n63504;
  assign n62279 = ~n63505;
  assign n63495 = n63513 ^ n60730;
  assign n63488 = n63521 & n63522;
  assign n63514 = ~n63513;
  assign n63134 = ~n61764;
  assign n63433 = n63482 & n63474;
  assign n63455 = ~n63485;
  assign n63478 = n63488 ^ n63489;
  assign n63436 = n63490 & n63491;
  assign n59504 = n63494 ^ n63495;
  assign n63476 = n63500 & n63501;
  assign n63492 = ~n63488;
  assign n63506 = n63514 & n63515;
  assign n63441 = ~n63433;
  assign n63459 = n63476 ^ n63477;
  assign n63424 = n63478 ^ n63479;
  assign n63468 = n59504 & n63483;
  assign n63470 = n59504 & n60748;
  assign n63469 = n63436 & n63484;
  assign n63480 = ~n63476;
  assign n63467 = ~n63436;
  assign n59545 = ~n59504;
  assign n63486 = n63492 & n63493;
  assign n63496 = ~n63506;
  assign n63434 = n424 ^ n63459;
  assign n63445 = n63424 & n439;
  assign n63456 = ~n63424;
  assign n63461 = n63467 & n63447;
  assign n62221 = ~n63468;
  assign n63452 = ~n63469;
  assign n63450 = ~n63470;
  assign n63463 = n59545 & n62222;
  assign n63462 = n59545 & n62108;
  assign n63460 = n63480 & n63481;
  assign n63465 = ~n63486;
  assign n63471 = n63496 & n63497;
  assign n61677 = n63433 ^ n63434;
  assign n63396 = n63434 & n63441;
  assign n63415 = ~n63445;
  assign n63443 = n63456 & n6709;
  assign n63454 = ~n63460;
  assign n63431 = ~n63461;
  assign n63451 = ~n63462;
  assign n62241 = ~n63463;
  assign n63446 = n63465 & n63466;
  assign n63458 = n63471 ^ n60649;
  assign n63472 = ~n63471;
  assign n63080 = ~n61677;
  assign n63439 = ~n63443;
  assign n63437 = n63446 ^ n63447;
  assign n63405 = n63450 & n63451;
  assign n63423 = n63454 & n63455;
  assign n59466 = n63457 ^ n63458;
  assign n63453 = ~n63446;
  assign n63464 = n63472 & n63473;
  assign n63413 = n63423 ^ n63424;
  assign n63393 = n63436 ^ n63437;
  assign n63427 = n59466 & n62182;
  assign n63425 = n63405 & n63442;
  assign n63426 = n59466 & n60698;
  assign n63438 = ~n63423;
  assign n59508 = ~n59466;
  assign n63435 = ~n63405;
  assign n63444 = n63452 & n63453;
  assign n63448 = ~n63464;
  assign n63399 = n439 ^ n63413;
  assign n63412 = n63393 & n438;
  assign n63403 = ~n63393;
  assign n63417 = ~n63425;
  assign n63411 = ~n63426;
  assign n62185 = ~n63427;
  assign n63420 = n59508 & n62100;
  assign n63418 = n63435 & n63398;
  assign n63422 = n63438 & n63439;
  assign n63419 = n59508 & n63440;
  assign n63430 = ~n63444;
  assign n63432 = n63448 & n63449;
  assign n61594 = n63396 ^ n63399;
  assign n63395 = ~n63399;
  assign n63401 = n63403 & n6678;
  assign n63365 = ~n63412;
  assign n63382 = ~n63418;
  assign n62199 = ~n63419;
  assign n63410 = ~n63420;
  assign n63414 = ~n63422;
  assign n63404 = n63430 & n63431;
  assign n63407 = n63432 ^ n60570;
  assign n63428 = ~n63432;
  assign n63001 = ~n61594;
  assign n63353 = n63395 & n63396;
  assign n63391 = ~n63401;
  assign n63397 = n63404 ^ n63405;
  assign n59424 = n63406 ^ n63407;
  assign n63354 = n63410 & n63411;
  assign n63392 = n63414 & n63415;
  assign n63416 = ~n63404;
  assign n63421 = n63428 & n63429;
  assign n63370 = n63392 ^ n63393;
  assign n63349 = n63397 ^ n63398;
  assign n63394 = n59424 & n63400;
  assign n63389 = n59424 & n62029;
  assign n63385 = n63354 & n63369;
  assign n63383 = ~n63354;
  assign n59455 = ~n59424;
  assign n63390 = ~n63392;
  assign n63402 = n63416 & n63417;
  assign n63408 = ~n63421;
  assign n63356 = n438 ^ n63370;
  assign n63361 = n63349 & n437;
  assign n63371 = ~n63349;
  assign n63377 = n63383 & n63384;
  assign n63379 = n59455 & n62138;
  assign n63367 = ~n63385;
  assign n63372 = ~n63389;
  assign n63376 = n63390 & n63391;
  assign n62160 = ~n63394;
  assign n63378 = n59455 & n60641;
  assign n63381 = ~n63402;
  assign n63386 = n63408 & n63409;
  assign n61563 = n63353 ^ n63356;
  assign n63352 = ~n63356;
  assign n63333 = ~n63361;
  assign n63359 = n63371 & n6625;
  assign n63364 = ~n63376;
  assign n63351 = ~n63377;
  assign n63373 = ~n63378;
  assign n62141 = ~n63379;
  assign n63368 = n63381 & n63382;
  assign n63375 = n63386 ^ n60488;
  assign n63387 = ~n63386;
  assign n62943 = ~n61563;
  assign n63311 = n63352 & n63353;
  assign n63358 = ~n63359;
  assign n63348 = n63364 & n63365;
  assign n63355 = n63368 ^ n63369;
  assign n63313 = n63372 & n63373;
  assign n59386 = n63374 ^ n63375;
  assign n63366 = ~n63368;
  assign n63380 = n63387 & n63388;
  assign n63328 = n63348 ^ n63349;
  assign n63298 = n63354 ^ n63355;
  assign n63343 = n63313 & n63321;
  assign n63344 = n59386 & n62089;
  assign n63342 = n59386 & n61986;
  assign n63357 = ~n63348;
  assign n63339 = ~n63313;
  assign n59411 = ~n59386;
  assign n63360 = n63366 & n63367;
  assign n63362 = ~n63380;
  assign n63312 = n437 ^ n63328;
  assign n63331 = n63298 & n6577;
  assign n63319 = ~n63298;
  assign n63335 = n63339 & n63340;
  assign n63336 = n59411 & n63341;
  assign n63338 = n59411 & n60546;
  assign n63329 = ~n63342;
  assign n63327 = ~n63343;
  assign n62114 = ~n63344;
  assign n63334 = n63357 & n63358;
  assign n63350 = ~n63360;
  assign n63345 = n63362 & n63363;
  assign n61430 = n63311 ^ n63312;
  assign n63310 = ~n63312;
  assign n63317 = n63319 & n436;
  assign n63304 = ~n63331;
  assign n63332 = ~n63334;
  assign n63306 = ~n63335;
  assign n62092 = ~n63336;
  assign n63330 = ~n63338;
  assign n63323 = n63345 ^ n60401;
  assign n63320 = n63350 & n63351;
  assign n63346 = ~n63345;
  assign n62880 = ~n61430;
  assign n63254 = n63310 & n63311;
  assign n63278 = ~n63317;
  assign n63314 = n63320 ^ n63321;
  assign n59347 = n63322 ^ n63323;
  assign n63256 = n63329 & n63330;
  assign n63297 = n63332 & n63333;
  assign n63326 = ~n63320;
  assign n63337 = n63346 & n63347;
  assign n63270 = ~n63254;
  assign n63285 = n63297 ^ n63298;
  assign n63273 = n63313 ^ n63314;
  assign n63299 = n59347 & n60401;
  assign n63301 = n59347 & n62034;
  assign n63309 = n63256 & n63316;
  assign n63302 = ~n63256;
  assign n59367 = ~n59347;
  assign n63303 = ~n63297;
  assign n63318 = n63326 & n63327;
  assign n63324 = ~n63337;
  assign n63255 = n436 ^ n63285;
  assign n63279 = n63273 & n6508;
  assign n63280 = ~n63273;
  assign n63294 = n59367 & n61939;
  assign n63286 = ~n63299;
  assign n62037 = ~n63301;
  assign n63296 = n63302 & n63282;
  assign n63292 = n63303 & n63304;
  assign n63291 = ~n63309;
  assign n63293 = n59367 & n63315;
  assign n63305 = ~n63318;
  assign n63300 = n63324 & n63325;
  assign n62827 = n63254 ^ n63255;
  assign n63269 = ~n63255;
  assign n63266 = ~n63279;
  assign n63275 = n63280 & n435;
  assign n63277 = ~n63292;
  assign n62068 = ~n63293;
  assign n63287 = ~n63294;
  assign n63264 = ~n63296;
  assign n63289 = n63300 ^ n60316;
  assign n63281 = n63305 & n63306;
  assign n63307 = ~n63300;
  assign n63222 = n63269 & n63270;
  assign n63248 = ~n63275;
  assign n63272 = n63277 & n63278;
  assign n63257 = n63281 ^ n63282;
  assign n63224 = n63286 & n63287;
  assign n59301 = n63288 ^ n63289;
  assign n63290 = ~n63281;
  assign n63295 = n63307 & n63308;
  assign n63230 = n63256 ^ n63257;
  assign n63243 = n63272 ^ n63273;
  assign n63258 = n59301 & n60384;
  assign n63259 = n63224 & n63245;
  assign n63274 = n59301 & n61975;
  assign n59327 = ~n59301;
  assign n63265 = ~n63272;
  assign n63267 = ~n63224;
  assign n63276 = n63290 & n63291;
  assign n63283 = ~n63295;
  assign n63223 = n435 ^ n63243;
  assign n63234 = n63230 & n434;
  assign n63246 = ~n63230;
  assign n63252 = n59327 & n61873;
  assign n63236 = ~n63258;
  assign n63238 = ~n63259;
  assign n63249 = n63265 & n63266;
  assign n63250 = n63267 & n63268;
  assign n63251 = n59327 & n63271;
  assign n61978 = ~n63274;
  assign n63263 = ~n63276;
  assign n63260 = n63283 & n63284;
  assign n63205 = n63222 ^ n63223;
  assign n63228 = ~n63223;
  assign n63190 = ~n63234;
  assign n63232 = n63246 & n6432;
  assign n63247 = ~n63249;
  assign n63221 = ~n63250;
  assign n62015 = ~n63251;
  assign n63235 = ~n63252;
  assign n63240 = n63260 ^ n60196;
  assign n63244 = n63263 & n63264;
  assign n63261 = ~n63260;
  assign n58974 = n63205 ^ n61004;
  assign n63086 = n63205 & n61004;
  assign n63204 = ~n63205;
  assign n63182 = n63228 & n63222;
  assign n63227 = ~n63232;
  assign n63171 = n63235 & n63236;
  assign n59240 = n63239 ^ n63240;
  assign n63225 = n63244 ^ n63245;
  assign n63229 = n63247 & n63248;
  assign n63237 = ~n63244;
  assign n63253 = n63261 & n63262;
  assign n58970 = ~n58974;
  assign n63187 = n63204 & n61004;
  assign n63179 = ~n63182;
  assign n63181 = n63224 ^ n63225;
  assign n63203 = n63229 ^ n63230;
  assign n63211 = n63171 & n63231;
  assign n63213 = n59240 & n61915;
  assign n63212 = n59240 & n60343;
  assign n63226 = ~n63229;
  assign n59286 = ~n59240;
  assign n63218 = ~n63171;
  assign n63233 = n63237 & n63238;
  assign n63241 = ~n63253;
  assign n63164 = n58970 & n62048;
  assign n63157 = ~n63187;
  assign n63183 = n434 ^ n63203;
  assign n63191 = n63181 & n6316;
  assign n63192 = ~n63181;
  assign n63196 = ~n63211;
  assign n63202 = ~n63212;
  assign n61914 = ~n63213;
  assign n63209 = n63218 & n63194;
  assign n63207 = n59286 & n61762;
  assign n63206 = n59286 & n63219;
  assign n63210 = n63226 & n63227;
  assign n63220 = ~n63233;
  assign n63214 = n63241 & n63242;
  assign n63156 = ~n63164;
  assign n63158 = n63182 ^ n63183;
  assign n63178 = ~n63183;
  assign n63176 = ~n63191;
  assign n63188 = n63192 & n433;
  assign n61945 = ~n63206;
  assign n63201 = ~n63207;
  assign n63174 = ~n63209;
  assign n63189 = ~n63210;
  assign n63197 = n63214 ^ n63215;
  assign n63193 = n63220 & n63221;
  assign n63216 = ~n63214;
  assign n63130 = n63156 & n63157;
  assign n63140 = n63158 & n60899;
  assign n63139 = ~n63158;
  assign n63132 = n63178 & n63179;
  assign n63142 = ~n63188;
  assign n63180 = n63189 & n63190;
  assign n63172 = n63193 ^ n63194;
  assign n59244 = n63197 ^ n60178;
  assign n63153 = n63201 & n63202;
  assign n63195 = ~n63193;
  assign n63198 = ~n63197;
  assign n63208 = n63216 & n63217;
  assign n63084 = n63130 ^ n63131;
  assign n63112 = ~n63130;
  assign n63136 = n63139 & n60904;
  assign n63105 = ~n63140;
  assign n63115 = n63171 ^ n63172;
  assign n63154 = n63180 ^ n63181;
  assign n63177 = n59244 & n63184;
  assign n63167 = n63153 & n63129;
  assign n63165 = ~n63153;
  assign n59220 = ~n59244;
  assign n63175 = ~n63180;
  assign n63185 = n63195 & n63196;
  assign n63186 = n63198 & n60178;
  assign n63199 = ~n63208;
  assign n60968 = n455 ^ n63084;
  assign n62800 = n63084 & n455;
  assign n62926 = n63112 & n63113;
  assign n63127 = ~n63136;
  assign n63133 = n433 ^ n63154;
  assign n63143 = n63115 & n432;
  assign n63155 = ~n63115;
  assign n63160 = n63165 & n63166;
  assign n63161 = n59220 & n61660;
  assign n63147 = ~n63167;
  assign n63162 = n59220 & n61880;
  assign n63159 = n63175 & n63176;
  assign n61836 = ~n63177;
  assign n63173 = ~n63185;
  assign n63145 = ~n63186;
  assign n63168 = n63199 & n63200;
  assign n62236 = ~n60968;
  assign n63085 = n63127 & n63105;
  assign n63106 = n63127 & n63086;
  assign n63048 = n63132 ^ n63133;
  assign n63076 = n63133 & n63132;
  assign n63101 = ~n63143;
  assign n63137 = n63155 & n6292;
  assign n63141 = ~n63159;
  assign n63124 = ~n63160;
  assign n63144 = ~n63161;
  assign n61878 = ~n63162;
  assign n63149 = n63168 ^ n60021;
  assign n63152 = n63173 & n63174;
  assign n63169 = ~n63168;
  assign n58927 = n63085 ^ n63086;
  assign n63088 = n63048 & n60847;
  assign n63104 = ~n63106;
  assign n63087 = ~n63048;
  assign n63079 = ~n63076;
  assign n63117 = ~n63137;
  assign n63114 = n63141 & n63142;
  assign n63074 = n63144 & n63145;
  assign n59175 = n63148 ^ n63149;
  assign n63128 = n63152 ^ n63153;
  assign n63146 = ~n63152;
  assign n63163 = n63169 & n63170;
  assign n63057 = n58927 & n60899;
  assign n58931 = ~n58927;
  assign n63081 = n63087 & n60817;
  assign n63040 = ~n63088;
  assign n63078 = n63104 & n63105;
  assign n63102 = n63114 ^ n63115;
  assign n63059 = n63128 ^ n63129;
  assign n63118 = n59175 & n63134;
  assign n63120 = n59175 & n61575;
  assign n63119 = n63074 & n63135;
  assign n63116 = ~n63114;
  assign n63122 = ~n63074;
  assign n59187 = ~n59175;
  assign n63138 = n63146 & n63147;
  assign n63150 = ~n63163;
  assign n63033 = ~n63057;
  assign n63050 = n58931 & n61956;
  assign n63049 = n63078 ^ n60817;
  assign n63073 = ~n63078;
  assign n63072 = ~n63081;
  assign n63077 = n432 ^ n63102;
  assign n63089 = n63059 & n6169;
  assign n63103 = ~n63059;
  assign n63107 = n63116 & n63117;
  assign n61800 = ~n63118;
  assign n63092 = ~n63119;
  assign n63109 = n59187 & n60021;
  assign n63096 = ~n63120;
  assign n63108 = n63122 & n63091;
  assign n63110 = n59187 & n61764;
  assign n63123 = ~n63138;
  assign n63121 = n63150 & n63151;
  assign n58893 = n63048 ^ n63049;
  assign n63034 = ~n63050;
  assign n63055 = n63072 & n63073;
  assign n62985 = n63076 ^ n63077;
  assign n63015 = n63077 & n63079;
  assign n63061 = ~n63089;
  assign n63082 = n63103 & n447;
  assign n63100 = ~n63107;
  assign n63063 = ~n63108;
  assign n63097 = ~n63109;
  assign n61767 = ~n63110;
  assign n63099 = n63121 ^ n59969;
  assign n63090 = n63123 & n63124;
  assign n63125 = ~n63121;
  assign n62995 = n58893 & n60847;
  assign n58903 = ~n58893;
  assign n63021 = n63033 & n63034;
  assign n63045 = n62985 & n60782;
  assign n63043 = ~n62985;
  assign n63039 = ~n63055;
  assign n63029 = ~n63082;
  assign n63075 = n63090 ^ n63091;
  assign n63008 = n63096 & n63097;
  assign n59117 = n63098 ^ n63099;
  assign n63058 = n63100 & n63101;
  assign n63093 = ~n63090;
  assign n63111 = n63125 & n63126;
  assign n62991 = n58903 & n61889;
  assign n62983 = ~n62995;
  assign n62996 = n63021 & n63022;
  assign n63019 = ~n63021;
  assign n62997 = n63039 & n63040;
  assign n63026 = n63043 & n60750;
  assign n62982 = ~n63045;
  assign n63027 = n63058 ^ n63059;
  assign n63011 = n63074 ^ n63075;
  assign n63069 = n59117 & n60043;
  assign n63066 = n59117 & n63080;
  assign n63067 = n63008 & n63047;
  assign n63064 = ~n63008;
  assign n59161 = ~n59117;
  assign n63060 = ~n63058;
  assign n63083 = n63092 & n63093;
  assign n63094 = ~n63111;
  assign n62984 = ~n62991;
  assign n62963 = ~n62996;
  assign n62986 = n62997 ^ n60750;
  assign n62994 = n63019 & n63020;
  assign n63013 = ~n62997;
  assign n63012 = ~n63026;
  assign n63016 = n447 ^ n63027;
  assign n63030 = n63011 & n446;
  assign n63044 = ~n63011;
  assign n63056 = n63060 & n63061;
  assign n63051 = n63064 & n63065;
  assign n61680 = ~n63066;
  assign n63053 = n59161 & n61677;
  assign n63042 = ~n63067;
  assign n63035 = ~n63069;
  assign n63052 = n59161 & n61491;
  assign n63062 = ~n63083;
  assign n63068 = n63094 & n63095;
  assign n62882 = n62983 & n62984;
  assign n58862 = n62985 ^ n62986;
  assign n62962 = n62963 & n62926;
  assign n62956 = ~n62994;
  assign n62992 = n63012 & n63013;
  assign n62890 = n63015 ^ n63016;
  assign n63014 = ~n63016;
  assign n62968 = ~n63030;
  assign n63024 = n63044 & n6144;
  assign n62999 = ~n63051;
  assign n63036 = ~n63052;
  assign n61725 = ~n63053;
  assign n63028 = ~n63056;
  assign n63046 = n63062 & n63063;
  assign n63038 = n63068 ^ n59885;
  assign n63070 = ~n63068;
  assign n62930 = n58862 & n60782;
  assign n62929 = n62882 & n62957;
  assign n62928 = ~n62882;
  assign n58878 = ~n58862;
  assign n62955 = ~n62962;
  assign n62958 = n62956 & n62963;
  assign n62965 = n62890 & n60656;
  assign n62964 = ~n62890;
  assign n62981 = ~n62992;
  assign n62949 = n63014 & n63015;
  assign n63017 = ~n63024;
  assign n63010 = n63028 & n63029;
  assign n62938 = n63035 & n63036;
  assign n59090 = n63037 ^ n63038;
  assign n63009 = n63046 ^ n63047;
  assign n63041 = ~n63046;
  assign n63054 = n63070 & n63071;
  assign n62918 = n62928 & n62915;
  assign n62916 = ~n62929;
  assign n62906 = ~n62930;
  assign n62919 = n58878 & n61811;
  assign n62914 = n62955 & n62956;
  assign n62927 = ~n62958;
  assign n62959 = n62964 & n60667;
  assign n62909 = ~n62965;
  assign n62931 = n62981 & n62982;
  assign n62935 = ~n62949;
  assign n62937 = n63008 ^ n63009;
  assign n62966 = n63010 ^ n63011;
  assign n63007 = n59090 & n61594;
  assign n63002 = n59090 & n61470;
  assign n63003 = n62938 & n63023;
  assign n63018 = ~n63010;
  assign n59114 = ~n59090;
  assign n63000 = ~n62938;
  assign n63025 = n63041 & n63042;
  assign n63031 = ~n63054;
  assign n62883 = n62914 ^ n62915;
  assign n62878 = ~n62918;
  assign n62907 = ~n62919;
  assign n62911 = n62926 ^ n62927;
  assign n62917 = ~n62914;
  assign n62891 = n62931 ^ n60656;
  assign n62932 = ~n62959;
  assign n62933 = ~n62931;
  assign n62950 = n446 ^ n62966;
  assign n62969 = n62937 & n6018;
  assign n62970 = ~n62937;
  assign n62990 = n63000 & n62972;
  assign n62989 = n59114 & n63001;
  assign n62978 = ~n63002;
  assign n62974 = ~n63003;
  assign n62987 = n59114 & n59885;
  assign n61648 = ~n63007;
  assign n62993 = n63017 & n63018;
  assign n62998 = ~n63025;
  assign n63004 = n63031 & n63032;
  assign n62797 = n62882 ^ n62883;
  assign n58827 = n62890 ^ n62891;
  assign n62803 = n62906 & n62907;
  assign n62884 = n62911 & n18650;
  assign n62888 = ~n62911;
  assign n62889 = n62916 & n62917;
  assign n62924 = n62932 & n62933;
  assign n62810 = n62949 ^ n62950;
  assign n62934 = ~n62950;
  assign n62951 = ~n62969;
  assign n62960 = n62970 & n445;
  assign n62977 = ~n62987;
  assign n61597 = ~n62989;
  assign n62941 = ~n62990;
  assign n62967 = ~n62993;
  assign n62971 = n62998 & n62999;
  assign n62980 = n63004 ^ n59806;
  assign n63005 = ~n63004;
  assign n62842 = n62797 & n453;
  assign n62835 = ~n62797;
  assign n62875 = n58827 & n61713;
  assign n62876 = n62803 & n62837;
  assign n62844 = ~n62884;
  assign n62852 = ~n62803;
  assign n58829 = ~n58827;
  assign n62879 = n62888 & n454;
  assign n62877 = ~n62889;
  assign n62893 = n62810 & n60556;
  assign n62892 = ~n62810;
  assign n62908 = ~n62924;
  assign n62871 = n62934 & n62935;
  assign n62913 = ~n62960;
  assign n62936 = n62967 & n62968;
  assign n62939 = n62971 ^ n62972;
  assign n62859 = n62977 & n62978;
  assign n59050 = n62979 ^ n62980;
  assign n62973 = ~n62971;
  assign n62988 = n63005 & n63006;
  assign n62828 = n62835 & n18542;
  assign n62764 = ~n62842;
  assign n62850 = n62852 & n62853;
  assign n62843 = n62844 & n62800;
  assign n62845 = n58829 & n60656;
  assign n62832 = ~n62875;
  assign n62839 = ~n62876;
  assign n62836 = n62877 & n62878;
  assign n62830 = ~n62879;
  assign n62885 = n62892 & n60590;
  assign n62813 = ~n62893;
  assign n62854 = n62908 & n62909;
  assign n62870 = ~n62871;
  assign n62894 = n62936 ^ n62937;
  assign n62856 = n62938 ^ n62939;
  assign n62942 = n59050 & n61415;
  assign n62947 = n59050 & n61563;
  assign n62953 = n62859 & n62954;
  assign n59070 = ~n59050;
  assign n62948 = ~n62859;
  assign n62952 = ~n62936;
  assign n62961 = n62973 & n62974;
  assign n62975 = ~n62988;
  assign n62777 = ~n62828;
  assign n62804 = n62836 ^ n62837;
  assign n62829 = ~n62843;
  assign n62841 = n62844 & n62830;
  assign n62833 = ~n62845;
  assign n62799 = ~n62850;
  assign n62811 = n62854 ^ n60556;
  assign n62840 = ~n62836;
  assign n62874 = ~n62885;
  assign n62873 = ~n62854;
  assign n62872 = n445 ^ n62894;
  assign n62910 = n62856 & n444;
  assign n62895 = ~n62856;
  assign n62904 = ~n62942;
  assign n62923 = n59070 & n62943;
  assign n62921 = n59070 & n59866;
  assign n61561 = ~n62947;
  assign n62920 = n62948 & n62897;
  assign n62925 = n62951 & n62952;
  assign n62899 = ~n62953;
  assign n62940 = ~n62961;
  assign n62944 = n62975 & n62976;
  assign n62728 = n62803 ^ n62804;
  assign n58783 = n62810 ^ n62811;
  assign n62796 = n62829 & n62830;
  assign n62735 = n62832 & n62833;
  assign n62809 = n62839 & n62840;
  assign n62801 = ~n62841;
  assign n62838 = n62871 ^ n62872;
  assign n62846 = n62873 & n62874;
  assign n62869 = ~n62872;
  assign n62886 = n62895 & n5930;
  assign n62817 = ~n62910;
  assign n62866 = ~n62920;
  assign n62905 = ~n62921;
  assign n61517 = ~n62923;
  assign n62912 = ~n62925;
  assign n62896 = n62940 & n62941;
  assign n62901 = n62944 ^ n59733;
  assign n62945 = ~n62944;
  assign n62765 = n62728 & n18500;
  assign n62770 = ~n62728;
  assign n62760 = n62796 ^ n62797;
  assign n62781 = n58783 & n61633;
  assign n60852 = n62800 ^ n62801;
  assign n62780 = n62735 & n62802;
  assign n62779 = ~n62735;
  assign n62778 = ~n62796;
  assign n58791 = ~n58783;
  assign n62798 = ~n62809;
  assign n62814 = n62838 & n60516;
  assign n62812 = ~n62846;
  assign n62831 = ~n62838;
  assign n62784 = n62869 & n62870;
  assign n62858 = ~n62886;
  assign n62860 = n62896 ^ n62897;
  assign n59014 = n62900 ^ n62901;
  assign n62786 = n62904 & n62905;
  assign n62855 = n62912 & n62913;
  assign n62898 = ~n62896;
  assign n62922 = n62945 & n62946;
  assign n62711 = n453 ^ n62760;
  assign n62712 = ~n62765;
  assign n62761 = n62770 & n452;
  assign n62775 = n62777 & n62778;
  assign n62771 = n62779 & n62769;
  assign n62766 = ~n62780;
  assign n62742 = ~n62781;
  assign n62772 = n58791 & n60556;
  assign n62768 = n62798 & n62799;
  assign n62740 = n62812 & n62813;
  assign n62783 = ~n62814;
  assign n62805 = n62831 & n60452;
  assign n62815 = n62855 ^ n62856;
  assign n62795 = n62859 ^ n62860;
  assign n62864 = n59014 & n59783;
  assign n62862 = n59014 & n62880;
  assign n62863 = n62786 & n62881;
  assign n62861 = ~n62786;
  assign n59039 = ~n59014;
  assign n62857 = ~n62855;
  assign n62887 = n62898 & n62899;
  assign n62902 = ~n62922;
  assign n60812 = n62711 ^ n60852;
  assign n62669 = n62711 & n60852;
  assign n62696 = ~n62761;
  assign n62736 = n62768 ^ n62769;
  assign n62731 = ~n62771;
  assign n62743 = ~n62772;
  assign n62763 = ~n62775;
  assign n62767 = ~n62768;
  assign n62782 = ~n62740;
  assign n62759 = ~n62805;
  assign n62785 = n444 ^ n62815;
  assign n62834 = n62795 & n443;
  assign n62818 = ~n62795;
  assign n62851 = n62857 & n62858;
  assign n62847 = n62861 & n62820;
  assign n61494 = ~n62862;
  assign n62822 = ~n62863;
  assign n62825 = ~n62864;
  assign n62849 = n59039 & n61322;
  assign n62848 = n59039 & n61430;
  assign n62865 = ~n62887;
  assign n62867 = n62902 & n62903;
  assign n62161 = ~n60812;
  assign n62667 = n62735 ^ n62736;
  assign n62675 = n62742 & n62743;
  assign n62727 = n62763 & n62764;
  assign n62762 = n62766 & n62767;
  assign n62774 = n62782 & n62783;
  assign n62776 = n62783 & n62759;
  assign n62684 = n62784 ^ n62785;
  assign n62718 = n62785 & n62784;
  assign n62808 = n62818 & n5860;
  assign n62756 = ~n62834;
  assign n62789 = ~n62847;
  assign n61447 = ~n62848;
  assign n62826 = ~n62849;
  assign n62816 = ~n62851;
  assign n62819 = n62865 & n62866;
  assign n58994 = n62867 ^ n62868;
  assign n62702 = n62667 & n451;
  assign n62705 = ~n62667;
  assign n62681 = n62727 ^ n62728;
  assign n62715 = n62675 & n62732;
  assign n62714 = ~n62675;
  assign n62713 = ~n62727;
  assign n62730 = ~n62762;
  assign n62744 = n62684 & n60432;
  assign n62757 = ~n62684;
  assign n62758 = ~n62774;
  assign n62741 = ~n62776;
  assign n62793 = ~n62808;
  assign n62794 = n62816 & n62817;
  assign n62787 = n62819 ^ n62820;
  assign n62720 = n62825 & n62826;
  assign n61413 = n62827 ^ n58994;
  assign n62823 = n58994 & n59709;
  assign n62821 = ~n62819;
  assign n59786 = ~n58994;
  assign n62670 = n452 ^ n62681;
  assign n62625 = ~n62702;
  assign n62682 = n62705 & n18450;
  assign n62706 = n62712 & n62713;
  assign n62707 = n62714 & n62698;
  assign n62703 = ~n62715;
  assign n62697 = n62730 & n62731;
  assign n58749 = n62740 ^ n62741;
  assign n62717 = ~n62744;
  assign n62737 = n62757 & n60370;
  assign n62729 = n62758 & n62759;
  assign n62724 = n62786 ^ n62787;
  assign n62745 = n62794 ^ n62795;
  assign n62792 = ~n62794;
  assign n62734 = ~n62720;
  assign n62806 = n62821 & n62822;
  assign n62791 = ~n62823;
  assign n62807 = n59786 & n62824;
  assign n60778 = n62669 ^ n62670;
  assign n62671 = ~n62670;
  assign n62655 = ~n62682;
  assign n62676 = n62697 ^ n62698;
  assign n62695 = ~n62706;
  assign n62673 = ~n62707;
  assign n62710 = n58749 & n60452;
  assign n62704 = ~n62697;
  assign n62685 = n62729 ^ n60370;
  assign n58757 = ~n58749;
  assign n62716 = ~n62729;
  assign n62687 = ~n62737;
  assign n62719 = n443 ^ n62745;
  assign n62747 = n62724 & n442;
  assign n62746 = ~n62724;
  assign n62773 = n62792 & n62793;
  assign n62788 = ~n62806;
  assign n62790 = ~n62807;
  assign n62115 = ~n60778;
  assign n62598 = n62671 & n62669;
  assign n62615 = n62675 ^ n62676;
  assign n58700 = n62684 ^ n62685;
  assign n62666 = n62695 & n62696;
  assign n62683 = n62703 & n62704;
  assign n62699 = n58757 & n61546;
  assign n62677 = ~n62710;
  assign n62708 = n62716 & n62717;
  assign n62632 = n62718 ^ n62719;
  assign n62660 = n62719 & n62718;
  assign n62738 = n62746 & n5793;
  assign n62692 = ~n62747;
  assign n62755 = ~n62773;
  assign n62748 = n62788 & n62789;
  assign n62753 = n62790 & n62791;
  assign n62619 = ~n62598;
  assign n62642 = n62615 & n450;
  assign n62634 = n62666 ^ n62667;
  assign n62641 = ~n62615;
  assign n62668 = n58700 & n60370;
  assign n62654 = ~n62666;
  assign n58719 = ~n58700;
  assign n62672 = ~n62683;
  assign n62678 = ~n62699;
  assign n62689 = n62632 & n60325;
  assign n62688 = ~n62632;
  assign n62686 = ~n62708;
  assign n62726 = ~n62738;
  assign n62721 = n62748 ^ n62749;
  assign n62647 = n62753 ^ n62754;
  assign n62723 = n62755 & n62756;
  assign n62752 = n62748 & n62749;
  assign n62750 = ~n62748;
  assign n62599 = n451 ^ n62634;
  assign n62639 = n62641 & n18410;
  assign n62590 = ~n62642;
  assign n62652 = n62654 & n62655;
  assign n62648 = n58719 & n61451;
  assign n62636 = ~n62668;
  assign n62643 = n62672 & n62673;
  assign n62620 = n62677 & n62678;
  assign n62657 = n62686 & n62687;
  assign n62680 = n62688 & n60290;
  assign n62658 = ~n62689;
  assign n62663 = n62720 ^ n62721;
  assign n62690 = n62723 ^ n62724;
  assign n62725 = ~n62723;
  assign n62739 = n62750 & n62751;
  assign n62733 = ~n62752;
  assign n60661 = n62598 ^ n62599;
  assign n62618 = ~n62599;
  assign n62616 = ~n62639;
  assign n62621 = n62643 ^ n62644;
  assign n62635 = ~n62648;
  assign n62624 = ~n62652;
  assign n62649 = n62620 & n62656;
  assign n62633 = n62657 ^ n60290;
  assign n62637 = ~n62643;
  assign n62653 = ~n62620;
  assign n62659 = ~n62657;
  assign n62631 = ~n62680;
  assign n62661 = n442 ^ n62690;
  assign n62693 = n62663 & n5708;
  assign n62694 = ~n62663;
  assign n62709 = n62725 & n62726;
  assign n62722 = n62733 & n62734;
  assign n62701 = ~n62739;
  assign n62079 = ~n60661;
  assign n62553 = n62618 & n62619;
  assign n62555 = n62620 ^ n62621;
  assign n62614 = n62624 & n62625;
  assign n58665 = n62632 ^ n62633;
  assign n62562 = n62635 & n62636;
  assign n62638 = ~n62649;
  assign n62645 = n62653 & n62644;
  assign n62651 = n62658 & n62659;
  assign n62579 = n62660 ^ n62661;
  assign n62610 = n62661 & n62660;
  assign n62665 = ~n62693;
  assign n62679 = n62694 & n441;
  assign n62691 = ~n62709;
  assign n62700 = ~n62722;
  assign n62593 = n62555 & n449;
  assign n62592 = ~n62555;
  assign n62591 = n62614 ^ n62615;
  assign n62604 = n58665 & n60290;
  assign n62605 = n62562 & n62588;
  assign n62602 = ~n62562;
  assign n58678 = ~n58665;
  assign n62617 = ~n62614;
  assign n62622 = n62637 & n62638;
  assign n62601 = ~n62645;
  assign n62627 = n62579 & n60243;
  assign n62626 = ~n62579;
  assign n62630 = ~n62651;
  assign n62629 = ~n62679;
  assign n62662 = n62691 & n62692;
  assign n62674 = n62700 & n62701;
  assign n62569 = n450 ^ n62591;
  assign n62576 = n62592 & n18389;
  assign n62536 = ~n62593;
  assign n62595 = n62602 & n62603;
  assign n62596 = n58678 & n61405;
  assign n62577 = ~n62604;
  assign n62575 = ~n62605;
  assign n62597 = n62616 & n62617;
  assign n62600 = ~n62622;
  assign n62623 = n62626 & n60184;
  assign n62608 = ~n62627;
  assign n62606 = n62630 & n62631;
  assign n62640 = n62662 ^ n62663;
  assign n62646 = n440 ^ n62674;
  assign n62664 = ~n62662;
  assign n60628 = n62553 ^ n62569;
  assign n62552 = ~n62569;
  assign n62570 = ~n62576;
  assign n62565 = ~n62595;
  assign n62578 = ~n62596;
  assign n62589 = ~n62597;
  assign n62587 = n62600 & n62601;
  assign n62580 = n62606 ^ n60184;
  assign n62607 = ~n62606;
  assign n62582 = ~n62623;
  assign n62613 = n441 ^ n62640;
  assign n62612 = n62646 ^ n62647;
  assign n62650 = n62664 & n62665;
  assign n62009 = ~n60628;
  assign n62512 = n62552 & n62553;
  assign n62524 = n62577 & n62578;
  assign n58617 = n62579 ^ n62580;
  assign n62563 = n62587 ^ n62588;
  assign n62554 = n62589 & n62590;
  assign n62574 = ~n62587;
  assign n62594 = n62607 & n62608;
  assign n62532 = n62610 ^ n62613;
  assign n62609 = ~n62613;
  assign n62628 = ~n62650;
  assign n62534 = n62554 ^ n62555;
  assign n62515 = n62562 ^ n62563;
  assign n62557 = n62524 & n62539;
  assign n62556 = n58617 & n60184;
  assign n62571 = ~n62554;
  assign n62567 = ~n62524;
  assign n58648 = ~n58617;
  assign n62573 = n62574 & n62575;
  assign n62584 = n62532 & n60093;
  assign n62581 = ~n62594;
  assign n62583 = ~n62532;
  assign n62585 = n62609 & n62610;
  assign n62611 = n62628 & n62629;
  assign n62513 = n449 ^ n62534;
  assign n62546 = n62515 & n18335;
  assign n62537 = ~n62515;
  assign n62548 = n58648 & n61289;
  assign n62542 = ~n62556;
  assign n62545 = ~n62557;
  assign n62551 = n62567 & n62568;
  assign n62547 = n62570 & n62571;
  assign n62564 = ~n62573;
  assign n62558 = n62581 & n62582;
  assign n62572 = n62583 & n60142;
  assign n62541 = ~n62584;
  assign n62586 = n62611 ^ n62612;
  assign n60506 = n62512 ^ n62513;
  assign n62526 = ~n62513;
  assign n62531 = n62537 & n448;
  assign n62527 = ~n62546;
  assign n62535 = ~n62547;
  assign n62543 = ~n62548;
  assign n62522 = ~n62551;
  assign n62533 = n62558 ^ n60093;
  assign n62538 = n62564 & n62565;
  assign n62559 = ~n62558;
  assign n62560 = ~n62572;
  assign n62500 = n62585 ^ n62586;
  assign n61948 = ~n60506;
  assign n62486 = n62526 & n62512;
  assign n62507 = ~n62531;
  assign n58579 = n62532 ^ n62533;
  assign n62514 = n62535 & n62536;
  assign n62525 = n62538 ^ n62539;
  assign n62484 = n62542 & n62543;
  assign n62544 = ~n62538;
  assign n62550 = n62559 & n62560;
  assign n62566 = n62500 & n60032;
  assign n62561 = ~n62500;
  assign n62473 = ~n62486;
  assign n62505 = n62514 ^ n62515;
  assign n62475 = n62524 ^ n62525;
  assign n62516 = n62484 & n62529;
  assign n62517 = n58579 & n61233;
  assign n62523 = ~n62484;
  assign n58588 = ~n58579;
  assign n62528 = ~n62514;
  assign n62530 = n62544 & n62545;
  assign n62540 = ~n62550;
  assign n62549 = n62561 & n60051;
  assign n62520 = ~n62566;
  assign n62487 = n448 ^ n62505;
  assign n62493 = n62475 & n18294;
  assign n62502 = ~n62475;
  assign n62497 = ~n62516;
  assign n62510 = n58588 & n60093;
  assign n62498 = ~n62517;
  assign n62509 = n62523 & n62495;
  assign n62508 = n62527 & n62528;
  assign n62521 = ~n62530;
  assign n62518 = n62540 & n62541;
  assign n62504 = ~n62549;
  assign n61896 = n62486 ^ n62487;
  assign n62472 = ~n62487;
  assign n62483 = ~n62493;
  assign n62491 = n62502 & n463;
  assign n62506 = ~n62508;
  assign n62489 = ~n62509;
  assign n62499 = ~n62510;
  assign n62501 = n62518 ^ n60032;
  assign n62494 = n62521 & n62522;
  assign n62519 = ~n62518;
  assign n61885 = ~n61896;
  assign n62436 = n62472 & n62473;
  assign n62465 = ~n62491;
  assign n62485 = n62494 ^ n62495;
  assign n62439 = n62498 & n62499;
  assign n58531 = n62500 ^ n62501;
  assign n62474 = n62506 & n62507;
  assign n62496 = ~n62494;
  assign n62511 = n62519 & n62520;
  assign n62454 = n62474 ^ n62475;
  assign n62438 = n62484 ^ n62485;
  assign n62476 = n58531 & n61156;
  assign n62477 = n62439 & n62458;
  assign n62480 = ~n62439;
  assign n58566 = ~n58531;
  assign n62482 = ~n62474;
  assign n62492 = n62496 & n62497;
  assign n62503 = ~n62511;
  assign n62448 = n463 ^ n62454;
  assign n62456 = n62438 & n462;
  assign n62455 = ~n62438;
  assign n62463 = ~n62476;
  assign n62461 = ~n62477;
  assign n62469 = n58566 & n60051;
  assign n62468 = n62480 & n62481;
  assign n62471 = n62482 & n62483;
  assign n62488 = ~n62492;
  assign n62490 = n62503 & n62504;
  assign n60382 = n62436 ^ n62448;
  assign n62435 = ~n62448;
  assign n62451 = n62455 & n18263;
  assign n62420 = ~n62456;
  assign n62445 = ~n62468;
  assign n62462 = ~n62469;
  assign n62464 = ~n62471;
  assign n62457 = n62488 & n62489;
  assign n62479 = n62490 & n59961;
  assign n62478 = ~n62490;
  assign n61804 = ~n60382;
  assign n62406 = n62435 & n62436;
  assign n62447 = ~n62451;
  assign n62440 = n62457 ^ n62458;
  assign n62408 = n62462 & n62463;
  assign n62437 = n62464 & n62465;
  assign n62460 = ~n62457;
  assign n62470 = n62478 & n59922;
  assign n62459 = ~n62479;
  assign n62418 = n62437 ^ n62438;
  assign n62401 = n62439 ^ n62440;
  assign n62441 = n62408 & n62425;
  assign n62442 = ~n62408;
  assign n62446 = ~n62437;
  assign n62453 = n62460 & n62461;
  assign n62466 = n62459 & n62467;
  assign n62450 = ~n62470;
  assign n62407 = n462 ^ n62418;
  assign n62426 = n62401 & n18218;
  assign n62427 = ~n62401;
  assign n62422 = ~n62441;
  assign n62432 = n62442 & n62443;
  assign n62431 = n62446 & n62447;
  assign n62444 = ~n62453;
  assign n62452 = n62450 & n62459;
  assign n62449 = ~n62466;
  assign n60247 = n62406 ^ n62407;
  assign n62361 = n62407 & n62406;
  assign n62405 = ~n62426;
  assign n62415 = n62427 & n461;
  assign n62419 = ~n62431;
  assign n62403 = ~n62432;
  assign n62424 = n62444 & n62445;
  assign n62430 = n62449 & n62450;
  assign n62433 = ~n62452;
  assign n61741 = ~n60247;
  assign n62370 = ~n62361;
  assign n62391 = ~n62415;
  assign n62400 = n62419 & n62420;
  assign n62409 = n62424 ^ n62425;
  assign n62411 = n62430 ^ n59827;
  assign n62421 = ~n62424;
  assign n58492 = n62433 ^ n62434;
  assign n62428 = ~n62430;
  assign n62392 = n62400 ^ n62401;
  assign n62364 = n62408 ^ n62409;
  assign n58444 = n62410 ^ n62411;
  assign n62404 = ~n62400;
  assign n62416 = n62421 & n62422;
  assign n62417 = n58492 & n59922;
  assign n62423 = n62428 & n62429;
  assign n58501 = ~n58492;
  assign n62362 = n461 ^ n62392;
  assign n62381 = n62364 & n18199;
  assign n62387 = ~n62364;
  assign n62393 = n58444 & n61048;
  assign n58495 = ~n58444;
  assign n62399 = n62404 & n62405;
  assign n62402 = ~n62416;
  assign n62412 = n58501 & n61084;
  assign n62397 = ~n62417;
  assign n62413 = ~n62423;
  assign n60162 = n62361 ^ n62362;
  assign n62327 = n62362 & n62370;
  assign n62369 = ~n62381;
  assign n62380 = n62387 & n460;
  assign n62384 = n58495 & n59827;
  assign n62371 = ~n62393;
  assign n62390 = ~n62399;
  assign n62388 = n62402 & n62403;
  assign n62398 = ~n62412;
  assign n62394 = n62413 & n62414;
  assign n61661 = ~n60162;
  assign n62349 = ~n62380;
  assign n62372 = ~n62384;
  assign n62367 = n62388 ^ n62389;
  assign n62363 = n62390 & n62391;
  assign n62386 = n62388 & n62389;
  assign n62376 = n62394 ^ n59752;
  assign n62382 = ~n62388;
  assign n62366 = n62397 & n62398;
  assign n62395 = ~n62394;
  assign n62347 = n62363 ^ n62364;
  assign n62325 = n62366 ^ n62367;
  assign n62320 = n62371 & n62372;
  assign n58399 = n62375 ^ n62376;
  assign n62368 = ~n62363;
  assign n62379 = n62382 & n62383;
  assign n62377 = ~n62386;
  assign n62385 = n62395 & n62396;
  assign n62378 = ~n62366;
  assign n62328 = n460 ^ n62347;
  assign n62342 = n62325 & n18144;
  assign n62343 = ~n62325;
  assign n62351 = n62320 & n62332;
  assign n62350 = n58399 & n59773;
  assign n62358 = ~n62320;
  assign n58419 = ~n58399;
  assign n62360 = n62368 & n62369;
  assign n62365 = n62377 & n62378;
  assign n62357 = ~n62379;
  assign n62373 = ~n62385;
  assign n60079 = n62327 ^ n62328;
  assign n62293 = n62328 & n62327;
  assign n62330 = ~n62342;
  assign n62341 = n62343 & n459;
  assign n62333 = ~n62350;
  assign n62340 = ~n62351;
  assign n62344 = n62358 & n62359;
  assign n62346 = n58419 & n61017;
  assign n62348 = ~n62360;
  assign n62356 = ~n62365;
  assign n62352 = n62373 & n62374;
  assign n61578 = ~n60079;
  assign n62312 = ~n62341;
  assign n62319 = ~n62344;
  assign n62334 = ~n62346;
  assign n62324 = n62348 & n62349;
  assign n62335 = n62352 ^ n62353;
  assign n62331 = n62356 & n62357;
  assign n62354 = ~n62352;
  assign n62307 = n62324 ^ n62325;
  assign n62321 = n62331 ^ n62332;
  assign n62274 = n62333 & n62334;
  assign n58350 = n59642 ^ n62335;
  assign n62329 = ~n62324;
  assign n62336 = n62335 & n59711;
  assign n62339 = ~n62331;
  assign n62345 = n62354 & n62355;
  assign n62294 = n459 ^ n62307;
  assign n62292 = n62320 ^ n62321;
  assign n62313 = n62274 & n62323;
  assign n62317 = ~n62274;
  assign n58423 = ~n58350;
  assign n62322 = n62329 & n62330;
  assign n62301 = ~n62336;
  assign n62326 = n62339 & n62340;
  assign n62337 = ~n62345;
  assign n59992 = n62293 ^ n62294;
  assign n62251 = n62294 & n62293;
  assign n62295 = n62292 & n18124;
  assign n62304 = ~n62292;
  assign n62299 = ~n62313;
  assign n62310 = n58423 & n60937;
  assign n62308 = n62317 & n62297;
  assign n62311 = ~n62322;
  assign n62318 = ~n62326;
  assign n62314 = n62337 & n62338;
  assign n61495 = ~n59992;
  assign n62287 = ~n62295;
  assign n62289 = n62304 & n458;
  assign n62285 = ~n62308;
  assign n62300 = ~n62310;
  assign n62291 = n62311 & n62312;
  assign n62306 = n62314 ^ n59614;
  assign n62296 = n62318 & n62319;
  assign n62315 = ~n62314;
  assign n62269 = ~n62289;
  assign n62273 = n62291 ^ n62292;
  assign n62275 = n62296 ^ n62297;
  assign n62242 = n62300 & n62301;
  assign n58324 = n62305 ^ n62306;
  assign n62288 = ~n62291;
  assign n62298 = ~n62296;
  assign n62309 = n62315 & n62316;
  assign n62252 = n458 ^ n62273;
  assign n62249 = n62274 ^ n62275;
  assign n62283 = n58324 & n60888;
  assign n62277 = n62242 & n62286;
  assign n62280 = n62287 & n62288;
  assign n62276 = ~n62242;
  assign n58321 = ~n58324;
  assign n62290 = n62298 & n62299;
  assign n62302 = ~n62309;
  assign n59902 = n62251 ^ n62252;
  assign n62209 = n62252 & n62251;
  assign n62263 = n62249 & n457;
  assign n62256 = ~n62249;
  assign n62270 = n62276 & n62258;
  assign n62264 = ~n62277;
  assign n62268 = ~n62280;
  assign n62271 = n58321 & n59614;
  assign n62259 = ~n62283;
  assign n62284 = ~n62290;
  assign n62281 = n62302 & n62303;
  assign n61395 = ~n59902;
  assign n62212 = ~n62209;
  assign n62253 = n62256 & n18059;
  assign n62225 = ~n62263;
  assign n62248 = n62268 & n62269;
  assign n62247 = ~n62270;
  assign n62260 = ~n62271;
  assign n62261 = n62281 ^ n62282;
  assign n62257 = n62284 & n62285;
  assign n62278 = ~n62281;
  assign n62229 = n62248 ^ n62249;
  assign n62244 = ~n62253;
  assign n62243 = n62257 ^ n62258;
  assign n62217 = n62259 & n62260;
  assign n58249 = n59587 ^ n62261;
  assign n62245 = ~n62248;
  assign n62262 = ~n62261;
  assign n62265 = ~n62257;
  assign n62272 = n62278 & n62279;
  assign n62210 = n457 ^ n62229;
  assign n62205 = n62242 ^ n62243;
  assign n62230 = n62244 & n62245;
  assign n62239 = n62217 & n62250;
  assign n62237 = n58249 & n60968;
  assign n62235 = ~n62217;
  assign n58347 = ~n58249;
  assign n62255 = n62262 & n59587;
  assign n62254 = n62264 & n62265;
  assign n62266 = ~n62272;
  assign n59821 = n62209 ^ n62210;
  assign n62164 = n62210 & n62212;
  assign n62215 = n62205 & n456;
  assign n62224 = ~n62230;
  assign n62228 = ~n62205;
  assign n62231 = n62235 & n62203;
  assign n62232 = n58347 & n62236;
  assign n60940 = ~n62237;
  assign n62233 = n58347 & n60780;
  assign n62219 = ~n62239;
  assign n62246 = ~n62254;
  assign n62227 = ~n62255;
  assign n62238 = n62266 & n62267;
  assign n62170 = ~n62164;
  assign n62178 = ~n62215;
  assign n62204 = n62224 & n62225;
  assign n62213 = n62228 & n18051;
  assign n62201 = ~n62231;
  assign n60972 = ~n62232;
  assign n62226 = ~n62233;
  assign n62223 = n62238 ^ n59504;
  assign n62216 = n62246 & n62247;
  assign n62240 = ~n62238;
  assign n62176 = n62204 ^ n62205;
  assign n62206 = ~n62213;
  assign n62207 = ~n62204;
  assign n62202 = n62216 ^ n62217;
  assign n58232 = n62222 ^ n62223;
  assign n62171 = n62226 & n62227;
  assign n62218 = ~n62216;
  assign n62234 = n62240 & n62241;
  assign n62165 = n456 ^ n62176;
  assign n62163 = n62202 ^ n62203;
  assign n62191 = n62206 & n62207;
  assign n62196 = n58232 & n59504;
  assign n62195 = n62171 & n62211;
  assign n62208 = ~n62171;
  assign n58237 = ~n58232;
  assign n62214 = n62218 & n62219;
  assign n62220 = ~n62234;
  assign n62147 = n62164 ^ n62165;
  assign n62169 = ~n62165;
  assign n62188 = n62163 & n471;
  assign n62177 = ~n62191;
  assign n62179 = ~n62163;
  assign n62193 = n58237 & n60748;
  assign n62186 = ~n62195;
  assign n62190 = ~n62196;
  assign n62192 = n62208 & n62181;
  assign n62200 = ~n62214;
  assign n62197 = n62220 & n62221;
  assign n62041 = n62147 & n58974;
  assign n62130 = n62147 & n58970;
  assign n62144 = ~n62147;
  assign n62123 = n62169 & n62170;
  assign n62162 = n62177 & n62178;
  assign n62174 = n62179 & n17983;
  assign n62143 = ~n62188;
  assign n62154 = ~n62192;
  assign n62189 = ~n62193;
  assign n62183 = n62197 ^ n59466;
  assign n62180 = n62200 & n62201;
  assign n62198 = ~n62197;
  assign n61030 = ~n62130;
  assign n62127 = n62144 & n58974;
  assign n62126 = ~n62123;
  assign n62146 = n62162 ^ n62163;
  assign n62166 = ~n62174;
  assign n62167 = ~n62162;
  assign n62172 = n62180 ^ n62181;
  assign n58173 = n62182 ^ n62183;
  assign n62133 = n62189 & n62190;
  assign n62187 = ~n62180;
  assign n62194 = n62198 & n62199;
  assign n62077 = ~n62127;
  assign n62124 = n471 ^ n62146;
  assign n62148 = n62166 & n62167;
  assign n62122 = n62171 ^ n62172;
  assign n62155 = n58173 & n60698;
  assign n62156 = n62133 & n62173;
  assign n62157 = n58173 & n60812;
  assign n62168 = ~n62133;
  assign n58271 = ~n58173;
  assign n62175 = n62186 & n62187;
  assign n62184 = ~n62194;
  assign n62101 = n62123 ^ n62124;
  assign n57840 = n62077 & n61030;
  assign n62072 = n62124 & n62126;
  assign n62131 = n62122 & n470;
  assign n62142 = ~n62148;
  assign n62145 = ~n62122;
  assign n62135 = ~n62155;
  assign n62137 = ~n62156;
  assign n60843 = ~n62157;
  assign n62150 = n58271 & n62161;
  assign n62151 = n58271 & n59466;
  assign n62149 = n62168 & n62108;
  assign n62153 = ~n62175;
  assign n62158 = n62184 & n62185;
  assign n62095 = n62101 & n58927;
  assign n62083 = n57840 & n61004;
  assign n57838 = ~n57840;
  assign n62096 = ~n62101;
  assign n62058 = ~n62072;
  assign n62085 = ~n62131;
  assign n62121 = n62142 & n62143;
  assign n62128 = n62145 & n17956;
  assign n62119 = ~n62149;
  assign n60808 = ~n62150;
  assign n62134 = ~n62151;
  assign n62132 = n62153 & n62154;
  assign n62139 = n62158 ^ n59424;
  assign n62159 = ~n62158;
  assign n62076 = ~n62083;
  assign n62046 = ~n62095;
  assign n62082 = n62096 & n58931;
  assign n62098 = n62121 ^ n62122;
  assign n62117 = ~n62128;
  assign n62116 = ~n62121;
  assign n62107 = n62132 ^ n62133;
  assign n62061 = n62134 & n62135;
  assign n58136 = n62138 ^ n62139;
  assign n62136 = ~n62132;
  assign n62152 = n62159 & n62160;
  assign n62049 = n62076 & n62077;
  assign n62056 = ~n62082;
  assign n62073 = n470 ^ n62098;
  assign n62060 = n62107 ^ n62108;
  assign n62102 = n62116 & n62117;
  assign n62110 = n58136 & n59455;
  assign n62111 = n58136 & n60778;
  assign n62109 = n62061 & n62125;
  assign n58150 = ~n58136;
  assign n62120 = ~n62061;
  assign n62129 = n62136 & n62137;
  assign n62140 = ~n62152;
  assign n62022 = n62049 ^ n62048;
  assign n62054 = n62056 & n62041;
  assign n61979 = n62072 ^ n62073;
  assign n62040 = n62046 & n62056;
  assign n62047 = ~n62049;
  assign n62057 = ~n62073;
  assign n62097 = n62060 & n469;
  assign n62084 = ~n62102;
  assign n62086 = ~n62060;
  assign n62088 = ~n62109;
  assign n62093 = ~n62110;
  assign n60734 = ~n62111;
  assign n62104 = n58150 & n62115;
  assign n62105 = n58150 & n60641;
  assign n62103 = n62120 & n62100;
  assign n62118 = ~n62129;
  assign n62112 = n62140 & n62141;
  assign n59414 = n487 ^ n62022;
  assign n62020 = ~n62022;
  assign n57756 = n62040 ^ n62041;
  assign n61891 = n62047 & n62048;
  assign n62026 = n61979 & n58893;
  assign n62044 = ~n61979;
  assign n62045 = ~n62054;
  assign n62000 = n62057 & n62058;
  assign n62059 = n62084 & n62085;
  assign n62081 = n62086 & n17901;
  assign n62043 = ~n62097;
  assign n62070 = ~n62103;
  assign n60776 = ~n62104;
  assign n62094 = ~n62105;
  assign n62090 = n62112 ^ n59386;
  assign n62099 = n62118 & n62119;
  assign n62113 = ~n62112;
  assign n61738 = ~n59414;
  assign n61772 = n62020 & n487;
  assign n61997 = n57756 & n58931;
  assign n61996 = n57756 & n58927;
  assign n57758 = ~n57756;
  assign n61984 = ~n62026;
  assign n62023 = n62044 & n58903;
  assign n62018 = n62045 & n62046;
  assign n62039 = n62059 ^ n62060;
  assign n62075 = ~n62081;
  assign n62074 = ~n62059;
  assign n58082 = n62089 ^ n62090;
  assign n62004 = n62093 & n62094;
  assign n62062 = n62099 ^ n62100;
  assign n62087 = ~n62099;
  assign n62106 = n62113 & n62114;
  assign n61981 = ~n61996;
  assign n60926 = ~n61997;
  assign n61980 = n62018 ^ n58893;
  assign n61995 = n57758 & n60899;
  assign n61998 = ~n62018;
  assign n61999 = ~n62023;
  assign n62001 = n469 ^ n62039;
  assign n62017 = n62061 ^ n62062;
  assign n62055 = n62074 & n62075;
  assign n62064 = n58082 & n60546;
  assign n62063 = n62004 & n62078;
  assign n62071 = n58082 & n62079;
  assign n62066 = ~n62004;
  assign n58191 = ~n58082;
  assign n62080 = n62087 & n62088;
  assign n62091 = ~n62106;
  assign n57692 = n61979 ^ n61980;
  assign n61982 = ~n61995;
  assign n61989 = n61998 & n61999;
  assign n61917 = n62000 ^ n62001;
  assign n62019 = ~n62001;
  assign n62027 = n62017 & n468;
  assign n62038 = ~n62017;
  assign n62042 = ~n62055;
  assign n62033 = ~n62063;
  assign n62030 = ~n62064;
  assign n62051 = n58191 & n59411;
  assign n62050 = n62066 & n62029;
  assign n60703 = ~n62071;
  assign n62053 = n58191 & n60661;
  assign n62069 = ~n62080;
  assign n62065 = n62091 & n62092;
  assign n61957 = n57692 & n60847;
  assign n57704 = ~n57692;
  assign n61961 = n61981 & n61982;
  assign n61967 = n61917 & n58878;
  assign n61983 = ~n61989;
  assign n61966 = ~n61917;
  assign n61953 = n62019 & n62000;
  assign n61970 = ~n62027;
  assign n62025 = n62038 & n17859;
  assign n62016 = n62042 & n62043;
  assign n62007 = ~n62050;
  assign n62031 = ~n62051;
  assign n60664 = ~n62053;
  assign n62035 = n62065 ^ n59347;
  assign n62028 = n62069 & n62070;
  assign n62067 = ~n62065;
  assign n61925 = n57704 & n58903;
  assign n61933 = n57704 & n58893;
  assign n61919 = ~n61957;
  assign n61934 = n61961 & n61962;
  assign n61955 = ~n61961;
  assign n61963 = n61966 & n58862;
  assign n61952 = ~n61967;
  assign n61935 = n61983 & n61984;
  assign n61960 = ~n61953;
  assign n61968 = n62016 ^ n62017;
  assign n62002 = ~n62016;
  assign n62003 = ~n62025;
  assign n62005 = n62028 ^ n62029;
  assign n61949 = n62030 & n62031;
  assign n58047 = n62034 ^ n62035;
  assign n62032 = ~n62028;
  assign n62052 = n62067 & n62068;
  assign n60874 = ~n61925;
  assign n61920 = ~n61933;
  assign n61901 = ~n61934;
  assign n61918 = n61935 ^ n58862;
  assign n61926 = n61955 & n61956;
  assign n61912 = ~n61963;
  assign n61951 = ~n61935;
  assign n61954 = n468 ^ n61968;
  assign n61990 = n62002 & n62003;
  assign n61937 = n62004 ^ n62005;
  assign n62012 = n58047 & n60401;
  assign n62011 = n58047 & n60628;
  assign n62010 = n61949 & n62021;
  assign n62008 = ~n61949;
  assign n58043 = ~n58047;
  assign n62024 = n62032 & n62033;
  assign n62036 = ~n62052;
  assign n57631 = n61917 ^ n61918;
  assign n61816 = n61919 & n61920;
  assign n61900 = n61901 & n61891;
  assign n61895 = ~n61926;
  assign n61932 = n61951 & n61952;
  assign n61826 = n61953 ^ n61954;
  assign n61868 = n61954 & n61960;
  assign n61972 = n61937 & n467;
  assign n61969 = ~n61990;
  assign n61971 = ~n61937;
  assign n61991 = n62008 & n61986;
  assign n61992 = n58043 & n62009;
  assign n61974 = ~n62010;
  assign n61993 = n58043 & n59347;
  assign n60626 = ~n62011;
  assign n61988 = ~n62012;
  assign n62006 = ~n62024;
  assign n62013 = n62036 & n62037;
  assign n61864 = n57631 & n58878;
  assign n61866 = n61816 & n61852;
  assign n61865 = n57631 & n58862;
  assign n61888 = ~n61816;
  assign n57640 = ~n57631;
  assign n61894 = ~n61900;
  assign n61890 = n61895 & n61901;
  assign n61902 = n61826 & n58829;
  assign n61922 = ~n61826;
  assign n61911 = ~n61932;
  assign n61936 = n61969 & n61970;
  assign n61964 = n61971 & n17816;
  assign n61924 = ~n61972;
  assign n61947 = ~n61991;
  assign n60586 = ~n61992;
  assign n61987 = ~n61993;
  assign n61985 = n62006 & n62007;
  assign n61976 = n62013 ^ n59301;
  assign n62014 = ~n62013;
  assign n60814 = ~n61864;
  assign n61846 = ~n61865;
  assign n61853 = ~n61866;
  assign n61857 = n57640 & n60782;
  assign n61856 = n61888 & n61889;
  assign n61855 = n61890 ^ n61891;
  assign n61851 = n61894 & n61895;
  assign n61842 = ~n61902;
  assign n61867 = n61911 & n61912;
  assign n61899 = n61922 & n58827;
  assign n61921 = n61936 ^ n61937;
  assign n61959 = ~n61964;
  assign n61958 = ~n61936;
  assign n57994 = n61975 ^ n61976;
  assign n61950 = n61985 ^ n61986;
  assign n61886 = n61987 & n61988;
  assign n61973 = ~n61985;
  assign n61994 = n62014 & n62015;
  assign n61817 = n61851 ^ n61852;
  assign n61825 = n61855 & n486;
  assign n61819 = ~n61856;
  assign n61845 = ~n61857;
  assign n61850 = ~n61855;
  assign n61854 = ~n61851;
  assign n61827 = n61867 ^ n58827;
  assign n61892 = ~n61867;
  assign n61893 = ~n61899;
  assign n61869 = n467 ^ n61921;
  assign n61882 = n61949 ^ n61950;
  assign n61927 = n61958 & n61959;
  assign n61940 = n57994 & n60384;
  assign n61941 = n57994 & n60506;
  assign n61942 = n61886 & n61906;
  assign n61938 = ~n61886;
  assign n58104 = ~n57994;
  assign n61965 = n61973 & n61974;
  assign n61977 = ~n61994;
  assign n61737 = n61816 ^ n61817;
  assign n61750 = ~n61825;
  assign n57560 = n61826 ^ n61827;
  assign n61743 = n61845 & n61846;
  assign n61820 = n61850 & n9791;
  assign n61844 = n61853 & n61854;
  assign n61752 = n61868 ^ n61869;
  assign n61858 = n61892 & n61893;
  assign n61807 = n61869 & n61868;
  assign n61904 = n61882 & n466;
  assign n61923 = ~n61927;
  assign n61903 = ~n61882;
  assign n61928 = n61938 & n61939;
  assign n61910 = ~n61940;
  assign n60542 = ~n61941;
  assign n61908 = ~n61942;
  assign n61930 = n58104 & n61948;
  assign n61931 = n58104 & n59301;
  assign n61946 = ~n61965;
  assign n61943 = n61977 & n61978;
  assign n61776 = n61737 & n9753;
  assign n61777 = ~n61737;
  assign n61815 = n57560 & n58829;
  assign n61793 = n61743 & n61779;
  assign n61809 = n57560 & n58827;
  assign n61792 = ~n61820;
  assign n57598 = ~n57560;
  assign n61810 = ~n61743;
  assign n61818 = ~n61844;
  assign n61828 = n61752 & n58783;
  assign n61841 = ~n61858;
  assign n61843 = ~n61752;
  assign n61897 = n61903 & n17747;
  assign n61849 = ~n61904;
  assign n61881 = n61923 & n61924;
  assign n61871 = ~n61928;
  assign n60505 = ~n61930;
  assign n61909 = ~n61931;
  assign n61916 = n61943 ^ n59240;
  assign n61905 = n61946 & n61947;
  assign n61944 = ~n61943;
  assign n61710 = ~n61776;
  assign n61748 = n61777 & n485;
  assign n61771 = n61792 & n61750;
  assign n61786 = n57598 & n60656;
  assign n61783 = ~n61793;
  assign n60692 = ~n61809;
  assign n61784 = n61810 & n61811;
  assign n61774 = ~n61815;
  assign n61785 = n61792 & n61772;
  assign n61778 = n61818 & n61819;
  assign n61813 = ~n61828;
  assign n61814 = n61841 & n61842;
  assign n61821 = n61843 & n58791;
  assign n61839 = n61881 ^ n61882;
  assign n61884 = ~n61897;
  assign n61883 = ~n61881;
  assign n61887 = n61905 ^ n61906;
  assign n61796 = n61909 & n61910;
  assign n57934 = n61915 ^ n61916;
  assign n61907 = ~n61905;
  assign n61929 = n61944 & n61945;
  assign n61670 = ~n61748;
  assign n61735 = n61771 ^ n61772;
  assign n61744 = n61778 ^ n61779;
  assign n61740 = ~n61784;
  assign n61749 = ~n61785;
  assign n61773 = ~n61786;
  assign n61782 = ~n61778;
  assign n61753 = n61814 ^ n58783;
  assign n61812 = ~n61814;
  assign n61755 = ~n61821;
  assign n61808 = n466 ^ n61839;
  assign n61859 = n61883 & n61884;
  assign n61806 = n61886 ^ n61887;
  assign n61876 = n61796 & n61831;
  assign n61875 = n57934 & n60196;
  assign n61874 = n57934 & n61896;
  assign n57960 = ~n57934;
  assign n61872 = ~n61796;
  assign n61898 = n61907 & n61908;
  assign n61913 = ~n61929;
  assign n59377 = n61735 ^ n59414;
  assign n61654 = n61735 & n61738;
  assign n61631 = n61743 ^ n61744;
  assign n61736 = n61749 & n61750;
  assign n57519 = n61752 ^ n61753;
  assign n61656 = n61773 & n61774;
  assign n61751 = n61782 & n61783;
  assign n61672 = n61807 ^ n61808;
  assign n61787 = n61812 & n61813;
  assign n61716 = n61808 & n61807;
  assign n61829 = n61806 & n17696;
  assign n61848 = ~n61859;
  assign n61847 = ~n61806;
  assign n61860 = n61872 & n61873;
  assign n60461 = ~n61874;
  assign n61833 = ~n61875;
  assign n61838 = ~n61876;
  assign n61863 = n57960 & n61885;
  assign n61861 = n57960 & n59286;
  assign n61870 = ~n61898;
  assign n61879 = n61913 & n61914;
  assign n60464 = ~n59377;
  assign n61692 = n61631 & n9721;
  assign n61693 = ~n61631;
  assign n61689 = n61736 ^ n61737;
  assign n61715 = n61656 & n61695;
  assign n61714 = n57519 & n60556;
  assign n61711 = ~n61736;
  assign n57538 = ~n57519;
  assign n61712 = ~n61656;
  assign n61739 = ~n61751;
  assign n61756 = n61672 & n58757;
  assign n61754 = ~n61787;
  assign n61775 = ~n61672;
  assign n61795 = ~n61829;
  assign n61822 = n61847 & n465;
  assign n61805 = n61848 & n61849;
  assign n61803 = ~n61860;
  assign n61832 = ~n61861;
  assign n60417 = ~n61863;
  assign n61830 = n61870 & n61871;
  assign n61840 = n61879 ^ n61880;
  assign n61877 = ~n61879;
  assign n61655 = n485 ^ n61689;
  assign n61628 = ~n61692;
  assign n61668 = n61693 & n484;
  assign n61700 = n61710 & n61711;
  assign n61709 = n61712 & n61713;
  assign n61702 = n57538 & n58783;
  assign n61687 = ~n61714;
  assign n61699 = ~n61715;
  assign n61701 = n57538 & n58791;
  assign n61694 = n61739 & n61740;
  assign n61734 = n61754 & n61755;
  assign n61732 = ~n61756;
  assign n61745 = n61775 & n58749;
  assign n61768 = n61805 ^ n61806;
  assign n61794 = ~n61805;
  assign n61770 = ~n61822;
  assign n61797 = n61830 ^ n61831;
  assign n61684 = n61832 & n61833;
  assign n60462 = n60461 & n60417;
  assign n57903 = n59244 ^ n61840;
  assign n61837 = ~n61830;
  assign n61834 = ~n61840;
  assign n61862 = n61877 & n61878;
  assign n59337 = n61654 ^ n61655;
  assign n61567 = n61655 & n61654;
  assign n61608 = ~n61668;
  assign n61657 = n61694 ^ n61695;
  assign n61669 = ~n61700;
  assign n61688 = ~n61701;
  assign n60613 = ~n61702;
  assign n61666 = ~n61709;
  assign n61673 = n61734 ^ n58749;
  assign n61698 = ~n61694;
  assign n61733 = ~n61734;
  assign n61675 = ~n61745;
  assign n61717 = n465 ^ n61768;
  assign n61788 = n61794 & n61795;
  assign n61731 = n61796 ^ n61797;
  assign n61798 = n57903 & n60382;
  assign n58034 = ~n57903;
  assign n61824 = n61834 & n59244;
  assign n61823 = n61837 & n61838;
  assign n61835 = ~n61862;
  assign n60433 = ~n59337;
  assign n61570 = n61656 ^ n61657;
  assign n61630 = n61669 & n61670;
  assign n57481 = n61672 ^ n61673;
  assign n61583 = n61687 & n61688;
  assign n61671 = n61698 & n61699;
  assign n61600 = n61716 ^ n61717;
  assign n61707 = n61732 & n61733;
  assign n61718 = ~n61717;
  assign n61757 = n61731 & n17666;
  assign n61769 = ~n61788;
  assign n61758 = ~n61731;
  assign n60338 = ~n61798;
  assign n61789 = n58034 & n61804;
  assign n61790 = n58034 & n60178;
  assign n61802 = ~n61823;
  assign n61760 = ~n61824;
  assign n61801 = n61835 & n61836;
  assign n61609 = n61570 & n9697;
  assign n61606 = n61630 ^ n61631;
  assign n61618 = ~n61570;
  assign n61653 = n57481 & n58757;
  assign n61635 = n61583 & n61611;
  assign n61634 = n57481 & n58749;
  assign n61632 = ~n61583;
  assign n57492 = ~n57481;
  assign n61629 = ~n61630;
  assign n61665 = ~n61671;
  assign n61676 = n61600 & n58700;
  assign n61674 = ~n61707;
  assign n61685 = ~n61600;
  assign n61651 = n61718 & n61716;
  assign n61728 = ~n61757;
  assign n61746 = n61758 & n464;
  assign n61730 = n61769 & n61770;
  assign n60380 = ~n61789;
  assign n61759 = ~n61790;
  assign n61765 = n61801 ^ n59175;
  assign n61780 = n61802 & n61803;
  assign n61799 = ~n61801;
  assign n61568 = n484 ^ n61606;
  assign n61571 = ~n61609;
  assign n61587 = n61618 & n483;
  assign n61627 = n61628 & n61629;
  assign n61626 = n61632 & n61633;
  assign n61619 = n57492 & n60452;
  assign n61604 = ~n61634;
  assign n61617 = ~n61635;
  assign n60552 = ~n61653;
  assign n61610 = n61665 & n61666;
  assign n61636 = n61674 & n61675;
  assign n61589 = ~n61676;
  assign n61667 = n61685 & n58719;
  assign n61658 = ~n61651;
  assign n61686 = n61730 ^ n61731;
  assign n61727 = ~n61730;
  assign n61691 = ~n61746;
  assign n61614 = n61759 & n61760;
  assign n57844 = n61764 ^ n61765;
  assign n61763 = n61780 & n61781;
  assign n61761 = ~n61780;
  assign n61791 = n61799 & n61800;
  assign n59317 = n61567 ^ n61568;
  assign n61483 = n61568 & n61567;
  assign n61525 = ~n61587;
  assign n61584 = n61610 ^ n61611;
  assign n61603 = ~n61619;
  assign n61580 = ~n61626;
  assign n61607 = ~n61627;
  assign n61601 = n61636 ^ n58700;
  assign n61616 = ~n61610;
  assign n61637 = ~n61667;
  assign n61638 = ~n61636;
  assign n61652 = n464 ^ n61686;
  assign n61703 = n61727 & n61728;
  assign n61720 = n57844 & n61741;
  assign n61721 = n57844 & n59187;
  assign n61722 = n61614 & n61742;
  assign n61726 = ~n61614;
  assign n57875 = ~n57844;
  assign n61747 = n61761 & n61762;
  assign n61729 = ~n61763;
  assign n61766 = ~n61791;
  assign n60267 = ~n59317;
  assign n61463 = n61583 ^ n61584;
  assign n57437 = n61600 ^ n61601;
  assign n61487 = n61603 & n61604;
  assign n61569 = n61607 & n61608;
  assign n61605 = n61616 & n61617;
  assign n61625 = n61637 & n61638;
  assign n61520 = n61651 ^ n61652;
  assign n61565 = n61652 & n61658;
  assign n61690 = ~n61703;
  assign n60252 = ~n61720;
  assign n61682 = ~n61721;
  assign n61664 = ~n61722;
  assign n61704 = n57875 & n60247;
  assign n61705 = n57875 & n60021;
  assign n61708 = n61726 & n61660;
  assign n61719 = n61729 & n61684;
  assign n61697 = ~n61747;
  assign n61723 = n61766 & n61767;
  assign n61526 = n61463 & n9663;
  assign n61535 = ~n61463;
  assign n61503 = n61569 ^ n61570;
  assign n61548 = n57437 & n60370;
  assign n61547 = n61487 & n61528;
  assign n57446 = ~n57437;
  assign n61545 = ~n61487;
  assign n61572 = ~n61569;
  assign n61579 = ~n61605;
  assign n61590 = n61520 & n58678;
  assign n61602 = ~n61520;
  assign n61588 = ~n61625;
  assign n61639 = n61690 & n61691;
  assign n60297 = ~n61704;
  assign n61681 = ~n61705;
  assign n61613 = ~n61708;
  assign n61696 = ~n61719;
  assign n61678 = n61723 ^ n59117;
  assign n61683 = n61697 & n61729;
  assign n61724 = ~n61723;
  assign n61484 = n483 ^ n61503;
  assign n61481 = ~n61526;
  assign n61504 = n61535 & n482;
  assign n61537 = n61545 & n61546;
  assign n61538 = n57446 & n58719;
  assign n61544 = n57446 & n58700;
  assign n61532 = ~n61547;
  assign n61522 = ~n61548;
  assign n61536 = n61571 & n61572;
  assign n61527 = n61579 & n61580;
  assign n61549 = n61588 & n61589;
  assign n61551 = ~n61590;
  assign n61585 = n61602 & n58665;
  assign n61593 = ~n61639;
  assign n57813 = n61677 ^ n61678;
  assign n61533 = n61681 & n61682;
  assign n61640 = n61683 ^ n61684;
  assign n61659 = n61696 & n61697;
  assign n61706 = n61724 & n61725;
  assign n59249 = n61483 ^ n61484;
  assign n61381 = n61484 & n61483;
  assign n61433 = ~n61504;
  assign n61488 = n61527 ^ n61528;
  assign n61524 = ~n61536;
  assign n61498 = ~n61537;
  assign n60456 = ~n61538;
  assign n61523 = ~n61544;
  assign n61521 = n61549 ^ n58665;
  assign n61531 = ~n61527;
  assign n61550 = ~n61549;
  assign n61519 = ~n61585;
  assign n61591 = n61639 ^ n61640;
  assign n61615 = n61659 ^ n61660;
  assign n61649 = n57813 & n59117;
  assign n61644 = n57813 & n61661;
  assign n61645 = n61533 & n61662;
  assign n61641 = n61640 & n479;
  assign n61650 = ~n61640;
  assign n61643 = ~n61533;
  assign n57969 = ~n57813;
  assign n61663 = ~n61659;
  assign n61679 = ~n61706;
  assign n60214 = ~n59249;
  assign n61403 = ~n61381;
  assign n61384 = n61487 ^ n61488;
  assign n57393 = n61520 ^ n61521;
  assign n61419 = n61522 & n61523;
  assign n61462 = n61524 & n61525;
  assign n61505 = n61531 & n61532;
  assign n61543 = n61550 & n61551;
  assign n61566 = n479 ^ n61591;
  assign n61511 = n61614 ^ n61615;
  assign n61554 = ~n61641;
  assign n61621 = n61643 & n61575;
  assign n60166 = ~n61644;
  assign n61577 = ~n61645;
  assign n61622 = n57969 & n60043;
  assign n61623 = n57969 & n60162;
  assign n61598 = ~n61649;
  assign n61620 = n61650 & n17570;
  assign n61642 = n61663 & n61664;
  assign n61646 = n61679 & n61680;
  assign n61441 = n61384 & n9619;
  assign n61438 = n61462 ^ n61463;
  assign n61455 = ~n61384;
  assign n61465 = n57393 & n58678;
  assign n61466 = n57393 & n58665;
  assign n61464 = n61419 & n61499;
  assign n61482 = ~n61462;
  assign n57407 = ~n57393;
  assign n61480 = ~n61419;
  assign n61497 = ~n61505;
  assign n61518 = ~n61543;
  assign n61439 = n61565 ^ n61566;
  assign n61564 = ~n61566;
  assign n61573 = n61511 & n478;
  assign n61582 = ~n61511;
  assign n61592 = ~n61620;
  assign n61530 = ~n61621;
  assign n61599 = ~n61622;
  assign n60220 = ~n61623;
  assign n61612 = ~n61642;
  assign n61595 = n61646 ^ n59090;
  assign n61647 = ~n61646;
  assign n61382 = n482 ^ n61438;
  assign n61401 = ~n61441;
  assign n61422 = n61455 & n481;
  assign n61453 = ~n61464;
  assign n60347 = ~n61465;
  assign n61456 = n57407 & n60290;
  assign n61437 = ~n61466;
  assign n61460 = n61480 & n61451;
  assign n61461 = n61481 & n61482;
  assign n61450 = n61497 & n61498;
  assign n61479 = n61518 & n61519;
  assign n61507 = n61439 & n58648;
  assign n61506 = ~n61439;
  assign n61424 = n61564 & n61565;
  assign n61478 = ~n61573;
  assign n61552 = n61582 & n17477;
  assign n61586 = n61592 & n61593;
  assign n57778 = n61594 ^ n61595;
  assign n61448 = n61598 & n61599;
  assign n61574 = n61612 & n61613;
  assign n61624 = n61647 & n61648;
  assign n59211 = n61381 ^ n61382;
  assign n61402 = ~n61382;
  assign n61363 = ~n61422;
  assign n61420 = n61450 ^ n61451;
  assign n61436 = ~n61456;
  assign n61407 = ~n61460;
  assign n61432 = ~n61461;
  assign n61452 = ~n61450;
  assign n61440 = n61479 ^ n58617;
  assign n61485 = ~n61479;
  assign n61500 = n61506 & n58617;
  assign n61486 = ~n61507;
  assign n61454 = ~n61424;
  assign n61508 = ~n61552;
  assign n61534 = n61574 ^ n61575;
  assign n61559 = n57778 & n59885;
  assign n61557 = n57778 & n61578;
  assign n61558 = n61448 & n61581;
  assign n61553 = ~n61586;
  assign n61556 = ~n61448;
  assign n57781 = ~n57778;
  assign n61576 = ~n61574;
  assign n61596 = ~n61624;
  assign n60136 = ~n59211;
  assign n61325 = n61402 & n61403;
  assign n61307 = n61419 ^ n61420;
  assign n61383 = n61432 & n61433;
  assign n61339 = n61436 & n61437;
  assign n57346 = n61439 ^ n61440;
  assign n61423 = n61452 & n61453;
  assign n61459 = n61485 & n61486;
  assign n61435 = ~n61500;
  assign n61427 = n61533 ^ n61534;
  assign n61510 = n61553 & n61554;
  assign n61539 = n61556 & n61491;
  assign n60128 = ~n61557;
  assign n61493 = ~n61558;
  assign n61540 = n57781 & n59114;
  assign n61541 = n57781 & n60079;
  assign n61512 = ~n61559;
  assign n61555 = n61576 & n61577;
  assign n61562 = n61596 & n61597;
  assign n61328 = ~n61325;
  assign n61364 = n61307 & n480;
  assign n61344 = n61383 ^ n61384;
  assign n61374 = ~n61307;
  assign n61386 = n57346 & n58617;
  assign n61387 = n61339 & n61371;
  assign n61385 = n57346 & n58648;
  assign n61404 = ~n61339;
  assign n61400 = ~n61383;
  assign n57375 = ~n57346;
  assign n61406 = ~n61423;
  assign n61434 = ~n61459;
  assign n61489 = n61427 & n477;
  assign n61467 = n61510 ^ n61511;
  assign n61496 = ~n61427;
  assign n61509 = ~n61510;
  assign n61443 = ~n61539;
  assign n61513 = ~n61540;
  assign n60082 = ~n61541;
  assign n61529 = ~n61555;
  assign n61514 = n61562 ^ n61563;
  assign n61560 = ~n61562;
  assign n61326 = n481 ^ n61344;
  assign n61287 = ~n61364;
  assign n61345 = n61374 & n9577;
  assign n60269 = ~n61385;
  assign n61346 = ~n61386;
  assign n61372 = ~n61387;
  assign n61377 = n57375 & n60184;
  assign n61375 = n61400 & n61401;
  assign n61376 = n61404 & n61405;
  assign n61370 = n61406 & n61407;
  assign n61388 = n61434 & n61435;
  assign n61425 = n478 ^ n61467;
  assign n61399 = ~n61489;
  assign n61468 = n61496 & n17431;
  assign n61501 = n61508 & n61509;
  assign n61368 = n61512 & n61513;
  assign n57718 = n59050 ^ n61514;
  assign n61490 = n61529 & n61530;
  assign n61515 = ~n61514;
  assign n61542 = n61560 & n61561;
  assign n59168 = n61325 ^ n61326;
  assign n61241 = n61326 & n61328;
  assign n61324 = ~n61345;
  assign n61340 = n61370 ^ n61371;
  assign n61362 = ~n61375;
  assign n61330 = ~n61376;
  assign n61347 = ~n61377;
  assign n61373 = ~n61370;
  assign n61350 = n61388 ^ n58579;
  assign n61361 = ~n61388;
  assign n61349 = n61424 ^ n61425;
  assign n61351 = n61425 & n61454;
  assign n61428 = ~n61468;
  assign n61449 = n61490 ^ n61491;
  assign n61472 = n61368 & n61410;
  assign n61471 = n57718 & n59866;
  assign n61476 = n57718 & n61495;
  assign n61469 = ~n61368;
  assign n57879 = ~n57718;
  assign n61477 = ~n61501;
  assign n61492 = ~n61490;
  assign n61502 = n61515 & n59070;
  assign n61516 = ~n61542;
  assign n60047 = ~n59168;
  assign n61243 = n61339 ^ n61340;
  assign n61260 = n61346 & n61347;
  assign n57309 = n61349 ^ n61350;
  assign n61306 = n61362 & n61363;
  assign n61348 = n61372 & n61373;
  assign n61390 = n61349 & n58588;
  assign n61389 = ~n61349;
  assign n61359 = n61448 ^ n61449;
  assign n61457 = n61469 & n61470;
  assign n61444 = ~n61471;
  assign n61417 = ~n61472;
  assign n61458 = n57879 & n59992;
  assign n60041 = ~n61476;
  assign n61426 = n61477 & n61478;
  assign n61475 = n61492 & n61493;
  assign n61445 = ~n61502;
  assign n61473 = n61516 & n61517;
  assign n61299 = n61243 & n9544;
  assign n61283 = n61306 ^ n61307;
  assign n61298 = ~n61243;
  assign n61308 = n61260 & n61341;
  assign n61310 = n57309 & n58579;
  assign n61309 = n57309 & n58588;
  assign n61327 = ~n61260;
  assign n57339 = ~n57309;
  assign n61323 = ~n61306;
  assign n61329 = ~n61348;
  assign n61378 = n61389 & n58579;
  assign n61318 = ~n61390;
  assign n61408 = n61359 & n476;
  assign n61391 = n61426 ^ n61427;
  assign n61418 = ~n61359;
  assign n61294 = n61444 & n61445;
  assign n61429 = ~n61426;
  assign n61366 = ~n61457;
  assign n59991 = ~n61458;
  assign n61431 = n61473 ^ n59014;
  assign n61442 = ~n61475;
  assign n61474 = n61473 & n61494;
  assign n61249 = n480 ^ n61283;
  assign n61274 = n61298 & n495;
  assign n61257 = ~n61299;
  assign n61291 = ~n61308;
  assign n61285 = ~n61309;
  assign n60182 = ~n61310;
  assign n61301 = n57339 & n60093;
  assign n61305 = n61323 & n61324;
  assign n61300 = n61327 & n61289;
  assign n61288 = n61329 & n61330;
  assign n61360 = ~n61378;
  assign n61352 = n477 ^ n61391;
  assign n61316 = ~n61408;
  assign n61392 = n61418 & n17352;
  assign n61411 = n61294 & n61336;
  assign n61421 = n61428 & n61429;
  assign n61414 = ~n61294;
  assign n57669 = n61430 ^ n61431;
  assign n61409 = n61442 & n61443;
  assign n61446 = ~n61474;
  assign n59147 = n61241 ^ n61249;
  assign n61240 = ~n61249;
  assign n61224 = ~n61274;
  assign n61261 = n61288 ^ n61289;
  assign n61259 = ~n61300;
  assign n61284 = ~n61301;
  assign n61286 = ~n61305;
  assign n61290 = ~n61288;
  assign n61238 = n61351 ^ n61352;
  assign n61343 = n61360 & n61361;
  assign n61272 = n61352 & n61351;
  assign n61354 = ~n61392;
  assign n61369 = n61409 ^ n61410;
  assign n61397 = n57669 & n59902;
  assign n61396 = n57669 & n59014;
  assign n61334 = ~n61411;
  assign n61394 = n61414 & n61415;
  assign n57678 = ~n57669;
  assign n61398 = ~n61421;
  assign n61416 = ~n61409;
  assign n61412 = n61446 & n61447;
  assign n59960 = ~n59147;
  assign n61183 = n61240 & n61241;
  assign n61186 = n61260 ^ n61261;
  assign n61206 = n61284 & n61285;
  assign n61242 = n61286 & n61287;
  assign n61282 = n61290 & n61291;
  assign n61311 = n61238 & n58531;
  assign n61320 = ~n61238;
  assign n61317 = ~n61343;
  assign n61276 = ~n61272;
  assign n61278 = n61368 ^ n61369;
  assign n61297 = ~n61394;
  assign n61380 = n57678 & n61395;
  assign n61355 = ~n61396;
  assign n59905 = ~n61397;
  assign n61358 = n61398 & n61399;
  assign n61379 = n57678 & n59783;
  assign n57799 = n61412 ^ n61413;
  assign n61393 = n61416 & n61417;
  assign n61234 = n61186 & n494;
  assign n61211 = n61242 ^ n61243;
  assign n61231 = ~n61186;
  assign n61245 = n61206 & n61268;
  assign n61244 = ~n61206;
  assign n61256 = ~n61242;
  assign n61258 = ~n61282;
  assign n61281 = ~n61311;
  assign n61303 = n61317 & n61318;
  assign n61302 = n61320 & n58566;
  assign n61337 = n61278 & n17233;
  assign n61338 = ~n61278;
  assign n61319 = n61358 ^ n61359;
  assign n61353 = ~n61358;
  assign n61356 = ~n61379;
  assign n59953 = ~n61380;
  assign n61367 = n57799 & n59709;
  assign n61365 = ~n61393;
  assign n59029 = ~n57799;
  assign n61184 = n495 ^ n61211;
  assign n61212 = n61231 & n9510;
  assign n61158 = ~n61234;
  assign n61239 = n61244 & n61233;
  assign n61230 = ~n61245;
  assign n61236 = n61256 & n61257;
  assign n61232 = n61258 & n61259;
  assign n61254 = ~n61302;
  assign n61270 = ~n61303;
  assign n61273 = n476 ^ n61319;
  assign n61280 = ~n61337;
  assign n61314 = n61338 & n475;
  assign n61342 = n61353 & n61354;
  assign n61225 = n61355 & n61356;
  assign n61335 = n61365 & n61366;
  assign n61331 = ~n61367;
  assign n61357 = n59029 & n59786;
  assign n59085 = n61183 ^ n61184;
  assign n61137 = n61184 & n61183;
  assign n61187 = ~n61212;
  assign n61207 = n61232 ^ n61233;
  assign n61223 = ~n61236;
  assign n61200 = ~n61239;
  assign n61229 = ~n61232;
  assign n61237 = n61270 ^ n58566;
  assign n61189 = n61272 ^ n61273;
  assign n61269 = n61281 & n61270;
  assign n61275 = ~n61273;
  assign n61252 = ~n61314;
  assign n61313 = n61225 & n61264;
  assign n61295 = n61335 ^ n61336;
  assign n61315 = ~n61342;
  assign n61321 = ~n61225;
  assign n61333 = ~n61335;
  assign n61332 = ~n61357;
  assign n59875 = ~n59085;
  assign n61128 = n61206 ^ n61207;
  assign n61185 = n61223 & n61224;
  assign n61220 = n61229 & n61230;
  assign n57286 = n61237 ^ n61238;
  assign n61246 = n61189 & n58492;
  assign n61253 = ~n61269;
  assign n61255 = ~n61189;
  assign n61221 = n61275 & n61276;
  assign n61217 = n61294 ^ n61295;
  assign n61267 = ~n61313;
  assign n61277 = n61315 & n61316;
  assign n61304 = n61321 & n61322;
  assign n61292 = n61331 & n61332;
  assign n61312 = n61333 & n61334;
  assign n61175 = n61128 & n493;
  assign n61171 = n61185 ^ n61186;
  assign n61174 = ~n61128;
  assign n61188 = ~n61185;
  assign n61210 = n57286 & n60051;
  assign n61199 = ~n61220;
  assign n57277 = ~n57286;
  assign n61192 = ~n61246;
  assign n61213 = n61253 & n61254;
  assign n61235 = n61255 & n58501;
  assign n61262 = n61217 & n17168;
  assign n61265 = ~n61217;
  assign n61247 = n61277 ^ n61278;
  assign n61178 = n61292 ^ n61293;
  assign n61279 = ~n61277;
  assign n61228 = ~n61304;
  assign n61296 = ~n61312;
  assign n61138 = n494 ^ n61171;
  assign n61172 = n61174 & n9459;
  assign n61119 = ~n61175;
  assign n61182 = n61187 & n61188;
  assign n61176 = n61199 & n61200;
  assign n61201 = n57277 & n58566;
  assign n61202 = n57277 & n58531;
  assign n61179 = ~n61210;
  assign n61190 = n61213 ^ n58492;
  assign n61215 = ~n61235;
  assign n61214 = ~n61213;
  assign n61222 = n475 ^ n61247;
  assign n61219 = ~n61262;
  assign n61248 = n61265 & n474;
  assign n61271 = n61279 & n61280;
  assign n61263 = n61296 & n61297;
  assign n59043 = n61137 ^ n61138;
  assign n61146 = ~n61138;
  assign n61145 = ~n61172;
  assign n61149 = n61176 ^ n61156;
  assign n61157 = ~n61182;
  assign n57231 = n61189 ^ n61190;
  assign n61142 = ~n61176;
  assign n61180 = ~n61201;
  assign n60088 = ~n61202;
  assign n61208 = n61214 & n61215;
  assign n61140 = n61221 ^ n61222;
  assign n61163 = n61222 & n61221;
  assign n61196 = ~n61248;
  assign n61226 = n61263 ^ n61264;
  assign n61251 = ~n61271;
  assign n61266 = ~n61263;
  assign n61095 = n61146 & n61137;
  assign n61127 = n61157 & n61158;
  assign n61159 = n57231 & n59922;
  assign n61148 = n61179 & n61180;
  assign n57265 = ~n57231;
  assign n61194 = n61140 & n58495;
  assign n61191 = ~n61208;
  assign n61193 = ~n61140;
  assign n61166 = ~n61163;
  assign n61168 = n61225 ^ n61226;
  assign n61216 = n61251 & n61252;
  assign n61250 = n61266 & n61267;
  assign n61117 = n61127 ^ n61128;
  assign n61080 = n61148 ^ n61149;
  assign n61144 = ~n61127;
  assign n61150 = n57265 & n58501;
  assign n61130 = ~n61159;
  assign n61154 = n57265 & n58492;
  assign n61153 = n61148 & n61173;
  assign n61155 = ~n61148;
  assign n61160 = n61191 & n61192;
  assign n61181 = n61193 & n58444;
  assign n61132 = ~n61194;
  assign n61203 = n61168 & n17141;
  assign n61198 = n61216 ^ n61217;
  assign n61205 = ~n61168;
  assign n61218 = ~n61216;
  assign n61227 = ~n61250;
  assign n61096 = n493 ^ n61117;
  assign n61120 = n61080 & n492;
  assign n61126 = n61144 & n61145;
  assign n61122 = ~n61080;
  assign n59997 = ~n61150;
  assign n61143 = ~n61153;
  assign n61129 = ~n61154;
  assign n61147 = n61155 & n61156;
  assign n61141 = n61160 ^ n58444;
  assign n61161 = ~n61160;
  assign n61162 = ~n61181;
  assign n61164 = n474 ^ n61198;
  assign n61170 = ~n61203;
  assign n61197 = n61205 & n473;
  assign n61209 = n61218 & n61219;
  assign n61204 = n61227 & n61228;
  assign n61057 = n61095 ^ n61096;
  assign n61097 = ~n61096;
  assign n61074 = ~n61120;
  assign n61103 = n61122 & n9421;
  assign n61118 = ~n61126;
  assign n61060 = n61129 & n61130;
  assign n57202 = n61140 ^ n61141;
  assign n61125 = n61142 & n61143;
  assign n61108 = ~n61147;
  assign n61151 = n61161 & n61162;
  assign n61081 = n61163 ^ n61164;
  assign n61165 = ~n61164;
  assign n61136 = ~n61197;
  assign n61177 = n472 ^ n61204;
  assign n61195 = ~n61209;
  assign n56789 = n57840 ^ n61057;
  assign n61058 = ~n61057;
  assign n61043 = n61097 & n61095;
  assign n61099 = ~n61103;
  assign n61079 = n61118 & n61119;
  assign n61106 = n57202 & n58495;
  assign n61116 = n57202 & n58444;
  assign n61105 = n61060 & n61123;
  assign n61104 = ~n61060;
  assign n61107 = ~n61125;
  assign n57197 = ~n57202;
  assign n61139 = n61081 & n58419;
  assign n61131 = ~n61151;
  assign n61133 = ~n61081;
  assign n61110 = n61165 & n61166;
  assign n61113 = n61177 ^ n61178;
  assign n61167 = n61195 & n61196;
  assign n61034 = n56789 & n58974;
  assign n56787 = ~n56789;
  assign n60970 = n61058 & n57838;
  assign n61052 = n61058 & n57840;
  assign n61051 = ~n61043;
  assign n61059 = n61079 ^ n61080;
  assign n61098 = ~n61079;
  assign n61102 = n61104 & n61084;
  assign n61093 = ~n61105;
  assign n61092 = ~n61106;
  assign n61100 = n57197 & n59827;
  assign n61083 = n61107 & n61108;
  assign n59909 = ~n61116;
  assign n61109 = n61131 & n61132;
  assign n61124 = n61133 & n58399;
  assign n61114 = ~n61139;
  assign n61121 = ~n61110;
  assign n61134 = n61167 ^ n61168;
  assign n61169 = ~n61167;
  assign n61029 = ~n61034;
  assign n58987 = ~n61052;
  assign n61044 = n492 ^ n61059;
  assign n61061 = n61083 ^ n61084;
  assign n61078 = n61098 & n61099;
  assign n61091 = ~n61100;
  assign n61094 = ~n61083;
  assign n61072 = ~n61102;
  assign n61082 = n61109 ^ n58399;
  assign n61115 = ~n61109;
  assign n61086 = ~n61124;
  assign n61111 = n473 ^ n61134;
  assign n61152 = n61169 & n61170;
  assign n61005 = n61029 & n61030;
  assign n61031 = n61043 ^ n61044;
  assign n60997 = n61044 & n61051;
  assign n61046 = n61060 ^ n61061;
  assign n61073 = ~n61078;
  assign n57187 = n61081 ^ n61082;
  assign n61014 = n61091 & n61092;
  assign n61076 = n61093 & n61094;
  assign n61041 = n61110 ^ n61111;
  assign n61101 = n61114 & n61115;
  assign n61089 = n61111 & n61121;
  assign n61135 = ~n61152;
  assign n60979 = n61005 ^ n61006;
  assign n61003 = ~n61005;
  assign n61028 = n61031 & n57756;
  assign n61012 = ~n61031;
  assign n60986 = ~n60997;
  assign n61035 = n61046 & n491;
  assign n61040 = ~n61046;
  assign n61045 = n61073 & n61074;
  assign n61064 = n57187 & n58419;
  assign n61065 = n57187 & n58399;
  assign n61063 = n61014 & n61075;
  assign n61071 = ~n61076;
  assign n61062 = ~n61014;
  assign n57136 = ~n57187;
  assign n61088 = n61041 & n58423;
  assign n61085 = ~n61101;
  assign n61087 = ~n61041;
  assign n61112 = n61135 & n61136;
  assign n58839 = n39 ^ n60979;
  assign n60741 = n60979 & n39;
  assign n60849 = n61003 & n61004;
  assign n61007 = n61012 & n57758;
  assign n60975 = ~n61028;
  assign n60989 = ~n61035;
  assign n61032 = n61040 & n9407;
  assign n61013 = n61045 ^ n61046;
  assign n61026 = ~n61045;
  assign n61056 = n61062 & n61048;
  assign n61050 = ~n61063;
  assign n59813 = ~n61064;
  assign n61036 = ~n61065;
  assign n61047 = n61071 & n61072;
  assign n61053 = n57136 & n59773;
  assign n61066 = n61085 & n61086;
  assign n61077 = n61087 & n58350;
  assign n61068 = ~n61088;
  assign n61090 = n61112 ^ n61113;
  assign n60668 = ~n58839;
  assign n60984 = ~n61007;
  assign n60998 = n491 ^ n61013;
  assign n61027 = ~n61032;
  assign n61015 = n61047 ^ n61048;
  assign n61049 = ~n61047;
  assign n61037 = ~n61053;
  assign n61025 = ~n61056;
  assign n61042 = n61066 ^ n58350;
  assign n61039 = ~n61077;
  assign n61067 = ~n61066;
  assign n60999 = n61089 ^ n61090;
  assign n60981 = n60984 & n60970;
  assign n60907 = n60997 ^ n60998;
  assign n60969 = n60975 & n60984;
  assign n60985 = ~n60998;
  assign n60961 = n61014 ^ n61015;
  assign n61008 = n61026 & n61027;
  assign n60976 = n61036 & n61037;
  assign n57105 = n61041 ^ n61042;
  assign n61033 = n61049 & n61050;
  assign n61054 = n61067 & n61068;
  assign n61070 = n60999 & n58324;
  assign n61069 = ~n60999;
  assign n56673 = n60969 ^ n60970;
  assign n60978 = n60907 & n57704;
  assign n60974 = ~n60981;
  assign n60957 = ~n60907;
  assign n60918 = n60985 & n60986;
  assign n60987 = n60961 & n490;
  assign n60988 = ~n61008;
  assign n60994 = ~n60961;
  assign n61020 = n57105 & n58350;
  assign n61019 = n60976 & n60991;
  assign n61018 = n57105 & n58423;
  assign n61016 = ~n60976;
  assign n61024 = ~n61033;
  assign n57111 = ~n57105;
  assign n61038 = ~n61054;
  assign n61055 = n61069 & n58321;
  assign n61023 = ~n61070;
  assign n60932 = n56673 & n58927;
  assign n60931 = n56673 & n57758;
  assign n56680 = ~n56673;
  assign n60956 = n60957 & n57692;
  assign n60949 = n60974 & n60975;
  assign n60921 = ~n60978;
  assign n60948 = ~n60987;
  assign n60960 = n60988 & n60989;
  assign n60982 = n60994 & n9340;
  assign n61009 = n61016 & n61017;
  assign n59746 = ~n61018;
  assign n60996 = ~n61019;
  assign n61002 = ~n61020;
  assign n60990 = n61024 & n61025;
  assign n61010 = n57111 & n59711;
  assign n61021 = n61038 & n61039;
  assign n60993 = ~n61055;
  assign n58935 = ~n60931;
  assign n60925 = ~n60932;
  assign n60908 = n60949 ^ n57692;
  assign n60933 = ~n60949;
  assign n60934 = ~n60956;
  assign n60946 = n60960 ^ n60961;
  assign n60958 = ~n60982;
  assign n60959 = ~n60960;
  assign n60977 = n60990 ^ n60991;
  assign n60995 = ~n60990;
  assign n60963 = ~n61009;
  assign n61001 = ~n61010;
  assign n61000 = n61021 ^ n58324;
  assign n61022 = ~n61021;
  assign n56610 = n60907 ^ n60908;
  assign n60903 = n60925 & n60926;
  assign n60930 = n60933 & n60934;
  assign n60919 = n490 ^ n60946;
  assign n60955 = n60958 & n60959;
  assign n60923 = n60976 ^ n60977;
  assign n60983 = n60995 & n60996;
  assign n57028 = n60999 ^ n61000;
  assign n60911 = n61001 & n61002;
  assign n61011 = n61022 & n61023;
  assign n60882 = n56610 & n58893;
  assign n60881 = n56610 & n57692;
  assign n60900 = n60903 & n60904;
  assign n56568 = ~n56610;
  assign n60862 = n60918 ^ n60919;
  assign n60898 = ~n60903;
  assign n60917 = ~n60919;
  assign n60920 = ~n60930;
  assign n60945 = n60923 & n9304;
  assign n60935 = ~n60923;
  assign n60947 = ~n60955;
  assign n60964 = n60911 & n60980;
  assign n60966 = n57028 & n58324;
  assign n60965 = n57028 & n59621;
  assign n60973 = ~n60911;
  assign n60962 = ~n60983;
  assign n57110 = ~n57028;
  assign n60992 = ~n61011;
  assign n58917 = ~n60881;
  assign n60873 = ~n60882;
  assign n60897 = n60898 & n60899;
  assign n60867 = ~n60900;
  assign n60883 = n60862 & n57640;
  assign n60895 = ~n60862;
  assign n60865 = n60917 & n60918;
  assign n60896 = n60920 & n60921;
  assign n60929 = n60935 & n489;
  assign n60909 = ~n60945;
  assign n60922 = n60947 & n60948;
  assign n60936 = n60962 & n60963;
  assign n60941 = ~n60964;
  assign n60943 = ~n60965;
  assign n59673 = ~n60966;
  assign n60953 = n57110 & n58324;
  assign n60952 = n60973 & n60937;
  assign n60967 = n60992 & n60993;
  assign n60783 = n60873 & n60874;
  assign n60872 = n60867 & n60849;
  assign n60871 = ~n60883;
  assign n60880 = n60895 & n57631;
  assign n60863 = n60896 ^ n57631;
  assign n60855 = ~n60897;
  assign n60870 = ~n60896;
  assign n60884 = n60922 ^ n60923;
  assign n60894 = ~n60929;
  assign n60910 = ~n60922;
  assign n60912 = n60936 ^ n60937;
  assign n60942 = ~n60936;
  assign n60916 = ~n60952;
  assign n60944 = ~n60953;
  assign n60951 = n60967 ^ n60968;
  assign n60971 = ~n60967;
  assign n60836 = n60783 & n60817;
  assign n56523 = n60862 ^ n60863;
  assign n60846 = ~n60783;
  assign n60848 = n60855 & n60867;
  assign n60861 = n60870 & n60871;
  assign n60854 = ~n60872;
  assign n60838 = ~n60880;
  assign n60866 = n489 ^ n60884;
  assign n60905 = n60909 & n60910;
  assign n60857 = n60911 ^ n60912;
  assign n60927 = n60941 & n60942;
  assign n60830 = n60943 & n60944;
  assign n60938 = n60951 & n58249;
  assign n60950 = ~n60951;
  assign n60954 = n60971 & n60972;
  assign n60821 = ~n60836;
  assign n60834 = n56523 & n57640;
  assign n60835 = n60846 & n60847;
  assign n60823 = n56523 & n58862;
  assign n60820 = n60848 ^ n60849;
  assign n56555 = ~n56523;
  assign n60816 = n60854 & n60855;
  assign n60837 = ~n60861;
  assign n60769 = n60865 ^ n60866;
  assign n60792 = n60866 & n60865;
  assign n60886 = n60857 & n488;
  assign n60893 = ~n60905;
  assign n60885 = ~n60857;
  assign n60915 = ~n60927;
  assign n60869 = ~n60938;
  assign n60928 = n60950 & n58347;
  assign n60939 = ~n60954;
  assign n60784 = n60816 ^ n60817;
  assign n60802 = n60820 & n38;
  assign n60813 = ~n60823;
  assign n60815 = ~n60820;
  assign n58883 = ~n60834;
  assign n60786 = ~n60835;
  assign n60822 = ~n60816;
  assign n60825 = n60769 & n57560;
  assign n60833 = n60837 & n60838;
  assign n60824 = ~n60769;
  assign n60879 = n60885 & n9262;
  assign n60832 = ~n60886;
  assign n60856 = n60893 & n60894;
  assign n60901 = n60915 & n60916;
  assign n59612 = ~n60928;
  assign n60924 = n60939 & n60940;
  assign n60694 = n60783 ^ n60784;
  assign n60743 = ~n60802;
  assign n60706 = n60813 & n60814;
  assign n60791 = n60815 & n12610;
  assign n60801 = n60821 & n60822;
  assign n60818 = n60824 & n57598;
  assign n60766 = ~n60825;
  assign n60799 = ~n60833;
  assign n60826 = n60856 ^ n60857;
  assign n60859 = ~n60856;
  assign n60858 = ~n60879;
  assign n60889 = n60901 & n60902;
  assign n60887 = ~n60901;
  assign n56994 = n59612 & n60869;
  assign n60914 = n60924 & n58237;
  assign n60913 = ~n60924;
  assign n60744 = n60694 & n12533;
  assign n60753 = ~n60694;
  assign n60771 = n60706 & n60750;
  assign n60770 = ~n60791;
  assign n60781 = ~n60706;
  assign n60768 = n60799 ^ n57598;
  assign n60785 = ~n60801;
  assign n60800 = ~n60818;
  assign n60793 = n488 ^ n60826;
  assign n60850 = n60858 & n60859;
  assign n60877 = n60887 & n60888;
  assign n60864 = ~n60889;
  assign n60890 = n56994 & n59587;
  assign n57059 = ~n56994;
  assign n60906 = n60913 & n58232;
  assign n60892 = ~n60914;
  assign n60704 = ~n60744;
  assign n60726 = n60753 & n37;
  assign n56440 = n60768 ^ n60769;
  assign n60755 = n60770 & n60741;
  assign n60752 = ~n60771;
  assign n60740 = n60770 & n60743;
  assign n60767 = n60781 & n60782;
  assign n60749 = n60785 & n60786;
  assign n60686 = n60792 ^ n60793;
  assign n60787 = n60799 & n60800;
  assign n60794 = ~n60793;
  assign n60831 = ~n60850;
  assign n60860 = n60864 & n60830;
  assign n60845 = ~n60877;
  assign n60868 = ~n60890;
  assign n60891 = n60892 & n60852;
  assign n60876 = ~n60906;
  assign n60666 = ~n60726;
  assign n58780 = n60740 ^ n60741;
  assign n56457 = ~n56440;
  assign n60707 = n60749 ^ n60750;
  assign n60742 = ~n60755;
  assign n60713 = ~n60767;
  assign n60756 = n60686 & n57519;
  assign n60751 = ~n60749;
  assign n60765 = ~n60787;
  assign n60764 = ~n60686;
  assign n60716 = n60794 & n60792;
  assign n60795 = n60831 & n60832;
  assign n60844 = ~n60860;
  assign n60829 = n60845 & n60864;
  assign n60804 = n60868 & n60869;
  assign n60875 = ~n60891;
  assign n60878 = n60876 & n60892;
  assign n60630 = n60706 ^ n60707;
  assign n60711 = n56457 & n57598;
  assign n60710 = n56457 & n58829;
  assign n58809 = ~n58780;
  assign n60693 = n60742 & n60743;
  assign n60727 = n60751 & n60752;
  assign n60724 = ~n60756;
  assign n60754 = n60764 & n57538;
  assign n60714 = n60765 & n60766;
  assign n60757 = n503 ^ n60795;
  assign n60760 = ~n60795;
  assign n60758 = n60829 ^ n60830;
  assign n60803 = n60844 & n60845;
  assign n60840 = n60804 & n60851;
  assign n60839 = ~n60804;
  assign n60841 = n60875 & n60876;
  assign n60853 = ~n60878;
  assign n60673 = n60630 & n12419;
  assign n60658 = n60693 ^ n60694;
  assign n60671 = ~n60630;
  assign n60691 = ~n60710;
  assign n58842 = ~n60711;
  assign n60705 = ~n60693;
  assign n60687 = n60714 ^ n57519;
  assign n60712 = ~n60727;
  assign n60723 = ~n60714;
  assign n60677 = ~n60754;
  assign n60725 = n60757 ^ n60758;
  assign n60779 = n60803 ^ n60804;
  assign n60796 = n60758 & n503;
  assign n60798 = ~n60758;
  assign n60805 = ~n60803;
  assign n60828 = n60839 & n60780;
  assign n60806 = ~n60840;
  assign n60811 = n60841 ^ n58173;
  assign n56968 = n60852 ^ n60853;
  assign n60842 = ~n60841;
  assign n60619 = n37 ^ n60658;
  assign n60657 = n60671 & n36;
  assign n60617 = ~n60673;
  assign n56365 = n60686 ^ n60687;
  assign n60631 = n60691 & n60692;
  assign n60690 = n60704 & n60705;
  assign n60672 = n60712 & n60713;
  assign n60708 = n60723 & n60724;
  assign n60610 = n60716 ^ n60725;
  assign n60715 = ~n60725;
  assign n60679 = n60779 ^ n60780;
  assign n60719 = ~n60796;
  assign n60788 = n60798 & n9219;
  assign n60797 = n60805 & n60806;
  assign n56917 = n60811 ^ n60812;
  assign n60819 = n56968 & n59504;
  assign n60773 = ~n60828;
  assign n60827 = n60842 & n60843;
  assign n56970 = ~n56968;
  assign n58761 = n60619 ^ n58780;
  assign n60536 = n60619 & n58780;
  assign n60588 = ~n60657;
  assign n60643 = n60631 & n60667;
  assign n60642 = n56365 & n60668;
  assign n56377 = ~n56365;
  assign n60655 = ~n60631;
  assign n60632 = n60672 ^ n60656;
  assign n60665 = ~n60690;
  assign n60689 = n60610 & n57492;
  assign n60620 = ~n60672;
  assign n60676 = ~n60708;
  assign n60688 = ~n60610;
  assign n60597 = n60715 & n60716;
  assign n60739 = n60679 & n502;
  assign n60728 = ~n60679;
  assign n60759 = ~n60788;
  assign n60774 = n56917 & n59466;
  assign n60772 = ~n60797;
  assign n56988 = ~n56917;
  assign n60809 = n56970 & n58237;
  assign n60789 = ~n60819;
  assign n60810 = n56970 & n58232;
  assign n60807 = ~n60827;
  assign n60483 = ~n58761;
  assign n60550 = n60631 ^ n60632;
  assign n58855 = ~n60642;
  assign n60633 = n56377 & n58791;
  assign n60621 = ~n60643;
  assign n60636 = n60655 & n60656;
  assign n60634 = n56377 & n58839;
  assign n60635 = n56377 & n57519;
  assign n60629 = n60665 & n60666;
  assign n60644 = n60676 & n60677;
  assign n60669 = n60688 & n57481;
  assign n60654 = ~n60689;
  assign n60717 = n60728 & n9190;
  assign n60652 = ~n60739;
  assign n60745 = n60759 & n60760;
  assign n60729 = n60772 & n60773;
  assign n60738 = ~n60774;
  assign n60763 = n56988 & n58173;
  assign n60761 = n56988 & n58271;
  assign n60777 = n60807 & n60808;
  assign n59565 = ~n60809;
  assign n60790 = ~n60810;
  assign n60595 = n60550 & n35;
  assign n60614 = n60620 & n60621;
  assign n60591 = n60629 ^ n60630;
  assign n60593 = ~n60550;
  assign n60612 = ~n60633;
  assign n58838 = ~n60634;
  assign n58808 = ~n60635;
  assign n60580 = ~n60636;
  assign n60611 = n60644 ^ n57481;
  assign n60618 = ~n60629;
  assign n60616 = ~n60669;
  assign n60653 = ~n60644;
  assign n60684 = ~n60717;
  assign n60696 = n60729 ^ n60730;
  assign n60718 = ~n60745;
  assign n60721 = ~n60729;
  assign n60737 = ~n60761;
  assign n59520 = ~n60763;
  assign n60731 = n60777 ^ n60778;
  assign n60695 = n60789 & n60790;
  assign n60775 = ~n60777;
  assign n60537 = n36 ^ n60591;
  assign n60592 = n60593 & n12343;
  assign n60503 = ~n60595;
  assign n56297 = n60610 ^ n60611;
  assign n60508 = n60612 & n60613;
  assign n60579 = ~n60614;
  assign n60596 = n60617 & n60618;
  assign n60637 = n60653 & n60654;
  assign n60600 = n60695 ^ n60696;
  assign n60678 = n60718 & n60719;
  assign n56874 = n58136 ^ n60731;
  assign n60601 = n60737 & n60738;
  assign n60732 = n60731 & n58136;
  assign n60746 = n60695 & n60730;
  assign n60736 = ~n60731;
  assign n60762 = n60775 & n60776;
  assign n60747 = ~n60695;
  assign n58722 = n60536 ^ n60537;
  assign n60471 = n60537 & n60536;
  assign n60555 = n60579 & n60580;
  assign n60561 = n56297 & n58749;
  assign n60575 = n56297 & n57492;
  assign n60574 = n60508 & n60590;
  assign n60553 = ~n60592;
  assign n56306 = ~n56297;
  assign n60576 = ~n60508;
  assign n60587 = ~n60596;
  assign n60615 = ~n60637;
  assign n60659 = n60600 & n9138;
  assign n60650 = n60678 ^ n60679;
  assign n60660 = ~n60600;
  assign n60685 = ~n60678;
  assign n60699 = n56874 & n59455;
  assign n60700 = n60601 & n60649;
  assign n56881 = ~n56874;
  assign n60697 = ~n60601;
  assign n60675 = ~n60732;
  assign n60720 = n60736 & n58150;
  assign n60722 = ~n60746;
  assign n60735 = n60747 & n60748;
  assign n60733 = ~n60762;
  assign n60366 = ~n58722;
  assign n60509 = n60555 ^ n60556;
  assign n60551 = ~n60561;
  assign n60547 = ~n60555;
  assign n60548 = ~n60574;
  assign n58756 = ~n60575;
  assign n60557 = n60576 & n60556;
  assign n60549 = n60587 & n60588;
  assign n60562 = n60615 & n60616;
  assign n60598 = n502 ^ n60650;
  assign n60607 = ~n60659;
  assign n60645 = n60660 & n501;
  assign n60670 = n60684 & n60685;
  assign n60682 = n60697 & n60698;
  assign n60674 = ~n60699;
  assign n60647 = ~n60700;
  assign n59475 = ~n60720;
  assign n60709 = n60721 & n60722;
  assign n60701 = n60733 & n60734;
  assign n60681 = ~n60735;
  assign n60475 = n60508 ^ n60509;
  assign n60517 = n60547 & n60548;
  assign n60510 = n60549 ^ n60550;
  assign n60420 = n60551 & n60552;
  assign n60512 = ~n60557;
  assign n60554 = ~n60549;
  assign n60543 = ~n60562;
  assign n60563 = n60597 ^ n60598;
  assign n60609 = ~n60598;
  assign n60578 = ~n60645;
  assign n60651 = ~n60670;
  assign n60525 = n60674 & n60675;
  assign n60605 = ~n60682;
  assign n60662 = n60701 ^ n58082;
  assign n60680 = ~n60709;
  assign n60702 = ~n60701;
  assign n60473 = n60475 & n34;
  assign n60469 = ~n60475;
  assign n60472 = n35 ^ n60510;
  assign n60499 = n60420 & n60516;
  assign n60511 = ~n60517;
  assign n60498 = ~n60420;
  assign n60535 = n60553 & n60554;
  assign n60518 = n60562 ^ n60563;
  assign n60565 = n60563 & n57437;
  assign n60564 = ~n60563;
  assign n60533 = n60609 & n60597;
  assign n60638 = n60525 & n60570;
  assign n60599 = n60651 & n60652;
  assign n60640 = ~n60525;
  assign n56823 = n60661 ^ n60662;
  assign n60648 = n60680 & n60681;
  assign n60683 = n60702 & n60703;
  assign n60434 = n60469 & n12231;
  assign n58709 = n60471 ^ n60472;
  assign n60391 = ~n60473;
  assign n60470 = ~n60472;
  assign n60497 = n60498 & n60452;
  assign n60454 = ~n60499;
  assign n60451 = n60511 & n60512;
  assign n56216 = n60518 ^ n57446;
  assign n60502 = ~n60535;
  assign n60519 = n60518 & n57437;
  assign n60558 = n60564 & n57446;
  assign n60544 = ~n60565;
  assign n60522 = ~n60533;
  assign n60566 = n60599 ^ n60600;
  assign n60572 = ~n60638;
  assign n60624 = n56823 & n58082;
  assign n60622 = n60640 & n60641;
  assign n60623 = n56823 & n58191;
  assign n60608 = ~n60599;
  assign n56904 = ~n56823;
  assign n60602 = n60648 ^ n60649;
  assign n60646 = ~n60648;
  assign n60663 = ~n60683;
  assign n60309 = ~n58709;
  assign n60413 = ~n60434;
  assign n60421 = n60451 ^ n60452;
  assign n60387 = n60470 & n60471;
  assign n60453 = ~n60451;
  assign n60426 = ~n60497;
  assign n60482 = n56216 & n58761;
  assign n60484 = n56216 & n58700;
  assign n60474 = n60502 & n60503;
  assign n56237 = ~n56216;
  assign n58727 = ~n60519;
  assign n60520 = n60543 & n60544;
  assign n60501 = ~n60558;
  assign n60534 = n501 ^ n60566;
  assign n60524 = n60601 ^ n60602;
  assign n60594 = n60607 & n60608;
  assign n60528 = ~n60622;
  assign n60582 = ~n60623;
  assign n59430 = ~n60624;
  assign n60606 = n56904 & n59411;
  assign n60639 = n60646 & n60647;
  assign n60627 = n60663 & n60664;
  assign n60300 = n60420 ^ n60421;
  assign n60392 = ~n60387;
  assign n60448 = n60453 & n60454;
  assign n60428 = n60474 ^ n60475;
  assign n58759 = ~n60482;
  assign n60476 = n56237 & n60483;
  assign n60455 = ~n60484;
  assign n60412 = ~n60474;
  assign n60500 = ~n60520;
  assign n60423 = n60533 ^ n60534;
  assign n60521 = ~n60534;
  assign n60567 = n60524 & n9098;
  assign n60577 = ~n60594;
  assign n60573 = ~n60524;
  assign n60581 = ~n60606;
  assign n60589 = n60627 ^ n60628;
  assign n60604 = ~n60639;
  assign n60625 = ~n60627;
  assign n60367 = n60300 & n33;
  assign n60389 = ~n60300;
  assign n60396 = n60412 & n60413;
  assign n60388 = n34 ^ n60428;
  assign n60425 = ~n60448;
  assign n60329 = n60455 & n60456;
  assign n58777 = ~n60476;
  assign n60467 = n60500 & n60501;
  assign n60485 = n60423 & n57407;
  assign n60496 = ~n60423;
  assign n60436 = n60521 & n60522;
  assign n60532 = ~n60567;
  assign n60559 = n60573 & n500;
  assign n60523 = n60577 & n60578;
  assign n60444 = n60581 & n60582;
  assign n56776 = n60589 ^ n58047;
  assign n60584 = n60589 & n58047;
  assign n60583 = ~n60589;
  assign n60569 = n60604 & n60605;
  assign n60603 = n60625 & n60626;
  assign n60304 = ~n60367;
  assign n58654 = n60387 ^ n60388;
  assign n60348 = n60389 & n12170;
  assign n60261 = n60388 & n60392;
  assign n60390 = ~n60396;
  assign n60369 = n60425 & n60426;
  assign n60422 = n60329 & n60432;
  assign n60427 = ~n60329;
  assign n60424 = n60467 ^ n57393;
  assign n60465 = ~n60485;
  assign n60466 = ~n60467;
  assign n60477 = n60496 & n57393;
  assign n60468 = ~n60436;
  assign n60486 = n60523 ^ n60524;
  assign n60495 = ~n60559;
  assign n60538 = n56776 & n59347;
  assign n60539 = n60444 & n60488;
  assign n60531 = ~n60523;
  assign n60545 = ~n60444;
  assign n56771 = ~n56776;
  assign n60526 = n60569 ^ n60570;
  assign n60568 = n60583 & n58043;
  assign n59382 = ~n60584;
  assign n60571 = ~n60569;
  assign n60585 = ~n60603;
  assign n60223 = ~n58654;
  assign n60327 = ~n60348;
  assign n60330 = n60369 ^ n60370;
  assign n60328 = n60390 & n60391;
  assign n60386 = ~n60369;
  assign n60385 = ~n60422;
  assign n56136 = n60423 ^ n60424;
  assign n60411 = n60427 & n60370;
  assign n60435 = n60465 & n60466;
  assign n60419 = ~n60477;
  assign n60437 = n500 ^ n60486;
  assign n60447 = n60525 ^ n60526;
  assign n60513 = n60531 & n60532;
  assign n60514 = ~n60538;
  assign n60490 = ~n60539;
  assign n60529 = n60545 & n60546;
  assign n60515 = ~n60568;
  assign n60560 = n60571 & n60572;
  assign n60540 = n60585 & n60586;
  assign n60299 = n33 ^ n60328;
  assign n60256 = n60329 ^ n60330;
  assign n60326 = ~n60328;
  assign n60350 = n60385 & n60386;
  assign n60371 = n56136 & n57407;
  assign n60372 = n56136 & n58665;
  assign n60368 = n56136 & n58722;
  assign n56160 = ~n56136;
  assign n60332 = ~n60411;
  assign n60418 = ~n60435;
  assign n60340 = n60436 ^ n60437;
  assign n60352 = n60437 & n60468;
  assign n60492 = n60447 & n9053;
  assign n60494 = ~n60513;
  assign n60493 = ~n60447;
  assign n60364 = n60514 & n60515;
  assign n60443 = ~n60529;
  assign n60507 = n60540 ^ n57994;
  assign n60527 = ~n60560;
  assign n60541 = ~n60540;
  assign n60262 = n60299 ^ n60300;
  assign n60288 = n60256 & n32;
  assign n60298 = ~n60256;
  assign n60311 = n60326 & n60327;
  assign n60331 = ~n60350;
  assign n60349 = n56160 & n60366;
  assign n58725 = ~n60368;
  assign n58689 = ~n60371;
  assign n60346 = ~n60372;
  assign n60410 = n60340 & n57375;
  assign n60373 = n60418 & n60419;
  assign n60397 = ~n60340;
  assign n60355 = ~n60352;
  assign n60479 = n60364 & n60491;
  assign n60450 = ~n60492;
  assign n60478 = n60493 & n499;
  assign n60446 = n60494 & n60495;
  assign n60481 = ~n60364;
  assign n56697 = n60506 ^ n60507;
  assign n60487 = n60527 & n60528;
  assign n60530 = n60541 & n60542;
  assign n58624 = n60261 ^ n60262;
  assign n60158 = n60262 & n60261;
  assign n60208 = ~n60288;
  assign n60270 = n60298 & n12118;
  assign n60303 = ~n60311;
  assign n60289 = n60331 & n60332;
  assign n60253 = n60346 & n60347;
  assign n58745 = ~n60349;
  assign n60341 = n60373 ^ n57346;
  assign n60374 = ~n60373;
  assign n60393 = n60397 & n57346;
  assign n60375 = ~n60410;
  assign n60398 = n60446 ^ n60447;
  assign n60409 = ~n60478;
  assign n60403 = ~n60479;
  assign n60457 = n60481 & n60401;
  assign n60459 = n56697 & n59377;
  assign n60449 = ~n60446;
  assign n60458 = n56697 & n59301;
  assign n60445 = n60487 ^ n60488;
  assign n56825 = ~n56697;
  assign n60489 = ~n60487;
  assign n60504 = ~n60530;
  assign n60137 = ~n58624;
  assign n60174 = ~n60158;
  assign n60258 = ~n60270;
  assign n60254 = n60289 ^ n60290;
  assign n60255 = n60303 & n60304;
  assign n60272 = ~n60289;
  assign n60305 = n60253 & n60325;
  assign n60307 = ~n60253;
  assign n56099 = n60340 ^ n60341;
  assign n60351 = n60374 & n60375;
  assign n60334 = ~n60393;
  assign n60353 = n499 ^ n60398;
  assign n60357 = n60444 ^ n60445;
  assign n60431 = n60449 & n60450;
  assign n60359 = ~n60457;
  assign n60440 = n56825 & n57994;
  assign n60430 = ~n60458;
  assign n59400 = ~n60459;
  assign n60438 = n56825 & n58104;
  assign n60439 = n56825 & n60464;
  assign n60480 = n60489 & n60490;
  assign n60463 = n60504 & n60505;
  assign n60168 = n60253 ^ n60254;
  assign n60206 = n60255 ^ n60256;
  assign n60257 = ~n60255;
  assign n60273 = ~n60305;
  assign n60293 = n60307 & n60290;
  assign n60292 = n56099 & n58617;
  assign n60291 = n56099 & n57375;
  assign n60287 = n56099 & n60309;
  assign n56080 = ~n56099;
  assign n60333 = ~n60351;
  assign n60259 = n60352 ^ n60353;
  assign n60354 = ~n60353;
  assign n60399 = n60357 & n9015;
  assign n60408 = ~n60431;
  assign n60407 = ~n60357;
  assign n60429 = ~n60438;
  assign n59380 = ~n60439;
  assign n59334 = ~n60440;
  assign n56607 = n60462 ^ n60463;
  assign n60442 = ~n60480;
  assign n60460 = ~n60463;
  assign n60159 = n32 ^ n60206;
  assign n60210 = n60168 & n47;
  assign n60209 = ~n60168;
  assign n60244 = n60257 & n60258;
  assign n60265 = n60272 & n60273;
  assign n58692 = ~n60287;
  assign n58659 = ~n60291;
  assign n60268 = ~n60292;
  assign n60246 = ~n60293;
  assign n60271 = n56080 & n58709;
  assign n60294 = n60333 & n60334;
  assign n60324 = n60259 & n57339;
  assign n60323 = ~n60259;
  assign n60276 = n60354 & n60355;
  assign n60363 = ~n60399;
  assign n60395 = n60407 & n498;
  assign n60356 = n60408 & n60409;
  assign n60284 = n60429 & n60430;
  assign n60415 = n56607 & n59240;
  assign n60414 = n56607 & n60433;
  assign n60400 = n60442 & n60443;
  assign n56638 = ~n56607;
  assign n60441 = n60460 & n60461;
  assign n58582 = n60158 ^ n60159;
  assign n60173 = ~n60159;
  assign n60193 = n60209 & n12057;
  assign n60126 = ~n60210;
  assign n60207 = ~n60244;
  assign n60245 = ~n60265;
  assign n60156 = n60268 & n60269;
  assign n58711 = ~n60271;
  assign n60260 = n60294 ^ n57309;
  assign n60301 = ~n60294;
  assign n60308 = n60323 & n57309;
  assign n60302 = ~n60324;
  assign n60321 = n60356 ^ n60357;
  assign n60320 = ~n60395;
  assign n60362 = ~n60356;
  assign n60376 = n60284 & n60316;
  assign n60365 = n60400 ^ n60401;
  assign n60383 = ~n60284;
  assign n59363 = ~n60414;
  assign n60377 = ~n60415;
  assign n60405 = n56638 & n59337;
  assign n60406 = n56638 & n57934;
  assign n60404 = n56638 & n57960;
  assign n60402 = ~n60400;
  assign n60416 = ~n60441;
  assign n60024 = ~n58582;
  assign n60073 = n60173 & n60174;
  assign n60171 = ~n60193;
  assign n60167 = n60207 & n60208;
  assign n60224 = n60156 & n60243;
  assign n60183 = n60245 & n60246;
  assign n60230 = ~n60156;
  assign n56041 = n60259 ^ n60260;
  assign n60274 = n60301 & n60302;
  assign n60264 = ~n60308;
  assign n60277 = n498 ^ n60321;
  assign n60344 = n60362 & n60363;
  assign n60283 = n60364 ^ n60365;
  assign n60318 = ~n60376;
  assign n60360 = n60383 & n60384;
  assign n60394 = n60402 & n60403;
  assign n60378 = ~n60404;
  assign n59336 = ~n60405;
  assign n59304 = ~n60406;
  assign n60381 = n60416 & n60417;
  assign n60086 = ~n60073;
  assign n60116 = n60167 ^ n60168;
  assign n60157 = n60183 ^ n60184;
  assign n60172 = ~n60167;
  assign n60211 = n56041 & n58654;
  assign n60212 = n56041 & n58588;
  assign n60203 = ~n60224;
  assign n60213 = n56041 & n57339;
  assign n60222 = n60230 & n60184;
  assign n60204 = ~n60183;
  assign n56058 = ~n56041;
  assign n60263 = ~n60274;
  assign n60169 = n60276 ^ n60277;
  assign n60286 = ~n60277;
  assign n60312 = n60283 & n497;
  assign n60319 = ~n60344;
  assign n60322 = ~n60283;
  assign n60281 = ~n60360;
  assign n60237 = n60377 & n60378;
  assign n60345 = n60381 ^ n60382;
  assign n60358 = ~n60394;
  assign n60379 = ~n60381;
  assign n60074 = n47 ^ n60116;
  assign n60076 = n60156 ^ n60157;
  assign n60139 = n60171 & n60172;
  assign n60180 = n60203 & n60204;
  assign n58657 = ~n60211;
  assign n60181 = ~n60212;
  assign n58623 = ~n60213;
  assign n60141 = ~n60222;
  assign n60205 = n56058 & n60223;
  assign n60231 = n60169 & n57277;
  assign n60221 = n60263 & n60264;
  assign n60241 = ~n60169;
  assign n60185 = n60286 & n60276;
  assign n60233 = ~n60312;
  assign n60282 = n60319 & n60320;
  assign n60306 = n60322 & n8981;
  assign n60336 = n60345 & n57903;
  assign n60339 = n60237 & n60196;
  assign n60315 = n60358 & n60359;
  assign n60342 = ~n60237;
  assign n60335 = ~n60345;
  assign n60361 = n60379 & n60380;
  assign n58541 = n60073 ^ n60074;
  assign n59994 = n60074 & n60086;
  assign n60091 = n60076 & n46;
  assign n60115 = ~n60076;
  assign n60125 = ~n60139;
  assign n60140 = ~n60180;
  assign n60052 = n60181 & n60182;
  assign n58676 = ~n60205;
  assign n60170 = n60221 ^ n57286;
  assign n60200 = ~n60221;
  assign n60144 = ~n60231;
  assign n60225 = n60241 & n57286;
  assign n60202 = ~n60185;
  assign n60242 = n60282 ^ n60283;
  assign n60278 = ~n60282;
  assign n60279 = ~n60306;
  assign n60285 = n60315 ^ n60316;
  assign n60314 = n60335 & n58034;
  assign n60229 = ~n60336;
  assign n60240 = ~n60339;
  assign n60313 = n60342 & n60343;
  assign n60317 = ~n60315;
  assign n60337 = ~n60361;
  assign n59919 = ~n58541;
  assign n59987 = ~n59994;
  assign n60030 = ~n60091;
  assign n60083 = n60115 & n12021;
  assign n60075 = n60125 & n60126;
  assign n60092 = n60140 & n60141;
  assign n60132 = n60052 & n60142;
  assign n56000 = n60169 ^ n60170;
  assign n60131 = ~n60052;
  assign n60199 = ~n60225;
  assign n60186 = n497 ^ n60242;
  assign n60266 = n60278 & n60279;
  assign n60188 = n60284 ^ n60285;
  assign n60190 = ~n60313;
  assign n59262 = ~n60314;
  assign n60310 = n60317 & n60318;
  assign n60295 = n60337 & n60338;
  assign n60033 = n60075 ^ n60076;
  assign n60072 = ~n60083;
  assign n60071 = ~n60075;
  assign n60053 = n60092 ^ n60093;
  assign n60129 = n60131 & n60093;
  assign n60118 = n56000 & n58566;
  assign n60112 = ~n60132;
  assign n60130 = n56000 & n57286;
  assign n60111 = ~n60092;
  assign n60117 = n56000 & n60137;
  assign n56005 = ~n56000;
  assign n60056 = n60185 ^ n60186;
  assign n60175 = n60199 & n60200;
  assign n60201 = ~n60186;
  assign n60234 = n60188 & n8944;
  assign n60232 = ~n60266;
  assign n60235 = ~n60188;
  assign n60248 = n60295 ^ n57844;
  assign n56731 = n60229 & n59262;
  assign n60280 = ~n60310;
  assign n60296 = ~n60295;
  assign n59995 = n46 ^ n60033;
  assign n59980 = n60052 ^ n60053;
  assign n60044 = n60071 & n60072;
  assign n60089 = n60111 & n60112;
  assign n58621 = ~n60117;
  assign n60090 = n56005 & n58624;
  assign n60087 = ~n60118;
  assign n60055 = ~n60129;
  assign n58590 = ~n60130;
  assign n60145 = n60056 & n57265;
  assign n60143 = ~n60175;
  assign n60155 = ~n60056;
  assign n60113 = n60201 & n60202;
  assign n60187 = n60232 & n60233;
  assign n60198 = ~n60234;
  assign n60226 = n60235 & n496;
  assign n56471 = n60247 ^ n60248;
  assign n60250 = n56731 & n59244;
  assign n60249 = n56731 & n60267;
  assign n56546 = ~n56731;
  assign n60236 = n60280 & n60281;
  assign n60275 = n60296 & n60297;
  assign n58507 = n59994 ^ n59995;
  assign n59986 = ~n59995;
  assign n60003 = n59980 & n45;
  assign n60029 = ~n60044;
  assign n60028 = ~n59980;
  assign n59963 = n60087 & n60088;
  assign n60054 = ~n60089;
  assign n58645 = ~n60090;
  assign n60094 = n60143 & n60144;
  assign n60068 = ~n60145;
  assign n60133 = n60155 & n57231;
  assign n60096 = ~n60113;
  assign n60154 = n60187 ^ n60188;
  assign n60153 = ~n60226;
  assign n60215 = n56471 & n57875;
  assign n60216 = n56471 & n57844;
  assign n60217 = n56471 & n59249;
  assign n60197 = ~n60187;
  assign n60195 = n60236 ^ n60237;
  assign n56674 = ~n56471;
  assign n59319 = ~n60249;
  assign n60228 = ~n60250;
  assign n60238 = n56546 & n59317;
  assign n60239 = ~n60236;
  assign n60251 = ~n60275;
  assign n59868 = ~n58507;
  assign n59895 = n59986 & n59987;
  assign n59943 = ~n60003;
  assign n59998 = n60028 & n11976;
  assign n59979 = n60029 & n60030;
  assign n60031 = n60054 & n60055;
  assign n60045 = n59963 & n60032;
  assign n60050 = ~n59963;
  assign n60057 = n60094 ^ n57231;
  assign n60109 = ~n60094;
  assign n60110 = ~n60133;
  assign n60114 = n496 ^ n60154;
  assign n60104 = n60195 ^ n60196;
  assign n60176 = n60197 & n60198;
  assign n60194 = n56674 & n60214;
  assign n60191 = n56674 & n59187;
  assign n59210 = ~n60215;
  assign n60161 = ~n60216;
  assign n59252 = ~n60217;
  assign n60148 = n60228 & n60229;
  assign n59294 = ~n60238;
  assign n60227 = n60239 & n60240;
  assign n60218 = n60251 & n60252;
  assign n59900 = ~n59895;
  assign n59916 = n59979 ^ n59980;
  assign n59984 = ~n59998;
  assign n59985 = ~n59979;
  assign n59964 = n60031 ^ n60032;
  assign n60026 = ~n60045;
  assign n60034 = n60050 & n60051;
  assign n60025 = ~n60031;
  assign n55967 = n60056 ^ n60057;
  assign n60084 = n60109 & n60110;
  assign n59977 = n60113 ^ n60114;
  assign n60095 = ~n60114;
  assign n60146 = n60104 & n8895;
  assign n60152 = ~n60176;
  assign n60151 = ~n60104;
  assign n60160 = ~n60191;
  assign n60179 = n60148 & n60098;
  assign n59275 = ~n60194;
  assign n60177 = ~n60148;
  assign n60163 = n60218 ^ n57813;
  assign n60189 = ~n60227;
  assign n60219 = ~n60218;
  assign n59896 = n45 ^ n59916;
  assign n59878 = n59963 ^ n59964;
  assign n59962 = n59984 & n59985;
  assign n60000 = n60025 & n60026;
  assign n59976 = ~n60034;
  assign n60006 = n55967 & n57231;
  assign n60004 = n55967 & n58582;
  assign n60005 = n55967 & n58492;
  assign n55947 = ~n55967;
  assign n60070 = n59977 & n57197;
  assign n60067 = ~n60084;
  assign n60066 = ~n59977;
  assign n60010 = n60095 & n60096;
  assign n60108 = ~n60146;
  assign n60134 = n60151 & n511;
  assign n60103 = n60152 & n60153;
  assign n60061 = n60160 & n60161;
  assign n56400 = n60162 ^ n60163;
  assign n60164 = n60177 & n60178;
  assign n60149 = ~n60179;
  assign n60147 = n60189 & n60190;
  assign n60192 = n60219 & n60220;
  assign n58461 = n59895 ^ n59896;
  assign n59795 = n59896 & n59900;
  assign n59917 = n59878 & n11934;
  assign n59918 = ~n59878;
  assign n59942 = ~n59962;
  assign n59975 = ~n60000;
  assign n58585 = ~n60004;
  assign n59996 = ~n60005;
  assign n58546 = ~n60006;
  assign n59999 = n55947 & n60024;
  assign n60049 = n60066 & n57202;
  assign n60007 = n60067 & n60068;
  assign n60009 = ~n60070;
  assign n60069 = n60103 ^ n60104;
  assign n60107 = ~n60103;
  assign n60063 = ~n60134;
  assign n60121 = n60061 & n60135;
  assign n60120 = n56400 & n60136;
  assign n60122 = n56400 & n57969;
  assign n60123 = n56400 & n57813;
  assign n60097 = n60147 ^ n60148;
  assign n56415 = ~n56400;
  assign n60119 = ~n60061;
  assign n60106 = ~n60164;
  assign n60150 = ~n60147;
  assign n60165 = ~n60192;
  assign n59756 = ~n58461;
  assign n59824 = ~n59795;
  assign n59897 = ~n59917;
  assign n59910 = n59918 & n44;
  assign n59877 = n59942 & n59943;
  assign n59921 = n59975 & n59976;
  assign n59893 = n59996 & n59997;
  assign n58605 = ~n59999;
  assign n59978 = n60007 ^ n57202;
  assign n60008 = ~n60007;
  assign n59982 = ~n60049;
  assign n60011 = n511 ^ n60069;
  assign n60013 = n60097 ^ n60098;
  assign n60085 = n60107 & n60108;
  assign n60099 = n60119 & n60021;
  assign n59214 = ~n60120;
  assign n60065 = ~n60121;
  assign n59179 = ~n60122;
  assign n60100 = n56415 & n59117;
  assign n60101 = n56415 & n59211;
  assign n60077 = ~n60123;
  assign n60138 = n60149 & n60150;
  assign n60124 = n60165 & n60166;
  assign n59859 = n59877 ^ n59878;
  assign n59898 = ~n59877;
  assign n59836 = ~n59910;
  assign n59894 = n59921 ^ n59922;
  assign n59914 = ~n59921;
  assign n59945 = n59893 & n59961;
  assign n59954 = ~n59893;
  assign n55924 = n59977 ^ n59978;
  assign n60002 = n60008 & n60009;
  assign n59888 = n60010 ^ n60011;
  assign n60027 = ~n60011;
  assign n60058 = n60013 & n8851;
  assign n60059 = ~n60013;
  assign n60062 = ~n60085;
  assign n60023 = ~n60099;
  assign n60078 = ~n60100;
  assign n59235 = ~n60101;
  assign n60080 = n60124 ^ n57778;
  assign n60105 = ~n60138;
  assign n60127 = ~n60124;
  assign n59796 = n44 ^ n59859;
  assign n59798 = n59893 ^ n59894;
  assign n59869 = n59897 & n59898;
  assign n59920 = n55924 & n58541;
  assign n59913 = ~n59945;
  assign n59924 = n55924 & n58495;
  assign n59923 = n59954 & n59922;
  assign n59925 = n55924 & n57197;
  assign n55929 = ~n55924;
  assign n59965 = n59888 & n57187;
  assign n59983 = ~n59888;
  assign n59981 = ~n60002;
  assign n59926 = n60027 & n60010;
  assign n60015 = ~n60058;
  assign n60046 = n60059 & n510;
  assign n60012 = n60062 & n60063;
  assign n59934 = n60077 & n60078;
  assign n56323 = n60079 ^ n60080;
  assign n60060 = n60105 & n60106;
  assign n60102 = n60127 & n60128;
  assign n58449 = n59795 ^ n59796;
  assign n59719 = n59796 & n59824;
  assign n59855 = n59798 & n43;
  assign n59835 = ~n59869;
  assign n59837 = ~n59798;
  assign n59901 = n59913 & n59914;
  assign n59915 = n55929 & n59919;
  assign n58539 = ~n59920;
  assign n59874 = ~n59923;
  assign n59908 = ~n59924;
  assign n58512 = ~n59925;
  assign n59892 = ~n59965;
  assign n59944 = n59981 & n59982;
  assign n59956 = n59983 & n57136;
  assign n59955 = ~n59926;
  assign n59970 = n60012 ^ n60013;
  assign n60014 = ~n60012;
  assign n59972 = ~n60046;
  assign n60035 = n56323 & n60047;
  assign n60037 = n59934 & n59969;
  assign n60036 = n56323 & n57781;
  assign n60038 = n56323 & n57778;
  assign n60020 = n60060 ^ n60061;
  assign n60042 = ~n59934;
  assign n56538 = ~n56323;
  assign n60064 = ~n60060;
  assign n60081 = ~n60102;
  assign n59683 = ~n58449;
  assign n59797 = n59835 & n59836;
  assign n59825 = n59837 & n11895;
  assign n59779 = ~n59855;
  assign n59873 = ~n59901;
  assign n59788 = n59908 & n59909;
  assign n58561 = ~n59915;
  assign n59889 = n59944 ^ n57187;
  assign n59940 = ~n59956;
  assign n59941 = ~n59944;
  assign n59927 = n510 ^ n59970;
  assign n60001 = n60014 & n60015;
  assign n59929 = n60020 ^ n60021;
  assign n59167 = ~n60035;
  assign n59988 = ~n60036;
  assign n59974 = ~n60037;
  assign n59135 = ~n60038;
  assign n60016 = n60042 & n60043;
  assign n60018 = n56538 & n59168;
  assign n60017 = n56538 & n59114;
  assign n60048 = n60064 & n60065;
  assign n60039 = n60081 & n60082;
  assign n59755 = n59797 ^ n59798;
  assign n59815 = ~n59825;
  assign n59814 = ~n59797;
  assign n59826 = n59873 & n59874;
  assign n59861 = n59788 & n59876;
  assign n59860 = ~n59788;
  assign n55879 = n59888 ^ n59889;
  assign n59799 = n59926 ^ n59927;
  assign n59911 = n59940 & n59941;
  assign n59845 = n59927 & n59955;
  assign n59967 = n59929 & n509;
  assign n59971 = ~n60001;
  assign n59966 = ~n59929;
  assign n59937 = ~n60016;
  assign n59989 = ~n60017;
  assign n59192 = ~n60018;
  assign n59993 = n60039 ^ n57718;
  assign n60022 = ~n60048;
  assign n60040 = ~n60039;
  assign n59720 = n43 ^ n59755;
  assign n59787 = n59814 & n59815;
  assign n59789 = n59826 ^ n59827;
  assign n59828 = ~n59826;
  assign n59838 = n59860 & n59827;
  assign n59829 = ~n59861;
  assign n59858 = n55879 & n59868;
  assign n55870 = ~n55879;
  assign n59879 = n59799 & n57111;
  assign n59891 = ~n59911;
  assign n59890 = ~n59799;
  assign n59957 = n59966 & n8797;
  assign n59881 = ~n59967;
  assign n59928 = n59971 & n59972;
  assign n59853 = n59988 & n59989;
  assign n56262 = n59992 ^ n59993;
  assign n59968 = n60022 & n60023;
  assign n60019 = n60040 & n60041;
  assign n58414 = n59719 ^ n59720;
  assign n59721 = ~n59720;
  assign n59778 = ~n59787;
  assign n59723 = n59788 ^ n59789;
  assign n59818 = n59828 & n59829;
  assign n59834 = n55870 & n58507;
  assign n59793 = ~n59838;
  assign n59830 = n55870 & n57136;
  assign n58527 = ~n59858;
  assign n59831 = n55870 & n58399;
  assign n59850 = ~n59879;
  assign n59870 = n59890 & n57105;
  assign n59856 = n59891 & n59892;
  assign n59899 = n59928 ^ n59929;
  assign n59938 = ~n59957;
  assign n59946 = n59853 & n59958;
  assign n59949 = n56262 & n57718;
  assign n59947 = n56262 & n59960;
  assign n59948 = n56262 & n57879;
  assign n59939 = ~n59928;
  assign n59935 = n59968 ^ n59969;
  assign n59950 = ~n59853;
  assign n56466 = ~n56262;
  assign n59973 = ~n59968;
  assign n59990 = ~n60019;
  assign n59640 = ~n58414;
  assign n59665 = n59721 & n59719;
  assign n59722 = n59778 & n59779;
  assign n59748 = n59723 & n42;
  assign n59753 = ~n59723;
  assign n59792 = ~n59818;
  assign n58469 = ~n59830;
  assign n59812 = ~n59831;
  assign n58506 = ~n59834;
  assign n59800 = n59856 ^ n57105;
  assign n59849 = ~n59856;
  assign n59802 = ~n59870;
  assign n59846 = n509 ^ n59899;
  assign n59840 = n59934 ^ n59935;
  assign n59912 = n59938 & n59939;
  assign n59887 = ~n59946;
  assign n59126 = ~n59947;
  assign n59906 = ~n59948;
  assign n59094 = ~n59949;
  assign n59932 = n56466 & n59147;
  assign n59930 = n59950 & n59885;
  assign n59931 = n56466 & n59070;
  assign n59959 = n59973 & n59974;
  assign n59951 = n59990 & n59991;
  assign n59674 = ~n59665;
  assign n59682 = n59722 ^ n59723;
  assign n59681 = ~n59748;
  assign n59717 = ~n59722;
  assign n59744 = n59753 & n11867;
  assign n59751 = n59792 & n59793;
  assign n55818 = n59799 ^ n59800;
  assign n59712 = n59812 & n59813;
  assign n59823 = n59845 ^ n59846;
  assign n59833 = n59849 & n59850;
  assign n59857 = ~n59846;
  assign n59882 = n59840 & n8745;
  assign n59880 = ~n59912;
  assign n59883 = ~n59840;
  assign n59852 = ~n59930;
  assign n59907 = ~n59931;
  assign n59149 = ~n59932;
  assign n59903 = n59951 ^ n57669;
  assign n59936 = ~n59959;
  assign n59952 = ~n59951;
  assign n59666 = n42 ^ n59682;
  assign n59716 = ~n59744;
  assign n59713 = n59751 ^ n59752;
  assign n59741 = ~n59751;
  assign n59757 = n55818 & n58461;
  assign n59759 = n55818 & n58350;
  assign n59760 = n59712 & n59752;
  assign n59758 = n55818 & n57111;
  assign n59772 = ~n59712;
  assign n55850 = ~n55818;
  assign n59810 = n59823 & n57028;
  assign n59811 = ~n59823;
  assign n59801 = ~n59833;
  assign n59761 = n59857 & n59845;
  assign n59839 = n59880 & n59881;
  assign n59847 = ~n59882;
  assign n59871 = n59883 & n508;
  assign n56207 = n59902 ^ n59903;
  assign n59770 = n59906 & n59907;
  assign n59884 = n59936 & n59937;
  assign n59933 = n59952 & n59953;
  assign n58353 = n59665 ^ n59666;
  assign n59591 = n59666 & n59674;
  assign n59647 = n59712 ^ n59713;
  assign n59704 = n59716 & n59717;
  assign n59747 = n55850 & n59756;
  assign n58464 = ~n59757;
  assign n58434 = ~n59758;
  assign n59745 = ~n59759;
  assign n59740 = ~n59760;
  assign n59749 = n59772 & n59773;
  assign n59726 = n59801 & n59802;
  assign n59775 = ~n59810;
  assign n59790 = n59811 & n57110;
  assign n59781 = ~n59761;
  assign n59809 = n59839 ^ n59840;
  assign n59863 = n59770 & n59806;
  assign n59817 = ~n59871;
  assign n59867 = n56207 & n59014;
  assign n59848 = ~n59839;
  assign n59862 = n56207 & n59875;
  assign n59854 = n59884 ^ n59885;
  assign n56212 = ~n56207;
  assign n59865 = ~n59770;
  assign n59886 = ~n59884;
  assign n59904 = ~n59933;
  assign n59577 = ~n58353;
  assign n59599 = ~n59591;
  assign n59675 = n59647 & n11822;
  assign n59680 = ~n59704;
  assign n59679 = ~n59647;
  assign n59724 = n59740 & n59741;
  assign n59669 = n59745 & n59746;
  assign n58486 = ~n59747;
  assign n59706 = ~n59749;
  assign n59774 = ~n59726;
  assign n59735 = ~n59790;
  assign n59762 = n508 ^ n59809;
  assign n59832 = n59847 & n59848;
  assign n59764 = n59853 ^ n59854;
  assign n59104 = ~n59862;
  assign n59842 = n56212 & n57678;
  assign n59844 = n56212 & n57669;
  assign n59808 = ~n59863;
  assign n59841 = n59865 & n59866;
  assign n59820 = ~n59867;
  assign n59843 = n56212 & n59085;
  assign n59872 = n59886 & n59887;
  assign n59864 = n59904 & n59905;
  assign n59648 = ~n59675;
  assign n59667 = n59679 & n41;
  assign n59646 = n59680 & n59681;
  assign n59707 = n59669 & n59642;
  assign n59705 = ~n59724;
  assign n59710 = ~n59669;
  assign n59703 = n59761 ^ n59762;
  assign n59754 = n59774 & n59775;
  assign n59725 = n59735 & n59775;
  assign n59780 = ~n59762;
  assign n59804 = n59764 & n507;
  assign n59816 = ~n59832;
  assign n59803 = ~n59764;
  assign n59777 = ~n59841;
  assign n59054 = ~n59842;
  assign n59082 = ~n59843;
  assign n59819 = ~n59844;
  assign n59822 = n59864 ^ n57799;
  assign n59851 = ~n59872;
  assign n59618 = n59646 ^ n59647;
  assign n59625 = ~n59667;
  assign n59649 = ~n59646;
  assign n59668 = n59705 & n59706;
  assign n59670 = ~n59707;
  assign n59684 = n59710 & n59711;
  assign n55810 = n59725 ^ n59726;
  assign n59728 = n59703 & n56994;
  assign n59727 = ~n59703;
  assign n59734 = ~n59754;
  assign n59697 = n59780 & n59781;
  assign n59791 = n59803 & n8665;
  assign n59737 = ~n59804;
  assign n59763 = n59816 & n59817;
  assign n59693 = n59819 & n59820;
  assign n56353 = n59821 ^ n59822;
  assign n59805 = n59851 & n59852;
  assign n59592 = n41 ^ n59618;
  assign n59645 = n59648 & n59649;
  assign n59641 = n59668 ^ n59669;
  assign n59644 = ~n59684;
  assign n59671 = ~n59668;
  assign n59701 = n55810 & n58449;
  assign n59686 = n55810 & n57028;
  assign n59685 = n55810 & n58321;
  assign n55754 = ~n55810;
  assign n59718 = n59727 & n57059;
  assign n59687 = ~n59728;
  assign n59702 = n59734 & n59735;
  assign n59690 = ~n59697;
  assign n59729 = n59763 ^ n59764;
  assign n59766 = ~n59791;
  assign n59785 = n56353 & n57799;
  assign n59784 = n59693 & n59733;
  assign n59765 = ~n59763;
  assign n59771 = n59805 ^ n59806;
  assign n59032 = ~n56353;
  assign n59782 = ~n59693;
  assign n59807 = ~n59805;
  assign n58314 = n59591 ^ n59592;
  assign n59547 = n59592 & n59599;
  assign n59594 = n59641 ^ n59642;
  assign n59624 = ~n59645;
  assign n59652 = n59670 & n59671;
  assign n59678 = n55754 & n59683;
  assign n59672 = ~n59685;
  assign n58395 = ~n59686;
  assign n58451 = ~n59701;
  assign n59653 = n59702 ^ n59703;
  assign n59688 = ~n59702;
  assign n59656 = ~n59718;
  assign n59698 = n507 ^ n59729;
  assign n59750 = n59765 & n59766;
  assign n59692 = n59770 ^ n59771;
  assign n59767 = n59782 & n59783;
  assign n59769 = n59032 & n57799;
  assign n59739 = ~n59784;
  assign n59743 = ~n59785;
  assign n59768 = n59032 & n59786;
  assign n59794 = n59807 & n59808;
  assign n59544 = ~n58314;
  assign n59617 = n59594 & n11752;
  assign n59593 = n59624 & n59625;
  assign n59615 = ~n59594;
  assign n59643 = ~n59652;
  assign n55758 = n59653 ^ n57059;
  assign n59654 = n59653 & n56994;
  assign n59562 = n59672 & n59673;
  assign n58432 = ~n59678;
  assign n59676 = n59687 & n59688;
  assign n59628 = n59697 ^ n59698;
  assign n59689 = ~n59698;
  assign n59730 = n59692 & n8632;
  assign n59736 = ~n59750;
  assign n59731 = ~n59692;
  assign n59696 = ~n59767;
  assign n59742 = ~n59768;
  assign n59009 = ~n59769;
  assign n59776 = ~n59794;
  assign n59566 = n59593 ^ n59594;
  assign n59600 = n59615 & n40;
  assign n59597 = ~n59593;
  assign n59598 = ~n59617;
  assign n59626 = n55758 & n59640;
  assign n59639 = n55758 & n58249;
  assign n59620 = n59643 & n59644;
  assign n55718 = ~n55758;
  assign n58363 = ~n59654;
  assign n59658 = n59628 & n56970;
  assign n59655 = ~n59676;
  assign n59657 = ~n59628;
  assign n59631 = n59689 & n59690;
  assign n59700 = ~n59730;
  assign n59714 = n59731 & n506;
  assign n59691 = n59736 & n59737;
  assign n59708 = n59742 & n59743;
  assign n59732 = n59776 & n59777;
  assign n59548 = n40 ^ n59566;
  assign n59585 = n59597 & n59598;
  assign n59572 = ~n59600;
  assign n59616 = n59620 & n59621;
  assign n58388 = ~n59626;
  assign n59611 = ~n59639;
  assign n59619 = n55718 & n58414;
  assign n59613 = ~n59620;
  assign n59627 = n59655 & n59656;
  assign n59650 = n59657 & n56968;
  assign n59605 = ~n59658;
  assign n59659 = n59691 ^ n59692;
  assign n59636 = n59708 ^ n59709;
  assign n59699 = ~n59691;
  assign n59664 = ~n59714;
  assign n59694 = n59732 ^ n59733;
  assign n59738 = ~n59732;
  assign n58283 = n59547 ^ n59548;
  assign n59500 = n59548 & n59547;
  assign n59571 = ~n59585;
  assign n59553 = n59611 & n59612;
  assign n59601 = n59613 & n59614;
  assign n59588 = ~n59616;
  assign n58416 = ~n59619;
  assign n59602 = n59627 ^ n59628;
  assign n59629 = ~n59627;
  assign n59630 = ~n59650;
  assign n59632 = n506 ^ n59659;
  assign n59634 = n59693 ^ n59694;
  assign n59677 = n59699 & n59700;
  assign n59715 = n59738 & n59739;
  assign n59499 = ~n58283;
  assign n59549 = n59571 & n59572;
  assign n59590 = n59588 & n59562;
  assign n59589 = n59553 & n59529;
  assign n59586 = ~n59553;
  assign n59569 = ~n59601;
  assign n55665 = n56968 ^ n59602;
  assign n59603 = ~n59602;
  assign n59622 = n59629 & n59630;
  assign n59560 = n59631 ^ n59632;
  assign n59579 = n59632 & n59631;
  assign n59660 = n59634 & n8583;
  assign n59663 = ~n59677;
  assign n59661 = ~n59634;
  assign n59695 = ~n59715;
  assign n59523 = n55 ^ n59549;
  assign n59518 = ~n59549;
  assign n59574 = n59586 & n59587;
  assign n59575 = n59569 & n59588;
  assign n59551 = ~n59589;
  assign n59578 = n55665 & n58232;
  assign n59568 = ~n59590;
  assign n59573 = n55665 & n58353;
  assign n55713 = ~n55665;
  assign n59595 = n59603 & n56968;
  assign n59607 = n59560 & n56988;
  assign n59604 = ~n59622;
  assign n59606 = ~n59560;
  assign n59584 = ~n59579;
  assign n59638 = ~n59660;
  assign n59651 = n59661 & n505;
  assign n59633 = n59663 & n59664;
  assign n59662 = n59695 & n59696;
  assign n59552 = n59568 & n59569;
  assign n58358 = ~n59573;
  assign n59527 = ~n59574;
  assign n59563 = ~n59575;
  assign n59567 = n55713 & n59577;
  assign n59564 = ~n59578;
  assign n58313 = ~n59595;
  assign n59576 = n59604 & n59605;
  assign n59596 = n59606 & n56917;
  assign n59555 = ~n59607;
  assign n59610 = n59633 ^ n59634;
  assign n59637 = ~n59633;
  assign n59609 = ~n59651;
  assign n59635 = n504 ^ n59662;
  assign n59528 = n59552 ^ n59553;
  assign n59524 = n59562 ^ n59563;
  assign n59550 = ~n59552;
  assign n59481 = n59564 & n59565;
  assign n58376 = ~n59567;
  assign n59561 = n59576 ^ n56917;
  assign n59581 = ~n59576;
  assign n59582 = ~n59596;
  assign n59580 = n505 ^ n59610;
  assign n59539 = n59635 ^ n59636;
  assign n59623 = n59637 & n59638;
  assign n59501 = n59523 ^ n59524;
  assign n59479 = n59528 ^ n59529;
  assign n59531 = n59524 & n11714;
  assign n59542 = n59481 & n59545;
  assign n59532 = ~n59524;
  assign n59541 = n59550 & n59551;
  assign n59543 = ~n59481;
  assign n55601 = n59560 ^ n59561;
  assign n59513 = n59579 ^ n59580;
  assign n59570 = n59581 & n59582;
  assign n59583 = ~n59580;
  assign n59608 = ~n59623;
  assign n58240 = n59500 ^ n59501;
  assign n59437 = n59501 & n59500;
  assign n59502 = n59479 & n11658;
  assign n59509 = ~n59479;
  assign n59517 = ~n59531;
  assign n59522 = n59532 & n55;
  assign n59526 = ~n59541;
  assign n59533 = n55601 & n58271;
  assign n59505 = ~n59542;
  assign n59540 = n59543 & n59504;
  assign n59534 = n55601 & n56917;
  assign n59530 = n55601 & n59544;
  assign n55656 = ~n55601;
  assign n59557 = n59513 & n56874;
  assign n59554 = ~n59570;
  assign n59556 = ~n59513;
  assign n59559 = n59583 & n59584;
  assign n59558 = n59608 & n59609;
  assign n59458 = ~n58240;
  assign n59476 = ~n59502;
  assign n59434 = ~n59437;
  assign n59493 = n59509 & n54;
  assign n59515 = n59517 & n59518;
  assign n59498 = ~n59522;
  assign n59503 = n59526 & n59527;
  assign n58319 = ~n59530;
  assign n59519 = ~n59533;
  assign n58288 = ~n59534;
  assign n59521 = n55656 & n58314;
  assign n59486 = ~n59540;
  assign n59535 = n59554 & n59555;
  assign n59546 = n59556 & n56881;
  assign n59537 = ~n59557;
  assign n59538 = n59558 ^ n59559;
  assign n59461 = ~n59493;
  assign n59482 = n59503 ^ n59504;
  assign n59497 = ~n59515;
  assign n59446 = n59519 & n59520;
  assign n59506 = ~n59503;
  assign n58340 = ~n59521;
  assign n59514 = n59535 ^ n56874;
  assign n59470 = n59538 ^ n59539;
  assign n59536 = ~n59535;
  assign n59512 = ~n59546;
  assign n59436 = n59481 ^ n59482;
  assign n59478 = n59497 & n59498;
  assign n59494 = n59505 & n59506;
  assign n59496 = n59446 & n59508;
  assign n59495 = ~n59446;
  assign n55521 = n59513 ^ n59514;
  assign n59510 = n59470 & n56823;
  assign n59516 = ~n59470;
  assign n59525 = n59536 & n59537;
  assign n59464 = n59436 & n53;
  assign n59462 = n59478 ^ n59479;
  assign n59463 = ~n59436;
  assign n59477 = ~n59478;
  assign n59485 = ~n59494;
  assign n59489 = n59495 & n59466;
  assign n59468 = ~n59496;
  assign n59488 = n55521 & n59499;
  assign n55561 = ~n55521;
  assign n59473 = ~n59510;
  assign n59507 = n59516 & n56904;
  assign n59511 = ~n59525;
  assign n59438 = n54 ^ n59462;
  assign n59456 = n59463 & n11582;
  assign n59421 = ~n59464;
  assign n59469 = n59476 & n59477;
  assign n59465 = n59485 & n59486;
  assign n58302 = ~n59488;
  assign n59443 = ~n59489;
  assign n59483 = n55561 & n58136;
  assign n59487 = n55561 & n56874;
  assign n59480 = n55561 & n58283;
  assign n59491 = ~n59507;
  assign n59492 = n59511 & n59512;
  assign n58201 = n59437 ^ n59438;
  assign n59433 = ~n59438;
  assign n59439 = ~n59456;
  assign n59447 = n59465 ^ n59466;
  assign n59460 = ~n59469;
  assign n59467 = ~n59465;
  assign n58277 = ~n59480;
  assign n59474 = ~n59483;
  assign n58247 = ~n59487;
  assign n59471 = n59492 ^ n56823;
  assign n59490 = ~n59492;
  assign n59395 = ~n58201;
  assign n59403 = n59433 & n59434;
  assign n59397 = n59446 ^ n59447;
  assign n59435 = n59460 & n59461;
  assign n59457 = n59467 & n59468;
  assign n55443 = n59470 ^ n59471;
  assign n59408 = n59474 & n59475;
  assign n59484 = n59490 & n59491;
  assign n59422 = n59397 & n52;
  assign n59419 = n59435 ^ n59436;
  assign n59425 = ~n59397;
  assign n59440 = ~n59435;
  assign n59442 = ~n59457;
  assign n59451 = n59408 & n59424;
  assign n59450 = n55443 & n59458;
  assign n59454 = ~n59408;
  assign n55483 = ~n55443;
  assign n59472 = ~n59484;
  assign n59404 = n53 ^ n59419;
  assign n59374 = ~n59422;
  assign n59415 = n59425 & n11500;
  assign n59428 = n59439 & n59440;
  assign n59423 = n59442 & n59443;
  assign n58265 = ~n59450;
  assign n59444 = n55483 & n56904;
  assign n59427 = ~n59451;
  assign n59441 = n55483 & n58240;
  assign n59449 = n59454 & n59455;
  assign n59448 = n55483 & n58191;
  assign n59459 = n59472 & n59473;
  assign n58169 = n59403 ^ n59404;
  assign n59354 = n59404 & n59403;
  assign n59401 = ~n59415;
  assign n59409 = n59423 ^ n59424;
  assign n59420 = ~n59428;
  assign n59426 = ~n59423;
  assign n58243 = ~n59441;
  assign n58209 = ~n59444;
  assign n59429 = ~n59448;
  assign n59406 = ~n59449;
  assign n59453 = n59459 & n56776;
  assign n59452 = ~n59459;
  assign n59364 = ~n58169;
  assign n59358 = n59408 ^ n59409;
  assign n59396 = n59420 & n59421;
  assign n59416 = n59426 & n59427;
  assign n59370 = n59429 & n59430;
  assign n59445 = n59452 & n56771;
  assign n59431 = ~n59453;
  assign n59389 = n59358 & n11429;
  assign n59372 = n59396 ^ n59397;
  assign n59383 = ~n59358;
  assign n59402 = ~n59396;
  assign n59405 = ~n59416;
  assign n59412 = n59370 & n59386;
  assign n59410 = ~n59370;
  assign n59432 = n59431 & n59414;
  assign n59418 = ~n59445;
  assign n59355 = n52 ^ n59372;
  assign n59375 = n59383 & n51;
  assign n59366 = ~n59389;
  assign n59391 = n59401 & n59402;
  assign n59385 = n59405 & n59406;
  assign n59407 = n59410 & n59411;
  assign n59388 = ~n59412;
  assign n59413 = n59418 & n59431;
  assign n59417 = ~n59432;
  assign n58147 = n59354 ^ n59355;
  assign n59309 = n59355 & n59354;
  assign n59341 = ~n59375;
  assign n59371 = n59385 ^ n59386;
  assign n59373 = ~n59391;
  assign n59387 = ~n59385;
  assign n59369 = ~n59407;
  assign n55362 = n59413 ^ n59414;
  assign n59398 = n59417 & n59418;
  assign n59330 = ~n58147;
  assign n59322 = n59370 ^ n59371;
  assign n59357 = n59373 & n59374;
  assign n59378 = n59387 & n59388;
  assign n59390 = n55362 & n59395;
  assign n59392 = n55362 & n58043;
  assign n59393 = n55362 & n56776;
  assign n59376 = n59398 ^ n56697;
  assign n55435 = ~n55362;
  assign n59399 = ~n59398;
  assign n59342 = n59322 & n11352;
  assign n59331 = n59357 ^ n59358;
  assign n59345 = ~n59322;
  assign n59365 = ~n59357;
  assign n55276 = n59376 ^ n59377;
  assign n59368 = ~n59378;
  assign n58203 = ~n59390;
  assign n59384 = n55435 & n58201;
  assign n59381 = ~n59392;
  assign n58164 = ~n59393;
  assign n59394 = n59399 & n59400;
  assign n59310 = n51 ^ n59331;
  assign n59312 = ~n59342;
  assign n59332 = n59345 & n50;
  assign n59349 = n59365 & n59366;
  assign n59356 = n55276 & n58169;
  assign n59346 = n59368 & n59369;
  assign n55339 = ~n55276;
  assign n59325 = n59381 & n59382;
  assign n58223 = ~n59384;
  assign n59379 = ~n59394;
  assign n58087 = n59309 ^ n59310;
  assign n59324 = ~n59310;
  assign n59289 = ~n59332;
  assign n59326 = n59346 ^ n59347;
  assign n59340 = ~n59349;
  assign n58186 = ~n59356;
  assign n59353 = n55339 & n58104;
  assign n59350 = n55339 & n56697;
  assign n59343 = ~n59346;
  assign n59348 = n55339 & n59364;
  assign n59360 = n59325 & n59367;
  assign n59359 = ~n59325;
  assign n59361 = n59379 & n59380;
  assign n59276 = ~n58087;
  assign n59277 = n59324 & n59309;
  assign n59268 = n59325 ^ n59326;
  assign n59321 = n59340 & n59341;
  assign n58166 = ~n59348;
  assign n58125 = ~n59350;
  assign n59333 = ~n59353;
  assign n59351 = n59359 & n59347;
  assign n59344 = ~n59360;
  assign n59338 = n59361 ^ n56607;
  assign n59362 = ~n59361;
  assign n59285 = ~n59277;
  assign n59302 = n59268 & n49;
  assign n59295 = n59321 ^ n59322;
  assign n59297 = ~n59268;
  assign n59311 = ~n59321;
  assign n59282 = n59333 & n59334;
  assign n55154 = n59337 ^ n59338;
  assign n59339 = n59343 & n59344;
  assign n59329 = ~n59351;
  assign n59352 = n59362 & n59363;
  assign n59278 = n50 ^ n59295;
  assign n59290 = n59297 & n11263;
  assign n59254 = ~n59302;
  assign n59306 = n59311 & n59312;
  assign n59313 = n59282 & n59327;
  assign n59314 = n55154 & n57960;
  assign n59315 = n55154 & n56607;
  assign n59323 = n55154 & n59330;
  assign n59320 = ~n59282;
  assign n55310 = ~n55154;
  assign n59328 = ~n59339;
  assign n59335 = ~n59352;
  assign n58067 = n59277 ^ n59278;
  assign n59226 = n59278 & n59285;
  assign n59271 = ~n59290;
  assign n59288 = ~n59306;
  assign n59299 = ~n59313;
  assign n59303 = ~n59314;
  assign n58090 = ~n59315;
  assign n59307 = n59320 & n59301;
  assign n58121 = ~n59323;
  assign n59305 = n55310 & n58147;
  assign n59300 = n59328 & n59329;
  assign n59316 = n59335 & n59336;
  assign n59238 = ~n58067;
  assign n59267 = n59288 & n59289;
  assign n59283 = n59300 ^ n59301;
  assign n59257 = n59303 & n59304;
  assign n58149 = ~n59305;
  assign n59280 = ~n59307;
  assign n59298 = ~n59300;
  assign n59296 = n59316 ^ n59317;
  assign n59318 = ~n59316;
  assign n59246 = n59267 ^ n59268;
  assign n59231 = n59282 ^ n59283;
  assign n59270 = ~n59267;
  assign n59284 = n59257 & n59286;
  assign n59281 = ~n59257;
  assign n55119 = n56731 ^ n59296;
  assign n59291 = n59298 & n59299;
  assign n59292 = ~n59296;
  assign n59308 = n59318 & n59319;
  assign n59227 = n49 ^ n59246;
  assign n59255 = n59231 & n48;
  assign n59264 = n59270 & n59271;
  assign n59260 = ~n59231;
  assign n59273 = n59281 & n59240;
  assign n59272 = n55119 & n57903;
  assign n59266 = n55119 & n58087;
  assign n59259 = ~n59284;
  assign n55192 = ~n55119;
  assign n59279 = ~n59291;
  assign n59287 = n59292 & n56731;
  assign n59293 = ~n59308;
  assign n58009 = n59226 ^ n59227;
  assign n59228 = ~n59227;
  assign n59207 = ~n59255;
  assign n59247 = n59260 & n11173;
  assign n59253 = ~n59264;
  assign n58086 = ~n59266;
  assign n59261 = ~n59272;
  assign n59242 = ~n59273;
  assign n59263 = n55192 & n59276;
  assign n59256 = n59279 & n59280;
  assign n58054 = ~n59287;
  assign n59269 = n59293 & n59294;
  assign n59199 = ~n58009;
  assign n59184 = n59228 & n59226;
  assign n59237 = ~n59247;
  assign n59230 = n59253 & n59254;
  assign n59239 = n59256 ^ n59257;
  assign n59200 = n59261 & n59262;
  assign n58109 = ~n59263;
  assign n59250 = n59269 ^ n56471;
  assign n59258 = ~n59256;
  assign n59274 = ~n59269;
  assign n59204 = n59230 ^ n59231;
  assign n59171 = n59239 ^ n59240;
  assign n59236 = ~n59230;
  assign n59245 = n59200 & n59220;
  assign n59243 = ~n59200;
  assign n54985 = n59249 ^ n59250;
  assign n59248 = n59258 & n59259;
  assign n59265 = n59274 & n59275;
  assign n59185 = n48 ^ n59204;
  assign n59216 = n59171 & n63;
  assign n59215 = ~n59171;
  assign n59222 = n59236 & n59237;
  assign n59229 = n54985 & n58067;
  assign n59232 = n59243 & n59244;
  assign n59217 = ~n59245;
  assign n55104 = ~n54985;
  assign n59241 = ~n59248;
  assign n59251 = ~n59265;
  assign n57972 = n59184 ^ n59185;
  assign n59195 = ~n59185;
  assign n59205 = n59215 & n11134;
  assign n59163 = ~n59216;
  assign n59206 = ~n59222;
  assign n58069 = ~n59229;
  assign n59203 = ~n59232;
  assign n59225 = n55104 & n57844;
  assign n59223 = n55104 & n56674;
  assign n59221 = n55104 & n59238;
  assign n59219 = n59241 & n59242;
  assign n59233 = n59251 & n59252;
  assign n59160 = ~n57972;
  assign n59139 = n59195 & n59184;
  assign n59197 = ~n59205;
  assign n59193 = n59206 & n59207;
  assign n59201 = n59219 ^ n59220;
  assign n58051 = ~n59221;
  assign n58008 = ~n59223;
  assign n59209 = ~n59225;
  assign n59218 = ~n59219;
  assign n59212 = n59233 ^ n56400;
  assign n59234 = ~n59233;
  assign n59170 = n63 ^ n59193;
  assign n59151 = n59200 ^ n59201;
  assign n59196 = ~n59193;
  assign n59154 = n59209 & n59210;
  assign n54992 = n59211 ^ n59212;
  assign n59208 = n59217 & n59218;
  assign n59224 = n59234 & n59235;
  assign n59140 = n59170 ^ n59171;
  assign n59172 = n59151 & n10999;
  assign n59173 = ~n59151;
  assign n59182 = n59196 & n59197;
  assign n59194 = n54992 & n59199;
  assign n59198 = n54992 & n56415;
  assign n59188 = n54992 & n57813;
  assign n59189 = n59154 & n59175;
  assign n54945 = ~n54992;
  assign n59186 = ~n59154;
  assign n59202 = ~n59208;
  assign n59213 = ~n59224;
  assign n57929 = n59139 ^ n59140;
  assign n59142 = ~n59140;
  assign n59153 = ~n59172;
  assign n59164 = n59173 & n62;
  assign n59162 = ~n59182;
  assign n59180 = n59186 & n59187;
  assign n59178 = ~n59188;
  assign n59177 = ~n59189;
  assign n58012 = ~n59194;
  assign n59183 = n54945 & n58009;
  assign n57976 = ~n59198;
  assign n59174 = n59202 & n59203;
  assign n59190 = n59213 & n59214;
  assign n59118 = ~n57929;
  assign n59098 = n59142 & n59139;
  assign n59150 = n59162 & n59163;
  assign n59121 = ~n59164;
  assign n59155 = n59174 ^ n59175;
  assign n59131 = n59178 & n59179;
  assign n59159 = ~n59180;
  assign n58028 = ~n59183;
  assign n59176 = ~n59174;
  assign n59169 = n59190 ^ n56323;
  assign n59191 = ~n59190;
  assign n59107 = ~n59098;
  assign n59119 = n59150 ^ n59151;
  assign n59084 = n59154 ^ n59155;
  assign n59152 = ~n59150;
  assign n59157 = n59131 & n59161;
  assign n59156 = ~n59131;
  assign n54861 = n59168 ^ n59169;
  assign n59165 = n59176 & n59177;
  assign n59181 = n59191 & n59192;
  assign n59099 = n62 ^ n59119;
  assign n59128 = n59084 & n10917;
  assign n59129 = ~n59084;
  assign n59138 = n59152 & n59153;
  assign n59143 = n59156 & n59117;
  assign n59144 = n54861 & n57781;
  assign n59133 = ~n59157;
  assign n59145 = n54861 & n56538;
  assign n59141 = n54861 & n59160;
  assign n54935 = ~n54861;
  assign n59158 = ~n59165;
  assign n59166 = ~n59181;
  assign n57891 = n59098 ^ n59099;
  assign n59106 = ~n59099;
  assign n59109 = ~n59128;
  assign n59122 = n59129 & n61;
  assign n59120 = ~n59138;
  assign n57971 = ~n59141;
  assign n59112 = ~n59143;
  assign n59134 = ~n59144;
  assign n57937 = ~n59145;
  assign n59136 = n54935 & n57972;
  assign n59130 = n59158 & n59159;
  assign n59146 = n59166 & n59167;
  assign n59072 = ~n57891;
  assign n59067 = n59106 & n59107;
  assign n59100 = n59120 & n59121;
  assign n59078 = ~n59122;
  assign n59116 = n59130 ^ n59131;
  assign n59075 = n59134 & n59135;
  assign n57991 = ~n59136;
  assign n59132 = ~n59130;
  assign n59123 = n59146 ^ n59147;
  assign n59148 = ~n59146;
  assign n59083 = n61 ^ n59100;
  assign n59059 = n59116 ^ n59117;
  assign n59110 = ~n59100;
  assign n59115 = n59075 & n59090;
  assign n59113 = ~n59075;
  assign n54834 = n56262 ^ n59123;
  assign n59127 = n59132 & n59133;
  assign n59124 = n59123 & n56466;
  assign n59137 = n59148 & n59149;
  assign n59068 = n59083 ^ n59084;
  assign n59088 = n59059 & n60;
  assign n59087 = ~n59059;
  assign n59096 = n59109 & n59110;
  assign n59101 = n59113 & n59114;
  assign n59105 = n54834 & n57879;
  assign n59092 = ~n59115;
  assign n59108 = n54834 & n59118;
  assign n54786 = ~n54834;
  assign n57898 = ~n59124;
  assign n59111 = ~n59127;
  assign n59125 = ~n59137;
  assign n57850 = n59067 ^ n59068;
  assign n59066 = ~n59068;
  assign n59079 = n59087 & n10873;
  assign n59046 = ~n59088;
  assign n59077 = ~n59096;
  assign n59095 = n54786 & n57929;
  assign n59074 = ~n59101;
  assign n59093 = ~n59105;
  assign n57928 = ~n59108;
  assign n59089 = n59111 & n59112;
  assign n59102 = n59125 & n59126;
  assign n59022 = n59066 & n59067;
  assign n59058 = n59077 & n59078;
  assign n59061 = ~n59079;
  assign n59076 = n59089 ^ n59090;
  assign n59036 = n59093 & n59094;
  assign n57953 = ~n59095;
  assign n59091 = ~n59089;
  assign n59086 = n59102 ^ n56207;
  assign n59103 = ~n59102;
  assign n59025 = ~n59022;
  assign n59040 = n59058 ^ n59059;
  assign n59031 = n59075 ^ n59076;
  assign n59060 = ~n59058;
  assign n59071 = n59036 & n59050;
  assign n59069 = ~n59036;
  assign n54719 = n59085 ^ n59086;
  assign n59080 = n59091 & n59092;
  assign n59097 = n59103 & n59104;
  assign n59023 = n60 ^ n59040;
  assign n59047 = n59031 & n10788;
  assign n59056 = n59060 & n59061;
  assign n59048 = ~n59031;
  assign n59062 = n59069 & n59070;
  assign n59051 = ~n59071;
  assign n59063 = n54719 & n57669;
  assign n59057 = n54719 & n59072;
  assign n59064 = n54719 & n56207;
  assign n54727 = ~n54719;
  assign n59073 = ~n59080;
  assign n59081 = ~n59097;
  assign n59004 = n59022 ^ n59023;
  assign n59024 = ~n59023;
  assign n59027 = ~n59047;
  assign n59041 = n59048 & n59;
  assign n59045 = ~n59056;
  assign n57890 = ~n59057;
  assign n59034 = ~n59062;
  assign n59053 = ~n59063;
  assign n57856 = ~n59064;
  assign n59055 = n54727 & n57891;
  assign n59049 = n59073 & n59074;
  assign n59065 = n59081 & n59082;
  assign n55803 = n56789 ^ n59004;
  assign n58950 = n59004 & n56789;
  assign n59005 = n59004 & n56787;
  assign n58998 = n59024 & n59025;
  assign n59012 = ~n59041;
  assign n59030 = n59045 & n59046;
  assign n59037 = n59049 ^ n59050;
  assign n59002 = n59053 & n59054;
  assign n57916 = ~n59055;
  assign n59052 = ~n59049;
  assign n59044 = n59065 ^ n56353;
  assign n58995 = n55803 & n57838;
  assign n57895 = ~n55803;
  assign n57859 = ~n59005;
  assign n58990 = ~n58998;
  assign n59006 = n59030 ^ n59031;
  assign n58997 = n59036 ^ n59037;
  assign n59026 = ~n59030;
  assign n59035 = n59002 & n59039;
  assign n54686 = n59043 ^ n59044;
  assign n59038 = ~n59002;
  assign n59042 = n59051 & n59052;
  assign n58986 = ~n58995;
  assign n58999 = n59 ^ n59006;
  assign n59018 = n58997 & n10703;
  assign n59019 = n59026 & n59027;
  assign n59015 = ~n58997;
  assign n59017 = ~n59035;
  assign n59028 = n59038 & n59014;
  assign n57836 = ~n54686;
  assign n59033 = ~n59042;
  assign n58969 = n58986 & n58987;
  assign n58983 = n58998 ^ n58999;
  assign n58989 = ~n58999;
  assign n59007 = n59015 & n58;
  assign n58992 = ~n59018;
  assign n59011 = ~n59019;
  assign n59001 = ~n59028;
  assign n59020 = n57836 & n59029;
  assign n59021 = n57836 & n59032;
  assign n59013 = n59033 & n59034;
  assign n58958 = n58969 ^ n58970;
  assign n58973 = ~n58969;
  assign n58976 = n58983 & n56680;
  assign n58977 = ~n58983;
  assign n58963 = n58989 & n58990;
  assign n58979 = ~n59007;
  assign n58996 = n59011 & n59012;
  assign n59003 = n59013 ^ n59014;
  assign n59008 = ~n59020;
  assign n57820 = ~n59021;
  assign n59016 = ~n59013;
  assign n57417 = n199 ^ n58958;
  assign n58850 = n58958 & n199;
  assign n58899 = n58973 & n58974;
  assign n58961 = ~n58976;
  assign n58975 = n58977 & n56673;
  assign n58980 = n58996 ^ n58997;
  assign n58965 = n59002 ^ n59003;
  assign n58991 = ~n58996;
  assign n58993 = n59008 & n59009;
  assign n59010 = n59016 & n59017;
  assign n58681 = ~n57417;
  assign n58960 = n58961 & n58950;
  assign n58957 = ~n58975;
  assign n58966 = n58 ^ n58980;
  assign n58985 = n58965 & n57;
  assign n58988 = n58991 & n58992;
  assign n58982 = ~n58965;
  assign n58972 = n58993 ^ n58994;
  assign n59000 = ~n59010;
  assign n58956 = ~n58960;
  assign n58949 = n58961 & n58957;
  assign n58938 = n58963 ^ n58966;
  assign n58962 = ~n58966;
  assign n58981 = n58982 & n10623;
  assign n58954 = ~n58985;
  assign n58978 = ~n58988;
  assign n58984 = n59000 & n59001;
  assign n55646 = n58949 ^ n58950;
  assign n58947 = n58956 & n58957;
  assign n58951 = n58938 & n56610;
  assign n58955 = ~n58938;
  assign n58945 = n58962 & n58963;
  assign n58964 = n58978 & n58979;
  assign n58967 = ~n58981;
  assign n58971 = n56 ^ n58984;
  assign n58942 = n55646 & n56680;
  assign n58939 = n58947 ^ n56610;
  assign n58941 = n55646 & n57756;
  assign n55784 = ~n55646;
  assign n58933 = ~n58951;
  assign n58944 = ~n58947;
  assign n58948 = n58955 & n56568;
  assign n58952 = n58964 ^ n58965;
  assign n58929 = n58971 ^ n58972;
  assign n58968 = ~n58964;
  assign n55611 = n58938 ^ n58939;
  assign n58934 = ~n58941;
  assign n57773 = ~n58942;
  assign n58943 = ~n58948;
  assign n58946 = n57 ^ n58952;
  assign n58959 = n58967 & n58968;
  assign n55613 = ~n55611;
  assign n58930 = n58934 & n58935;
  assign n58940 = n58943 & n58944;
  assign n58908 = n58945 ^ n58946;
  assign n58936 = n58946 & n58945;
  assign n58953 = ~n58959;
  assign n58922 = n55613 & n56568;
  assign n58923 = n55613 & n57704;
  assign n58925 = n58930 & n58931;
  assign n58926 = ~n58930;
  assign n58932 = ~n58940;
  assign n58914 = ~n58908;
  assign n58937 = n58953 & n58954;
  assign n57734 = ~n58922;
  assign n58916 = ~n58923;
  assign n58910 = ~n58925;
  assign n58924 = n58926 & n58927;
  assign n58919 = n58932 & n58933;
  assign n58928 = n58936 ^ n58937;
  assign n58874 = n58916 & n58917;
  assign n58915 = n58910 & n58899;
  assign n58909 = n58919 ^ n56523;
  assign n58905 = ~n58924;
  assign n58921 = n58919 & n56555;
  assign n58872 = n58928 ^ n58929;
  assign n58920 = ~n58919;
  assign n58897 = n58874 & n58903;
  assign n55502 = n58908 ^ n58909;
  assign n58902 = ~n58874;
  assign n58898 = n58905 & n58910;
  assign n58904 = ~n58915;
  assign n58912 = n58872 & n56457;
  assign n58911 = ~n58872;
  assign n58918 = n58920 & n56523;
  assign n58913 = ~n58921;
  assign n58890 = ~n58897;
  assign n58895 = n55502 & n56555;
  assign n58889 = n58898 ^ n58899;
  assign n58896 = n55502 & n57631;
  assign n58894 = n58902 & n58893;
  assign n55508 = ~n55502;
  assign n58892 = n58904 & n58905;
  assign n58906 = n58911 & n56440;
  assign n58871 = ~n58912;
  assign n58907 = n58913 & n58914;
  assign n58901 = ~n58918;
  assign n58884 = n58889 & n198;
  assign n58875 = n58892 ^ n58893;
  assign n58877 = ~n58894;
  assign n57662 = ~n58895;
  assign n58882 = ~n58896;
  assign n58888 = ~n58889;
  assign n58891 = ~n58892;
  assign n58887 = ~n58906;
  assign n58900 = ~n58907;
  assign n58836 = n58874 ^ n58875;
  assign n58845 = n58882 & n58883;
  assign n58857 = ~n58884;
  assign n58879 = n58888 & n8617;
  assign n58881 = n58890 & n58891;
  assign n58885 = n58900 & n58901;
  assign n58860 = n58836 & n197;
  assign n58859 = ~n58836;
  assign n58869 = n58845 & n58878;
  assign n58868 = ~n58845;
  assign n58867 = ~n58879;
  assign n58876 = ~n58881;
  assign n58873 = n58885 ^ n56440;
  assign n58886 = ~n58885;
  assign n58848 = n58859 & n8554;
  assign n58822 = ~n58860;
  assign n58865 = n58867 & n58850;
  assign n58866 = n58868 & n58862;
  assign n58849 = n58867 & n58857;
  assign n58863 = ~n58869;
  assign n55459 = n58872 ^ n58873;
  assign n58861 = n58876 & n58877;
  assign n58880 = n58886 & n58887;
  assign n58833 = ~n58848;
  assign n57379 = n58849 ^ n58850;
  assign n58846 = n58861 ^ n58862;
  assign n58858 = n55459 & n56440;
  assign n58852 = n55459 & n57560;
  assign n58856 = ~n58865;
  assign n58844 = ~n58866;
  assign n55382 = ~n55459;
  assign n58864 = ~n58861;
  assign n58870 = ~n58880;
  assign n58801 = n58845 ^ n58846;
  assign n58646 = ~n57379;
  assign n58841 = ~n58852;
  assign n58835 = n58856 & n58857;
  assign n57615 = ~n58858;
  assign n58851 = n58863 & n58864;
  assign n58853 = n58870 & n58871;
  assign n58825 = n58801 & n196;
  assign n58824 = ~n58801;
  assign n58819 = n58835 ^ n58836;
  assign n58810 = n58841 & n58842;
  assign n58834 = ~n58835;
  assign n58843 = ~n58851;
  assign n58840 = n58853 ^ n56365;
  assign n58854 = ~n58853;
  assign n57349 = n197 ^ n58819;
  assign n58823 = n58824 & n8495;
  assign n58788 = ~n58825;
  assign n58832 = n58833 & n58834;
  assign n58814 = ~n58810;
  assign n55312 = n58839 ^ n58840;
  assign n58826 = n58843 & n58844;
  assign n58847 = n58854 & n58855;
  assign n58607 = ~n57349;
  assign n58804 = ~n58823;
  assign n58811 = n58826 ^ n58827;
  assign n58815 = n55312 & n57538;
  assign n58816 = n55312 & n56365;
  assign n58831 = n58826 & n58827;
  assign n55348 = ~n55312;
  assign n58821 = ~n58832;
  assign n58828 = ~n58826;
  assign n58837 = ~n58847;
  assign n58771 = n58810 ^ n58811;
  assign n58807 = ~n58815;
  assign n57553 = ~n58816;
  assign n58800 = n58821 & n58822;
  assign n58820 = n58828 & n58829;
  assign n58813 = ~n58831;
  assign n58830 = n58837 & n58838;
  assign n58789 = n58771 & n8474;
  assign n58795 = ~n58771;
  assign n58786 = n58800 ^ n58801;
  assign n58762 = n58807 & n58808;
  assign n58805 = ~n58800;
  assign n58806 = n58813 & n58814;
  assign n58798 = ~n58820;
  assign n58818 = n58830 & n56306;
  assign n58817 = ~n58830;
  assign n57312 = n196 ^ n58786;
  assign n58772 = ~n58789;
  assign n58784 = n58795 & n195;
  assign n58792 = n58762 & n58783;
  assign n58790 = ~n58762;
  assign n58796 = n58804 & n58805;
  assign n58797 = ~n58806;
  assign n58812 = n58817 & n56297;
  assign n58803 = ~n58818;
  assign n58567 = ~n57312;
  assign n58754 = ~n58784;
  assign n58785 = n58790 & n58791;
  assign n58778 = ~n58792;
  assign n58787 = ~n58796;
  assign n58782 = n58797 & n58798;
  assign n58802 = n58803 & n58809;
  assign n58794 = ~n58812;
  assign n58763 = n58782 ^ n58783;
  assign n58766 = ~n58785;
  assign n58770 = n58787 & n58788;
  assign n58779 = ~n58782;
  assign n58793 = ~n58802;
  assign n58799 = n58794 & n58803;
  assign n58735 = n58762 ^ n58763;
  assign n58752 = n58770 ^ n58771;
  assign n58773 = ~n58770;
  assign n58774 = n58778 & n58779;
  assign n58775 = n58793 & n58794;
  assign n58781 = ~n58799;
  assign n57282 = n195 ^ n58752;
  assign n58746 = n58735 & n8425;
  assign n58747 = ~n58735;
  assign n58764 = n58772 & n58773;
  assign n58765 = ~n58774;
  assign n58760 = n58775 ^ n56237;
  assign n55195 = n58780 ^ n58781;
  assign n58776 = ~n58775;
  assign n58732 = ~n58746;
  assign n58739 = n58747 & n194;
  assign n58528 = ~n57282;
  assign n55140 = n58760 ^ n58761;
  assign n58753 = ~n58764;
  assign n58748 = n58765 & n58766;
  assign n58767 = n55195 & n57481;
  assign n58768 = n55195 & n56306;
  assign n58769 = n58776 & n58777;
  assign n55266 = ~n55195;
  assign n58721 = ~n58739;
  assign n58731 = n58748 ^ n58749;
  assign n58742 = n55140 & n56237;
  assign n58741 = n55140 & n57446;
  assign n58734 = n58753 & n58754;
  assign n55191 = ~n55140;
  assign n58750 = n58748 & n58757;
  assign n58751 = ~n58748;
  assign n58755 = ~n58767;
  assign n57502 = ~n58768;
  assign n58758 = ~n58769;
  assign n58716 = n58734 ^ n58735;
  assign n58726 = ~n58741;
  assign n57459 = ~n58742;
  assign n58736 = ~n58750;
  assign n58740 = n58751 & n58749;
  assign n58733 = ~n58734;
  assign n58730 = n58755 & n58756;
  assign n58743 = n58758 & n58759;
  assign n57240 = n194 ^ n58716;
  assign n58685 = n58726 & n58727;
  assign n58698 = n58730 ^ n58731;
  assign n58728 = n58732 & n58733;
  assign n58718 = ~n58740;
  assign n58723 = n58743 ^ n56136;
  assign n58737 = ~n58730;
  assign n58744 = ~n58743;
  assign n58484 = ~n57240;
  assign n58713 = n58685 & n58719;
  assign n58714 = n58698 & n193;
  assign n58715 = ~n58698;
  assign n58712 = ~n58685;
  assign n55046 = n58722 ^ n58723;
  assign n58720 = ~n58728;
  assign n58729 = n58736 & n58737;
  assign n58738 = n58744 & n58745;
  assign n58707 = n58712 & n58700;
  assign n58701 = ~n58713;
  assign n58680 = ~n58714;
  assign n58706 = n58715 & n8392;
  assign n55099 = ~n55046;
  assign n58697 = n58720 & n58721;
  assign n58717 = ~n58729;
  assign n58724 = ~n58738;
  assign n58684 = n58697 ^ n58698;
  assign n58695 = ~n58706;
  assign n58683 = ~n58707;
  assign n58704 = n55099 & n56160;
  assign n58703 = n55099 & n57393;
  assign n58696 = ~n58697;
  assign n58699 = n58717 & n58718;
  assign n58708 = n58724 & n58725;
  assign n57179 = n193 ^ n58684;
  assign n58687 = n58695 & n58696;
  assign n58686 = n58699 ^ n58700;
  assign n58688 = ~n58703;
  assign n57420 = ~n58704;
  assign n58690 = n58708 ^ n58709;
  assign n58702 = ~n58699;
  assign n58710 = ~n58708;
  assign n58614 = ~n57179;
  assign n58677 = n58685 ^ n58686;
  assign n58679 = ~n58687;
  assign n58651 = n58688 & n58689;
  assign n54957 = n58690 ^ n56080;
  assign n58693 = n58690 & n56080;
  assign n58694 = n58701 & n58702;
  assign n58705 = n58710 & n58711;
  assign n58669 = n58677 & n192;
  assign n58636 = n58679 & n58680;
  assign n58673 = n54957 & n58681;
  assign n58671 = ~n58677;
  assign n54976 = ~n54957;
  assign n58661 = ~n58651;
  assign n57389 = ~n58693;
  assign n58682 = ~n58694;
  assign n58691 = ~n58705;
  assign n58628 = ~n58669;
  assign n58662 = n58671 & n8358;
  assign n57441 = ~n58673;
  assign n58667 = n54976 & n57417;
  assign n58668 = n54976 & n57346;
  assign n58650 = ~n58636;
  assign n58664 = n58682 & n58683;
  assign n58674 = n58691 & n58692;
  assign n58649 = ~n58662;
  assign n58652 = n58664 ^ n58665;
  assign n57416 = ~n58667;
  assign n58658 = ~n58668;
  assign n58655 = n58674 ^ n56041;
  assign n58666 = n58664 & n58678;
  assign n58672 = ~n58664;
  assign n58675 = ~n58674;
  assign n58647 = n58649 & n58650;
  assign n58609 = n58651 ^ n58652;
  assign n58635 = n58649 & n58628;
  assign n54897 = n58654 ^ n58655;
  assign n58596 = n58658 & n58659;
  assign n58660 = ~n58666;
  assign n58663 = n58672 & n58665;
  assign n58670 = n58675 & n58676;
  assign n58615 = n58635 ^ n58636;
  assign n58629 = n58609 & n207;
  assign n58637 = ~n58609;
  assign n58640 = n54897 & n58646;
  assign n58627 = ~n58647;
  assign n58639 = n58596 & n58648;
  assign n58638 = ~n58596;
  assign n54872 = ~n54897;
  assign n58653 = n58660 & n58661;
  assign n58643 = ~n58663;
  assign n58656 = ~n58670;
  assign n57172 = n58615 ^ n57179;
  assign n58613 = ~n58615;
  assign n58608 = n58627 & n58628;
  assign n58595 = ~n58629;
  assign n58626 = n58637 & n8317;
  assign n58632 = n54872 & n57309;
  assign n58630 = n58638 & n58617;
  assign n58619 = ~n58639;
  assign n58631 = n54872 & n56058;
  assign n57409 = ~n58640;
  assign n58633 = n54872 & n57379;
  assign n58642 = ~n58653;
  assign n58641 = n58656 & n58657;
  assign n58420 = ~n57172;
  assign n58593 = n58608 ^ n58609;
  assign n58571 = n58613 & n58614;
  assign n58611 = ~n58626;
  assign n58612 = ~n58608;
  assign n58599 = ~n58630;
  assign n57352 = ~n58631;
  assign n58622 = ~n58632;
  assign n57382 = ~n58633;
  assign n58625 = n58641 ^ n56000;
  assign n58616 = n58642 & n58643;
  assign n58644 = ~n58641;
  assign n58572 = n207 ^ n58593;
  assign n58577 = ~n58571;
  assign n58606 = n58611 & n58612;
  assign n58597 = n58616 ^ n58617;
  assign n58563 = n58622 & n58623;
  assign n54777 = n58624 ^ n58625;
  assign n58618 = ~n58616;
  assign n58634 = n58644 & n58645;
  assign n57134 = n58571 ^ n58572;
  assign n58535 = n58572 & n58577;
  assign n58576 = n58596 ^ n58597;
  assign n58594 = ~n58606;
  assign n58600 = n54777 & n57277;
  assign n58602 = n54777 & n56005;
  assign n58601 = n54777 & n58607;
  assign n58570 = ~n58563;
  assign n54828 = ~n54777;
  assign n58610 = n58618 & n58619;
  assign n58620 = ~n58634;
  assign n58374 = ~n57134;
  assign n58586 = n58576 & n206;
  assign n58583 = ~n58576;
  assign n58575 = n58594 & n58595;
  assign n58589 = ~n58600;
  assign n57348 = ~n58601;
  assign n57320 = ~n58602;
  assign n58592 = n54828 & n57349;
  assign n58598 = ~n58610;
  assign n58603 = n58620 & n58621;
  assign n58552 = n58575 ^ n58576;
  assign n58573 = n58583 & n8278;
  assign n58544 = ~n58586;
  assign n58513 = n58589 & n58590;
  assign n58554 = ~n58575;
  assign n57368 = ~n58592;
  assign n58578 = n58598 & n58599;
  assign n58581 = n58603 ^ n55947;
  assign n58604 = ~n58603;
  assign n58536 = n206 ^ n58552;
  assign n58553 = ~n58573;
  assign n58568 = n58513 & n58531;
  assign n58564 = n58578 ^ n58579;
  assign n54708 = n58581 ^ n58582;
  assign n58565 = ~n58513;
  assign n58580 = n58578 & n58579;
  assign n58587 = ~n58578;
  assign n58591 = n58604 & n58605;
  assign n57072 = n58535 ^ n58536;
  assign n58487 = n58536 & n58535;
  assign n58549 = n58553 & n58554;
  assign n58519 = n58563 ^ n58564;
  assign n58556 = n58565 & n58566;
  assign n58557 = n54708 & n58567;
  assign n58533 = ~n58568;
  assign n58558 = n54708 & n57265;
  assign n58559 = n54708 & n55947;
  assign n54728 = ~n54708;
  assign n58569 = ~n58580;
  assign n58574 = n58587 & n58588;
  assign n58584 = ~n58591;
  assign n58336 = ~n57072;
  assign n58500 = ~n58487;
  assign n58537 = n58519 & n8239;
  assign n58543 = ~n58549;
  assign n58542 = ~n58519;
  assign n58510 = ~n58556;
  assign n57315 = ~n58557;
  assign n58545 = ~n58558;
  assign n57288 = ~n58559;
  assign n58550 = n54728 & n57312;
  assign n58555 = n58569 & n58570;
  assign n58548 = ~n58574;
  assign n58562 = n58584 & n58585;
  assign n58521 = ~n58537;
  assign n58534 = n58542 & n205;
  assign n58518 = n58543 & n58544;
  assign n58465 = n58545 & n58546;
  assign n57331 = ~n58550;
  assign n58547 = ~n58555;
  assign n58540 = n58562 ^ n55929;
  assign n58560 = ~n58562;
  assign n58502 = n58518 ^ n58519;
  assign n58520 = ~n58518;
  assign n58504 = ~n58534;
  assign n58472 = ~n58465;
  assign n54625 = n58540 ^ n58541;
  assign n58530 = n58547 & n58548;
  assign n58551 = n58560 & n58561;
  assign n58488 = n205 ^ n58502;
  assign n58517 = n58520 & n58521;
  assign n58514 = n58530 ^ n58531;
  assign n58523 = n54625 & n57202;
  assign n58525 = n54625 & n55929;
  assign n58524 = n54625 & n57282;
  assign n54631 = ~n54625;
  assign n58532 = ~n58530;
  assign n58538 = ~n58551;
  assign n57031 = n58487 ^ n58488;
  assign n58452 = n58488 & n58500;
  assign n58490 = n58513 ^ n58514;
  assign n58503 = ~n58517;
  assign n58511 = ~n58523;
  assign n57279 = ~n58524;
  assign n57248 = ~n58525;
  assign n58515 = n54631 & n58528;
  assign n58522 = n58532 & n58533;
  assign n58529 = n58538 & n58539;
  assign n58303 = ~n57031;
  assign n58499 = n58490 & n8227;
  assign n58489 = n58503 & n58504;
  assign n58497 = ~n58490;
  assign n58427 = n58511 & n58512;
  assign n57296 = ~n58515;
  assign n58509 = ~n58522;
  assign n58508 = n58529 ^ n55879;
  assign n58526 = ~n58529;
  assign n58460 = n58489 ^ n58490;
  assign n58477 = n58497 & n204;
  assign n58475 = ~n58499;
  assign n58496 = n58427 & n58444;
  assign n58476 = ~n58489;
  assign n58494 = ~n58427;
  assign n54582 = n58507 ^ n58508;
  assign n58491 = n58509 & n58510;
  assign n58516 = n58526 & n58527;
  assign n58453 = n204 ^ n58460;
  assign n58470 = n58475 & n58476;
  assign n58457 = ~n58477;
  assign n58466 = n58491 ^ n58492;
  assign n58479 = n58494 & n58495;
  assign n58446 = ~n58496;
  assign n58481 = n54582 & n57240;
  assign n58480 = n54582 & n57187;
  assign n58482 = n54582 & n55879;
  assign n58498 = n58491 & n58501;
  assign n54545 = ~n54582;
  assign n58493 = ~n58491;
  assign n58505 = ~n58516;
  assign n56998 = n58452 ^ n58453;
  assign n58407 = n58453 & n58452;
  assign n58439 = n58465 ^ n58466;
  assign n58456 = ~n58470;
  assign n58425 = ~n58479;
  assign n58468 = ~n58480;
  assign n57239 = ~n58481;
  assign n57206 = ~n58482;
  assign n58473 = n54545 & n58484;
  assign n58478 = n58493 & n58492;
  assign n58471 = ~n58498;
  assign n58483 = n58505 & n58506;
  assign n58257 = ~n56998;
  assign n58418 = ~n58407;
  assign n58438 = n58456 & n58457;
  assign n58454 = n58439 & n203;
  assign n58455 = ~n58439;
  assign n58381 = n58468 & n58469;
  assign n58467 = n58471 & n58472;
  assign n57261 = ~n58473;
  assign n58459 = ~n58478;
  assign n58462 = n58483 ^ n55818;
  assign n58485 = ~n58483;
  assign n58426 = n58438 ^ n58439;
  assign n58437 = ~n58438;
  assign n58422 = ~n58454;
  assign n58447 = n58455 & n8167;
  assign n58391 = ~n58381;
  assign n54530 = n58461 ^ n58462;
  assign n58458 = ~n58467;
  assign n58474 = n58485 & n58486;
  assign n58408 = n203 ^ n58426;
  assign n58436 = ~n58447;
  assign n54496 = ~n54530;
  assign n58443 = n58458 & n58459;
  assign n58463 = ~n58474;
  assign n56951 = n58407 ^ n58408;
  assign n58359 = n58408 & n58418;
  assign n58429 = n58436 & n58437;
  assign n58428 = n58443 ^ n58444;
  assign n58441 = n54496 & n57105;
  assign n58440 = n54496 & n55850;
  assign n58445 = ~n58443;
  assign n58448 = n58463 & n58464;
  assign n58224 = ~n56951;
  assign n58397 = n58427 ^ n58428;
  assign n58421 = ~n58429;
  assign n57141 = ~n58440;
  assign n58433 = ~n58441;
  assign n58435 = n58445 & n58446;
  assign n58430 = n58448 ^ n58449;
  assign n58450 = ~n58448;
  assign n58400 = n58397 & n8128;
  assign n58396 = n58421 & n58422;
  assign n58404 = ~n58397;
  assign n54449 = n55810 ^ n58430;
  assign n58331 = n58433 & n58434;
  assign n58424 = ~n58435;
  assign n58442 = n58450 & n58451;
  assign n58379 = n58396 ^ n58397;
  assign n58384 = ~n58400;
  assign n58392 = n58404 & n202;
  assign n58385 = ~n58396;
  assign n58410 = n54449 & n58420;
  assign n58411 = n54449 & n57110;
  assign n58412 = n54449 & n55810;
  assign n58409 = n58331 & n58423;
  assign n58401 = n58424 & n58425;
  assign n54510 = ~n54449;
  assign n58417 = ~n58331;
  assign n58431 = ~n58442;
  assign n58360 = n202 ^ n58379;
  assign n58380 = n58384 & n58385;
  assign n58378 = ~n58392;
  assign n58382 = n58401 ^ n58399;
  assign n58352 = ~n58409;
  assign n57174 = ~n58410;
  assign n58394 = ~n58411;
  assign n57119 = ~n58412;
  assign n58405 = n54510 & n57172;
  assign n58403 = n58417 & n58350;
  assign n58402 = n58401 & n58419;
  assign n58398 = ~n58401;
  assign n58413 = n58431 & n58432;
  assign n56922 = n58359 ^ n58360;
  assign n58364 = ~n58360;
  assign n58377 = ~n58380;
  assign n58356 = n58381 ^ n58382;
  assign n58282 = n58394 & n58395;
  assign n58393 = n58398 & n58399;
  assign n58390 = ~n58402;
  assign n58334 = ~n58403;
  assign n57156 = ~n58405;
  assign n58386 = n58413 ^ n58414;
  assign n58415 = ~n58413;
  assign n58192 = ~n56922;
  assign n58308 = n58364 & n58359;
  assign n58365 = n58356 & n201;
  assign n58355 = n58377 & n58378;
  assign n58368 = ~n58356;
  assign n54420 = n55758 ^ n58386;
  assign n58383 = n58390 & n58391;
  assign n58373 = ~n58393;
  assign n58389 = n58386 & n55718;
  assign n58406 = n58415 & n58416;
  assign n58341 = n58355 ^ n58356;
  assign n58317 = ~n58308;
  assign n58346 = ~n58355;
  assign n58326 = ~n58365;
  assign n58361 = n58368 & n8107;
  assign n58369 = n54420 & n57059;
  assign n58370 = n54420 & n57134;
  assign n54433 = ~n54420;
  assign n58372 = ~n58383;
  assign n57080 = ~n58389;
  assign n58387 = ~n58406;
  assign n58309 = n201 ^ n58341;
  assign n58345 = ~n58361;
  assign n58362 = ~n58369;
  assign n57115 = ~n58370;
  assign n58349 = n58372 & n58373;
  assign n58366 = n54433 & n58374;
  assign n58371 = n58387 & n58388;
  assign n56878 = n58308 ^ n58309;
  assign n58316 = ~n58309;
  assign n58342 = n58345 & n58346;
  assign n58332 = n58349 ^ n58350;
  assign n58273 = n58362 & n58363;
  assign n58351 = ~n58349;
  assign n57132 = ~n58366;
  assign n58354 = n58371 ^ n55665;
  assign n58375 = ~n58371;
  assign n58153 = ~n56878;
  assign n58274 = n58316 & n58317;
  assign n58305 = n58331 ^ n58332;
  assign n58325 = ~n58342;
  assign n58344 = n58273 & n58347;
  assign n58348 = n58351 & n58352;
  assign n58343 = ~n58273;
  assign n54370 = n58353 ^ n58354;
  assign n58367 = n58375 & n58376;
  assign n58280 = ~n58274;
  assign n58310 = n58305 & n200;
  assign n58304 = n58325 & n58326;
  assign n58322 = ~n58305;
  assign n58335 = n58343 & n58249;
  assign n58269 = ~n58344;
  assign n58337 = n54370 & n57072;
  assign n54411 = ~n54370;
  assign n58333 = ~n58348;
  assign n58357 = ~n58367;
  assign n58289 = n58304 ^ n58305;
  assign n58279 = ~n58310;
  assign n58306 = n58322 & n8067;
  assign n58299 = ~n58304;
  assign n58323 = n58333 & n58334;
  assign n58251 = ~n58335;
  assign n58327 = n54411 & n58336;
  assign n57093 = ~n58337;
  assign n58328 = n54411 & n56970;
  assign n58329 = n54411 & n55713;
  assign n58338 = n58357 & n58358;
  assign n58275 = n200 ^ n58289;
  assign n58298 = ~n58306;
  assign n58311 = n58323 & n58324;
  assign n58320 = ~n58323;
  assign n57071 = ~n58327;
  assign n58312 = ~n58328;
  assign n57036 = ~n58329;
  assign n58315 = n58338 ^ n55601;
  assign n58339 = ~n58338;
  assign n56836 = n58274 ^ n58275;
  assign n58215 = n58275 & n58280;
  assign n58290 = n58298 & n58299;
  assign n58300 = ~n58311;
  assign n58205 = n58312 & n58313;
  assign n54327 = n58314 ^ n58315;
  assign n58307 = n58320 & n58321;
  assign n58330 = n58339 & n58340;
  assign n58112 = ~n56836;
  assign n58226 = ~n58215;
  assign n58278 = ~n58290;
  assign n58293 = n58300 & n58282;
  assign n58294 = n54327 & n58303;
  assign n58296 = n54327 & n55656;
  assign n58295 = n54327 & n56988;
  assign n58213 = ~n58205;
  assign n54373 = ~n54327;
  assign n58286 = ~n58307;
  assign n58318 = ~n58330;
  assign n58262 = n58278 & n58279;
  assign n58285 = ~n58293;
  assign n57034 = ~n58294;
  assign n58287 = ~n58295;
  assign n57002 = ~n58296;
  assign n58281 = n58286 & n58300;
  assign n58291 = n54373 & n57031;
  assign n58297 = n58318 & n58319;
  assign n58244 = n215 ^ n58262;
  assign n58239 = ~n58262;
  assign n58245 = n58281 ^ n58282;
  assign n58272 = n58285 & n58286;
  assign n58154 = n58287 & n58288;
  assign n57055 = ~n58291;
  assign n58284 = n58297 ^ n55521;
  assign n58301 = ~n58297;
  assign n58216 = n58244 ^ n58245;
  assign n58263 = n58245 & n215;
  assign n58248 = n58272 ^ n58273;
  assign n58266 = ~n58245;
  assign n58267 = n58154 & n58173;
  assign n58270 = ~n58154;
  assign n54329 = n58283 ^ n58284;
  assign n58268 = ~n58272;
  assign n58292 = n58301 & n58302;
  assign n56812 = n58215 ^ n58216;
  assign n58225 = ~n58216;
  assign n58197 = n58248 ^ n58249;
  assign n58228 = ~n58263;
  assign n58252 = n58266 & n8015;
  assign n58258 = n54329 & n56881;
  assign n58178 = ~n58267;
  assign n58259 = n54329 & n55521;
  assign n58260 = n54329 & n56998;
  assign n58255 = n58268 & n58269;
  assign n58256 = n58270 & n58271;
  assign n54290 = ~n54329;
  assign n58276 = ~n58292;
  assign n58075 = ~n56812;
  assign n58159 = n58225 & n58226;
  assign n58230 = n58197 & n214;
  assign n58235 = ~n58197;
  assign n58238 = ~n58252;
  assign n58250 = ~n58255;
  assign n58158 = ~n58256;
  assign n58253 = n54290 & n58257;
  assign n58246 = ~n58258;
  assign n56959 = ~n58259;
  assign n56996 = ~n58260;
  assign n58261 = n58276 & n58277;
  assign n58188 = ~n58230;
  assign n58229 = n58235 & n7981;
  assign n58236 = n58238 & n58239;
  assign n58114 = n58246 & n58247;
  assign n58231 = n58250 & n58251;
  assign n57021 = ~n58253;
  assign n58241 = n58261 ^ n55443;
  assign n58264 = ~n58261;
  assign n58204 = ~n58229;
  assign n58206 = n58231 ^ n58232;
  assign n58227 = ~n58236;
  assign n58234 = n58231 & n58237;
  assign n58127 = ~n58114;
  assign n54259 = n58240 ^ n58241;
  assign n58233 = ~n58231;
  assign n58254 = n58264 & n58265;
  assign n58168 = n58205 ^ n58206;
  assign n58210 = n58227 & n58228;
  assign n58217 = n58233 & n58232;
  assign n58212 = ~n58234;
  assign n58221 = n54259 & n56951;
  assign n58219 = n54259 & n55443;
  assign n58218 = n54259 & n56823;
  assign n54257 = ~n54259;
  assign n58242 = ~n58254;
  assign n58189 = n58168 & n213;
  assign n58194 = ~n58168;
  assign n58196 = ~n58210;
  assign n58207 = n58212 & n58213;
  assign n58199 = ~n58217;
  assign n58208 = ~n58218;
  assign n56921 = ~n58219;
  assign n56954 = ~n58221;
  assign n58211 = n54257 & n58224;
  assign n58220 = n58242 & n58243;
  assign n58152 = ~n58189;
  assign n58181 = n58194 & n7930;
  assign n58180 = n58196 ^ n58197;
  assign n58195 = n58204 & n58196;
  assign n58198 = ~n58207;
  assign n58070 = n58208 & n58209;
  assign n56981 = ~n58211;
  assign n58200 = n58220 ^ n55435;
  assign n58222 = ~n58220;
  assign n58160 = n214 ^ n58180;
  assign n58161 = ~n58181;
  assign n58187 = ~n58195;
  assign n58193 = n58070 & n58082;
  assign n58172 = n58198 & n58199;
  assign n58190 = ~n58070;
  assign n54196 = n58200 ^ n58201;
  assign n58214 = n58222 & n58223;
  assign n56736 = n58159 ^ n58160;
  assign n58122 = n58160 & n58159;
  assign n58155 = n58172 ^ n58173;
  assign n58167 = n58187 & n58188;
  assign n58177 = ~n58172;
  assign n58182 = n58190 & n58191;
  assign n58183 = n54196 & n58192;
  assign n58084 = ~n58193;
  assign n54232 = ~n54196;
  assign n58202 = ~n58214;
  assign n58035 = ~n56736;
  assign n58130 = n58154 ^ n58155;
  assign n58144 = n58167 ^ n58168;
  assign n58171 = n58177 & n58178;
  assign n58162 = ~n58167;
  assign n58073 = ~n58182;
  assign n58176 = n54232 & n56771;
  assign n56942 = ~n58183;
  assign n58174 = n54232 & n56922;
  assign n58179 = n54232 & n55435;
  assign n58184 = n58202 & n58203;
  assign n58123 = n213 ^ n58144;
  assign n58134 = n58130 & n7900;
  assign n58141 = ~n58130;
  assign n58156 = n58161 & n58162;
  assign n58157 = ~n58171;
  assign n56925 = ~n58174;
  assign n58163 = ~n58176;
  assign n56885 = ~n58179;
  assign n58170 = n58184 ^ n55276;
  assign n58185 = ~n58184;
  assign n56710 = n58122 ^ n58123;
  assign n58131 = ~n58123;
  assign n58117 = ~n58134;
  assign n58132 = n58141 & n212;
  assign n58151 = ~n58156;
  assign n58135 = n58157 & n58158;
  assign n58029 = n58163 & n58164;
  assign n54159 = n58169 ^ n58170;
  assign n58175 = n58185 & n58186;
  assign n57995 = ~n56710;
  assign n58091 = n58131 & n58122;
  assign n58101 = ~n58132;
  assign n58115 = n58135 ^ n58136;
  assign n58137 = n58135 & n58150;
  assign n58129 = n58151 & n58152;
  assign n58143 = ~n58135;
  assign n58145 = n54159 & n58153;
  assign n58033 = ~n58029;
  assign n54186 = ~n54159;
  assign n58165 = ~n58175;
  assign n58080 = n58114 ^ n58115;
  assign n58102 = n58129 ^ n58130;
  assign n58118 = ~n58129;
  assign n58126 = ~n58137;
  assign n58133 = n58143 & n58136;
  assign n56901 = ~n58145;
  assign n58138 = n54186 & n56825;
  assign n58139 = n54186 & n55276;
  assign n58142 = n54186 & n56878;
  assign n58146 = n58165 & n58166;
  assign n58092 = n212 ^ n58102;
  assign n58094 = n58080 & n211;
  assign n58099 = ~n58080;
  assign n58113 = n58117 & n58118;
  assign n58116 = n58126 & n58127;
  assign n58111 = ~n58133;
  assign n58124 = ~n58138;
  assign n56844 = ~n58139;
  assign n56876 = ~n58142;
  assign n58128 = n58146 ^ n58147;
  assign n58148 = ~n58146;
  assign n56620 = n58091 ^ n58092;
  assign n58044 = n58092 & n58091;
  assign n58059 = ~n58094;
  assign n58093 = n58099 & n7845;
  assign n58100 = ~n58113;
  assign n58110 = ~n58116;
  assign n57981 = n58124 & n58125;
  assign n54099 = n58128 ^ n55310;
  assign n58119 = n58128 & n55310;
  assign n58140 = n58148 & n58149;
  assign n57946 = ~n56620;
  assign n58077 = ~n58093;
  assign n58079 = n58100 & n58101;
  assign n58081 = n58110 & n58111;
  assign n58107 = n54099 & n58112;
  assign n58105 = n57981 & n57994;
  assign n58103 = ~n57981;
  assign n54174 = ~n54099;
  assign n56796 = ~n58119;
  assign n58120 = ~n58140;
  assign n58064 = n58079 ^ n58080;
  assign n58071 = n58081 ^ n58082;
  assign n58078 = ~n58079;
  assign n58083 = ~n58081;
  assign n58095 = n58103 & n58104;
  assign n58096 = n54174 & n56638;
  assign n57997 = ~n58105;
  assign n56861 = ~n58107;
  assign n58097 = n54174 & n56836;
  assign n58106 = n58120 & n58121;
  assign n58045 = n211 ^ n58064;
  assign n58039 = n58070 ^ n58071;
  assign n58074 = n58077 & n58078;
  assign n58076 = n58083 & n58084;
  assign n57978 = ~n58095;
  assign n58089 = ~n58096;
  assign n56839 = ~n58097;
  assign n58088 = n58106 ^ n55119;
  assign n58108 = ~n58106;
  assign n56587 = n58044 ^ n58045;
  assign n58052 = n58039 & n7794;
  assign n58056 = ~n58039;
  assign n58057 = ~n58045;
  assign n58058 = ~n58074;
  assign n58072 = ~n58076;
  assign n54056 = n58087 ^ n58088;
  assign n57957 = n58089 & n58090;
  assign n58098 = n58108 & n58109;
  assign n57919 = ~n56587;
  assign n58036 = ~n58052;
  assign n58040 = n58056 & n210;
  assign n58003 = n58057 & n58044;
  assign n58038 = n58058 & n58059;
  assign n58046 = n58072 & n58073;
  assign n58065 = n54056 & n58075;
  assign n57943 = ~n57957;
  assign n54080 = ~n54056;
  assign n58085 = ~n58098;
  assign n58021 = n58038 ^ n58039;
  assign n58016 = ~n58040;
  assign n58030 = n58046 ^ n58047;
  assign n58048 = n58046 & n58047;
  assign n58037 = ~n58038;
  assign n58042 = ~n58046;
  assign n56816 = ~n58065;
  assign n58061 = n54080 & n56812;
  assign n58062 = n54080 & n55192;
  assign n58060 = n54080 & n56546;
  assign n58066 = n58085 & n58086;
  assign n58004 = n210 ^ n58021;
  assign n58001 = n58029 ^ n58030;
  assign n58031 = n58036 & n58037;
  assign n58041 = n58042 & n58043;
  assign n58032 = ~n58048;
  assign n58053 = ~n58060;
  assign n56785 = ~n58061;
  assign n56749 = ~n58062;
  assign n58055 = n58066 ^ n58067;
  assign n58068 = ~n58066;
  assign n56473 = n58003 ^ n58004;
  assign n57954 = n58004 & n58003;
  assign n58005 = n58001 & n7739;
  assign n58006 = ~n58001;
  assign n58015 = ~n58031;
  assign n58022 = n58032 & n58033;
  assign n58014 = ~n58041;
  assign n57887 = n58053 & n58054;
  assign n54020 = n54985 ^ n58055;
  assign n58049 = n58055 & n54985;
  assign n58063 = n58068 & n58069;
  assign n57869 = ~n56473;
  assign n57965 = ~n57954;
  assign n57999 = ~n58005;
  assign n58002 = n58006 & n209;
  assign n58000 = n58015 & n58016;
  assign n58013 = ~n58022;
  assign n58024 = n57887 & n58034;
  assign n58025 = n54020 & n58035;
  assign n54085 = ~n54020;
  assign n58023 = ~n57887;
  assign n56691 = ~n58049;
  assign n58050 = ~n58063;
  assign n57974 = n58000 ^ n58001;
  assign n57980 = ~n58002;
  assign n57998 = ~n58000;
  assign n57993 = n58013 & n58014;
  assign n58019 = n58023 & n57903;
  assign n57905 = ~n58024;
  assign n58020 = n54085 & n56471;
  assign n56760 = ~n58025;
  assign n58017 = n54085 & n56736;
  assign n58026 = n58050 & n58051;
  assign n57955 = n209 ^ n57974;
  assign n57982 = n57993 ^ n57994;
  assign n57985 = n57998 & n57999;
  assign n57996 = ~n57993;
  assign n56734 = ~n58017;
  assign n57886 = ~n58019;
  assign n58007 = ~n58020;
  assign n58010 = n58026 ^ n54992;
  assign n58027 = ~n58026;
  assign n57828 = n57954 ^ n57955;
  assign n57964 = ~n57955;
  assign n57968 = n57981 ^ n57982;
  assign n57979 = ~n57985;
  assign n57986 = n57996 & n57997;
  assign n57863 = n58007 & n58008;
  assign n53980 = n58009 ^ n58010;
  assign n58018 = n58027 & n58028;
  assign n57920 = n57964 & n57965;
  assign n57956 = n57968 & n7684;
  assign n57963 = ~n57968;
  assign n57967 = n57979 & n57980;
  assign n57977 = ~n57986;
  assign n57992 = n53980 & n57995;
  assign n57987 = n53980 & n54945;
  assign n57988 = n53980 & n56400;
  assign n57849 = ~n57863;
  assign n54042 = ~n53980;
  assign n58011 = ~n58018;
  assign n57926 = ~n57920;
  assign n57938 = ~n57956;
  assign n57944 = n57963 & n208;
  assign n57931 = n57967 ^ n57968;
  assign n57939 = ~n57967;
  assign n57958 = n57977 & n57978;
  assign n57983 = n54042 & n56710;
  assign n56618 = ~n57987;
  assign n57975 = ~n57988;
  assign n56678 = ~n57992;
  assign n57989 = n58011 & n58012;
  assign n57921 = n208 ^ n57931;
  assign n57932 = n57938 & n57939;
  assign n57923 = ~n57944;
  assign n57933 = n57957 ^ n57958;
  assign n57961 = n57958 & n57934;
  assign n57959 = ~n57958;
  assign n57791 = n57975 & n57976;
  assign n56713 = ~n57983;
  assign n57973 = n57989 ^ n54861;
  assign n57990 = ~n57989;
  assign n57899 = n57920 ^ n57921;
  assign n57860 = n57921 & n57926;
  assign n57922 = ~n57932;
  assign n57882 = n57933 ^ n57934;
  assign n57945 = n57959 & n57960;
  assign n57942 = ~n57961;
  assign n57966 = n57791 & n57969;
  assign n57962 = ~n57791;
  assign n53997 = n57972 ^ n57973;
  assign n57984 = n57990 & n57991;
  assign n53846 = n57899 ^ n55803;
  assign n57894 = ~n57899;
  assign n57901 = n57922 & n57923;
  assign n57917 = n57882 & n7559;
  assign n57918 = ~n57882;
  assign n57935 = n57942 & n57943;
  assign n57925 = ~n57945;
  assign n57948 = n57962 & n57813;
  assign n57949 = n53997 & n54935;
  assign n57950 = n53997 & n56323;
  assign n57815 = ~n57966;
  assign n57947 = n53997 & n56620;
  assign n53944 = ~n53997;
  assign n57970 = ~n57984;
  assign n53849 = ~n53846;
  assign n57893 = n57894 & n57895;
  assign n57803 = n57894 & n55803;
  assign n57881 = n223 ^ n57901;
  assign n57908 = ~n57901;
  assign n57909 = ~n57917;
  assign n57910 = n57918 & n223;
  assign n57924 = ~n57935;
  assign n57940 = n53944 & n57946;
  assign n56614 = ~n57947;
  assign n57794 = ~n57948;
  assign n56561 = ~n57949;
  assign n57936 = ~n57950;
  assign n57951 = n57970 & n57971;
  assign n57873 = n53849 & n56789;
  assign n57861 = n57881 ^ n57882;
  assign n56814 = ~n57893;
  assign n57900 = n57908 & n57909;
  assign n57884 = ~n57910;
  assign n57902 = n57924 & n57925;
  assign n57752 = n57936 & n57937;
  assign n56655 = ~n57940;
  assign n57930 = n57951 ^ n54834;
  assign n57952 = ~n57951;
  assign n57852 = n57860 ^ n57861;
  assign n57816 = n57861 & n57860;
  assign n57858 = ~n57873;
  assign n57883 = ~n57900;
  assign n57888 = n57902 ^ n57903;
  assign n57904 = ~n57902;
  assign n57762 = ~n57752;
  assign n53915 = n57929 ^ n57930;
  assign n57941 = n57952 & n57953;
  assign n57842 = n57852 & n55646;
  assign n57841 = ~n57852;
  assign n57839 = n57858 & n57859;
  assign n57877 = n57883 & n57884;
  assign n57857 = n57887 ^ n57888;
  assign n57896 = n57904 & n57905;
  assign n57912 = n53915 & n56262;
  assign n57913 = n53915 & n54786;
  assign n57911 = n53915 & n57919;
  assign n53959 = ~n53915;
  assign n57927 = ~n57941;
  assign n57822 = n57839 ^ n57840;
  assign n57833 = n57841 & n55784;
  assign n57811 = ~n57842;
  assign n57837 = ~n57839;
  assign n57862 = n57857 & n222;
  assign n57847 = ~n57877;
  assign n57868 = ~n57857;
  assign n57885 = ~n57896;
  assign n56552 = ~n57911;
  assign n57906 = n53959 & n56587;
  assign n57897 = ~n57912;
  assign n56487 = ~n57913;
  assign n57914 = n57927 & n57928;
  assign n55920 = n359 ^ n57822;
  assign n57686 = n57822 & n359;
  assign n57825 = ~n57833;
  assign n57714 = n57837 & n57838;
  assign n57834 = n57847 ^ n57857;
  assign n57827 = ~n57862;
  assign n57853 = n57868 & n7536;
  assign n57864 = n57885 & n57886;
  assign n57694 = n57897 & n57898;
  assign n56589 = ~n57906;
  assign n57892 = n57914 ^ n54719;
  assign n57915 = ~n57914;
  assign n55948 = ~n55920;
  assign n57801 = n57686 & n358;
  assign n57809 = ~n57686;
  assign n57821 = n57825 & n57803;
  assign n57802 = n57825 & n57811;
  assign n57817 = n222 ^ n57834;
  assign n57846 = ~n57853;
  assign n57843 = n57863 ^ n57864;
  assign n57866 = n57864 & n57875;
  assign n57865 = ~n57864;
  assign n57880 = n57694 & n57718;
  assign n57878 = ~n57694;
  assign n53884 = n57891 ^ n57892;
  assign n57907 = n57915 & n57916;
  assign n57666 = ~n57801;
  assign n53796 = n57802 ^ n57803;
  assign n57795 = n57809 & n4928;
  assign n57770 = n57816 ^ n57817;
  assign n57810 = ~n57821;
  assign n57764 = n57817 & n57816;
  assign n57808 = n57843 ^ n57844;
  assign n57835 = n57846 & n57847;
  assign n57854 = n57865 & n57844;
  assign n57848 = ~n57866;
  assign n57876 = n53884 & n56473;
  assign n57870 = n57878 & n57879;
  assign n57720 = ~n57880;
  assign n57874 = n53884 & n56212;
  assign n57871 = n53884 & n54727;
  assign n53890 = ~n53884;
  assign n57889 = ~n57907;
  assign n57785 = n53796 & n55784;
  assign n57784 = n53796 & n56673;
  assign n57698 = ~n57795;
  assign n53801 = ~n53796;
  assign n57789 = n57810 & n57811;
  assign n57797 = n57770 & n55613;
  assign n57796 = ~n57770;
  assign n57824 = n57808 & n221;
  assign n57826 = ~n57835;
  assign n57823 = ~n57808;
  assign n57845 = n57848 & n57849;
  assign n57832 = ~n57854;
  assign n57867 = n53890 & n57869;
  assign n57697 = ~n57870;
  assign n56417 = ~n57871;
  assign n57855 = ~n57874;
  assign n56477 = ~n57876;
  assign n57872 = n57889 & n57890;
  assign n57772 = ~n57784;
  assign n56703 = ~n57785;
  assign n57771 = n57789 ^ n55611;
  assign n57783 = ~n57789;
  assign n57790 = n57796 & n55611;
  assign n57760 = ~n57797;
  assign n57818 = n57823 & n7384;
  assign n57788 = ~n57824;
  assign n57807 = n57826 & n57827;
  assign n57831 = ~n57845;
  assign n57641 = n57855 & n57856;
  assign n56514 = ~n57867;
  assign n57851 = n57872 ^ n54686;
  assign n53756 = n57770 ^ n57771;
  assign n57757 = n57772 & n57773;
  assign n57782 = ~n57790;
  assign n57786 = n57807 ^ n57808;
  assign n57805 = ~n57807;
  assign n57806 = ~n57818;
  assign n57812 = n57831 & n57832;
  assign n57646 = ~n57641;
  assign n53909 = n57850 ^ n57851;
  assign n57742 = n53756 & n55611;
  assign n57741 = n53756 & n56610;
  assign n57748 = n57757 & n57758;
  assign n53778 = ~n53756;
  assign n57755 = ~n57757;
  assign n57774 = n57782 & n57783;
  assign n57769 = n221 ^ n57786;
  assign n57800 = n57805 & n57806;
  assign n57792 = n57812 ^ n57813;
  assign n57814 = ~n57812;
  assign n56437 = n57828 ^ n53909;
  assign n57830 = n53909 & n57836;
  assign n57829 = n53909 & n56353;
  assign n54760 = ~n53909;
  assign n57733 = ~n57741;
  assign n56648 = ~n57742;
  assign n57728 = ~n57748;
  assign n57743 = n57755 & n57756;
  assign n57711 = n57764 ^ n57769;
  assign n57759 = ~n57774;
  assign n57763 = ~n57769;
  assign n57768 = n57791 ^ n57792;
  assign n57787 = ~n57800;
  assign n57804 = n57814 & n57815;
  assign n57819 = ~n57829;
  assign n56385 = ~n57830;
  assign n57672 = n57733 & n57734;
  assign n57736 = n57728 & n57714;
  assign n57722 = ~n57743;
  assign n57744 = n57711 & n55508;
  assign n57749 = n57759 & n57760;
  assign n57747 = ~n57711;
  assign n57725 = n57763 & n57764;
  assign n57776 = n57768 & n220;
  assign n57767 = n57787 & n57788;
  assign n57775 = ~n57768;
  assign n57793 = ~n57804;
  assign n57798 = n57819 & n57820;
  assign n57705 = n57672 & n57692;
  assign n57703 = ~n57672;
  assign n57713 = n57722 & n57728;
  assign n57721 = ~n57736;
  assign n57732 = ~n57744;
  assign n57740 = n57747 & n55502;
  assign n57729 = ~n57749;
  assign n57746 = n57767 ^ n57768;
  assign n57765 = n57775 & n7394;
  assign n57731 = ~n57776;
  assign n57751 = ~n57767;
  assign n57777 = n57793 & n57794;
  assign n57570 = n57798 ^ n57799;
  assign n57702 = n57703 & n57704;
  assign n57689 = ~n57705;
  assign n57687 = n57713 ^ n57714;
  assign n57691 = n57721 & n57722;
  assign n57712 = n57729 ^ n55502;
  assign n57723 = n57732 & n57729;
  assign n57707 = ~n57740;
  assign n57727 = n220 ^ n57746;
  assign n57750 = ~n57765;
  assign n57753 = n57777 ^ n57778;
  assign n57779 = n57777 & n57778;
  assign n57780 = ~n57777;
  assign n57650 = n57686 ^ n57687;
  assign n57673 = n57691 ^ n57692;
  assign n57680 = n57687 & n57698;
  assign n57664 = ~n57702;
  assign n57690 = ~n57691;
  assign n53729 = n57711 ^ n57712;
  assign n57706 = ~n57723;
  assign n57651 = n57725 ^ n57727;
  assign n57724 = ~n57727;
  assign n57745 = n57750 & n57751;
  assign n57716 = n57752 ^ n57753;
  assign n57761 = ~n57779;
  assign n57766 = n57780 & n57781;
  assign n57634 = n358 ^ n57650;
  assign n57637 = n57672 ^ n57673;
  assign n57665 = ~n57680;
  assign n57679 = n57689 & n57690;
  assign n53741 = ~n53729;
  assign n57700 = n57651 & n55382;
  assign n57688 = n57706 & n57707;
  assign n57699 = ~n57651;
  assign n57659 = n57724 & n57725;
  assign n57737 = n57716 & n7342;
  assign n57730 = ~n57745;
  assign n57735 = ~n57716;
  assign n57754 = n57761 & n57762;
  assign n57739 = ~n57766;
  assign n55894 = n57634 ^ n55920;
  assign n57590 = n57634 & n55920;
  assign n57638 = n57637 & n4867;
  assign n57644 = ~n57637;
  assign n57636 = n57665 & n57666;
  assign n57663 = ~n57679;
  assign n57676 = n53741 & n56523;
  assign n57677 = n53741 & n55508;
  assign n57652 = n57688 ^ n55459;
  assign n57683 = ~n57688;
  assign n57693 = n57699 & n55459;
  assign n57682 = ~n57700;
  assign n57715 = n57730 & n57731;
  assign n57726 = n57735 & n219;
  assign n57708 = ~n57737;
  assign n57738 = ~n57754;
  assign n57166 = ~n55894;
  assign n57607 = n57636 ^ n57637;
  assign n57621 = ~n57638;
  assign n57625 = n57644 & n357;
  assign n53705 = n57651 ^ n57652;
  assign n57622 = ~n57636;
  assign n57639 = n57663 & n57664;
  assign n57661 = ~n57676;
  assign n56575 = ~n57677;
  assign n57675 = n57682 & n57683;
  assign n57654 = ~n57693;
  assign n57681 = n57715 ^ n57716;
  assign n57709 = ~n57715;
  assign n57685 = ~n57726;
  assign n57717 = n57738 & n57739;
  assign n57591 = n357 ^ n57607;
  assign n57616 = n57621 & n57622;
  assign n57593 = ~n57625;
  assign n57609 = n57639 ^ n57631;
  assign n57626 = n53705 & n56457;
  assign n57627 = n53705 & n55382;
  assign n53692 = ~n53705;
  assign n57612 = ~n57639;
  assign n57608 = n57661 & n57662;
  assign n57653 = ~n57675;
  assign n57660 = n219 ^ n57681;
  assign n57701 = n57708 & n57709;
  assign n57695 = n57717 ^ n57718;
  assign n57719 = ~n57717;
  assign n55885 = n57590 ^ n57591;
  assign n57529 = n57591 & n57590;
  assign n57572 = n57608 ^ n57609;
  assign n57592 = ~n57616;
  assign n57614 = ~n57626;
  assign n56495 = ~n57627;
  assign n57628 = n57608 & n57640;
  assign n57630 = ~n57608;
  assign n57649 = n57653 & n57654;
  assign n57599 = n57659 ^ n57660;
  assign n57604 = n57660 & n57659;
  assign n57656 = n57694 ^ n57695;
  assign n57684 = ~n57701;
  assign n57710 = n57719 & n57720;
  assign n57139 = ~n55885;
  assign n57571 = n57592 & n57593;
  assign n57582 = n57572 & n356;
  assign n57589 = ~n57572;
  assign n57541 = n57614 & n57615;
  assign n57611 = ~n57628;
  assign n57617 = n57630 & n57631;
  assign n57629 = n57599 & n55312;
  assign n57632 = ~n57599;
  assign n57603 = ~n57649;
  assign n57667 = n57656 & n7252;
  assign n57674 = ~n57656;
  assign n57655 = n57684 & n57685;
  assign n57696 = ~n57710;
  assign n57548 = n57571 ^ n57572;
  assign n57546 = ~n57582;
  assign n57564 = ~n57571;
  assign n57575 = n57589 & n4824;
  assign n57583 = n57541 & n57598;
  assign n57588 = ~n57541;
  assign n57601 = n57611 & n57612;
  assign n57585 = ~n57617;
  assign n57600 = n57603 ^ n55312;
  assign n57581 = ~n57629;
  assign n57618 = n57632 & n55348;
  assign n57633 = n57655 ^ n57656;
  assign n57647 = ~n57667;
  assign n57657 = n57674 & n218;
  assign n57648 = ~n57655;
  assign n57668 = n57696 & n57697;
  assign n57530 = n356 ^ n57548;
  assign n57563 = ~n57575;
  assign n57565 = ~n57583;
  assign n57576 = n57588 & n57560;
  assign n53643 = n57599 ^ n57600;
  assign n57584 = ~n57601;
  assign n57602 = ~n57618;
  assign n57605 = n218 ^ n57633;
  assign n57635 = n57647 & n57648;
  assign n57624 = ~n57657;
  assign n57642 = n57668 ^ n57669;
  assign n57671 = n57668 & n57678;
  assign n57670 = ~n57668;
  assign n55840 = n57529 ^ n57530;
  assign n57531 = ~n57530;
  assign n57551 = n57563 & n57564;
  assign n57544 = ~n57576;
  assign n57567 = n53643 & n56377;
  assign n57574 = n53643 & n55348;
  assign n57559 = n57584 & n57585;
  assign n53646 = ~n53643;
  assign n57594 = n57602 & n57603;
  assign n57540 = n57604 ^ n57605;
  assign n57549 = n57605 & n57604;
  assign n57623 = ~n57635;
  assign n57596 = n57641 ^ n57642;
  assign n57658 = n57670 & n57669;
  assign n57645 = ~n57671;
  assign n57101 = ~n55840;
  assign n57484 = n57531 & n57529;
  assign n57545 = ~n57551;
  assign n57542 = n57559 ^ n57560;
  assign n57552 = ~n57567;
  assign n56408 = ~n57574;
  assign n57566 = ~n57559;
  assign n57577 = n57540 & n55195;
  assign n57580 = ~n57594;
  assign n57579 = ~n57540;
  assign n57555 = ~n57549;
  assign n57610 = n57596 & n217;
  assign n57595 = n57623 & n57624;
  assign n57613 = ~n57596;
  assign n57643 = n57645 & n57646;
  assign n57620 = ~n57658;
  assign n57491 = ~n57484;
  assign n57523 = n57541 ^ n57542;
  assign n57522 = n57545 & n57546;
  assign n57504 = n57552 & n57553;
  assign n57554 = n57565 & n57566;
  assign n57536 = ~n57577;
  assign n57573 = n57579 & n55266;
  assign n57558 = n57580 & n57581;
  assign n57568 = n57595 ^ n57596;
  assign n57587 = ~n57595;
  assign n57562 = ~n57610;
  assign n57606 = n57613 & n7185;
  assign n57619 = ~n57643;
  assign n57498 = n57522 ^ n57523;
  assign n57516 = n57523 & n355;
  assign n57507 = ~n57522;
  assign n57524 = ~n57523;
  assign n57532 = n57504 & n57519;
  assign n57537 = ~n57504;
  assign n57543 = ~n57554;
  assign n57539 = n57558 ^ n55266;
  assign n57557 = ~n57558;
  assign n57550 = n217 ^ n57568;
  assign n57556 = ~n57573;
  assign n57586 = ~n57606;
  assign n57597 = n57619 & n57620;
  assign n57485 = n355 ^ n57498;
  assign n57479 = ~n57516;
  assign n57510 = n57524 & n4762;
  assign n57520 = ~n57532;
  assign n57525 = n57537 & n57538;
  assign n53621 = n57539 ^ n57540;
  assign n57518 = n57543 & n57544;
  assign n57489 = n57549 ^ n57550;
  assign n57534 = n57550 & n57555;
  assign n57547 = n57556 & n57557;
  assign n57578 = n57586 & n57587;
  assign n57569 = n216 ^ n57597;
  assign n55780 = n57484 ^ n57485;
  assign n57432 = n57485 & n57491;
  assign n57506 = ~n57510;
  assign n57513 = n53621 & n55266;
  assign n57505 = n57518 ^ n57519;
  assign n57512 = n53621 & n56297;
  assign n57500 = ~n57525;
  assign n53585 = ~n53621;
  assign n57521 = ~n57518;
  assign n57527 = n57489 & n55140;
  assign n57526 = ~n57489;
  assign n57535 = ~n57547;
  assign n57515 = n57569 ^ n57570;
  assign n57561 = ~n57578;
  assign n57060 = ~n55780;
  assign n57439 = ~n57432;
  assign n57464 = n57504 ^ n57505;
  assign n57495 = n57506 & n57507;
  assign n57501 = ~n57512;
  assign n56331 = ~n57513;
  assign n57511 = n57520 & n57521;
  assign n57517 = n57526 & n55191;
  assign n57494 = ~n57527;
  assign n57528 = n57535 & n57536;
  assign n57533 = n57561 & n57562;
  assign n57477 = n57464 & n4727;
  assign n57478 = ~n57495;
  assign n57487 = ~n57464;
  assign n57468 = n57501 & n57502;
  assign n57499 = ~n57511;
  assign n57508 = ~n57517;
  assign n57509 = ~n57528;
  assign n57514 = n57533 ^ n57534;
  assign n57461 = ~n57477;
  assign n57463 = n57478 & n57479;
  assign n57475 = n57487 & n354;
  assign n57482 = n57468 & n57492;
  assign n57486 = ~n57468;
  assign n57480 = n57499 & n57500;
  assign n57503 = n57508 & n57509;
  assign n57490 = n57509 ^ n55140;
  assign n57449 = n57514 ^ n57515;
  assign n57447 = n57463 ^ n57464;
  assign n57452 = ~n57475;
  assign n57462 = ~n57463;
  assign n57469 = n57480 ^ n57481;
  assign n57472 = ~n57482;
  assign n57476 = n57486 & n57481;
  assign n53555 = n57489 ^ n57490;
  assign n57473 = ~n57480;
  assign n57497 = n57449 & n55046;
  assign n57493 = ~n57503;
  assign n57496 = ~n57449;
  assign n57433 = n354 ^ n57447;
  assign n57460 = n57461 & n57462;
  assign n57430 = n57468 ^ n57469;
  assign n57465 = n57472 & n57473;
  assign n57455 = ~n57476;
  assign n57471 = n53555 & n55191;
  assign n57470 = n53555 & n56216;
  assign n53587 = ~n53555;
  assign n57483 = n57493 & n57494;
  assign n57488 = n57496 & n55099;
  assign n57474 = ~n57497;
  assign n55721 = n57432 ^ n57433;
  assign n57399 = n57433 & n57439;
  assign n57448 = n57430 & n353;
  assign n57453 = ~n57430;
  assign n57451 = ~n57460;
  assign n57454 = ~n57465;
  assign n57458 = ~n57470;
  assign n56256 = ~n57471;
  assign n57467 = ~n57483;
  assign n57457 = ~n57488;
  assign n57022 = ~n55721;
  assign n57401 = ~n57399;
  assign n57414 = ~n57448;
  assign n57429 = n57451 & n57452;
  assign n57443 = n57453 & n4683;
  assign n57436 = n57454 & n57455;
  assign n57421 = n57458 & n57459;
  assign n57450 = n57467 ^ n55046;
  assign n57466 = n57467 & n57474;
  assign n57410 = n57429 ^ n57430;
  assign n57422 = n57436 ^ n57437;
  assign n57434 = ~n57443;
  assign n57435 = ~n57429;
  assign n57426 = ~n57436;
  assign n53520 = n57449 ^ n57450;
  assign n57444 = n57421 & n57437;
  assign n57445 = ~n57421;
  assign n57456 = ~n57466;
  assign n57400 = n353 ^ n57410;
  assign n57397 = n57421 ^ n57422;
  assign n57423 = n57434 & n57435;
  assign n57431 = n53520 & n56136;
  assign n57427 = n53520 & n55046;
  assign n57425 = ~n57444;
  assign n53553 = ~n53520;
  assign n57442 = n57445 & n57446;
  assign n57438 = n57456 & n57457;
  assign n55666 = n57399 ^ n57400;
  assign n57359 = n57400 & n57401;
  assign n57402 = n57397 & n4635;
  assign n57403 = ~n57397;
  assign n57413 = ~n57423;
  assign n57424 = n57425 & n57426;
  assign n56184 = ~n57427;
  assign n57419 = ~n57431;
  assign n57418 = n57438 ^ n54957;
  assign n57412 = ~n57442;
  assign n57440 = ~n57438;
  assign n56976 = ~n55666;
  assign n57361 = ~n57359;
  assign n57386 = ~n57402;
  assign n57391 = n57403 & n352;
  assign n57396 = n57413 & n57414;
  assign n53477 = n57417 ^ n57418;
  assign n57376 = n57419 & n57420;
  assign n57411 = ~n57424;
  assign n57428 = n57440 & n57441;
  assign n57372 = ~n57391;
  assign n57374 = n57396 ^ n57397;
  assign n57387 = ~n57396;
  assign n57405 = n53477 & n54957;
  assign n57404 = n53477 & n56099;
  assign n53516 = ~n53477;
  assign n57384 = ~n57376;
  assign n57392 = n57411 & n57412;
  assign n57415 = ~n57428;
  assign n57360 = n352 ^ n57374;
  assign n57385 = n57386 & n57387;
  assign n57377 = n57392 ^ n57393;
  assign n57388 = ~n57404;
  assign n56124 = ~n57405;
  assign n57394 = n57392 & n57407;
  assign n57398 = ~n57392;
  assign n57406 = n57415 & n57416;
  assign n55606 = n57359 ^ n57360;
  assign n57318 = n57360 & n57361;
  assign n57355 = n57376 ^ n57377;
  assign n57371 = ~n57385;
  assign n57332 = n57388 & n57389;
  assign n57383 = ~n57394;
  assign n57390 = n57398 & n57393;
  assign n57380 = n57406 ^ n54897;
  assign n57408 = ~n57406;
  assign n56938 = ~n55606;
  assign n57358 = n57355 & n367;
  assign n57356 = ~n57355;
  assign n57354 = n57371 & n57372;
  assign n57373 = n57332 & n57375;
  assign n57370 = ~n57332;
  assign n53472 = n57379 ^ n57380;
  assign n57378 = n57383 & n57384;
  assign n57365 = ~n57390;
  assign n57395 = n57408 & n57409;
  assign n57337 = n57354 ^ n57355;
  assign n57353 = n57356 & n4592;
  assign n57323 = ~n57358;
  assign n57342 = ~n57354;
  assign n57362 = n57370 & n57346;
  assign n57363 = n53472 & n56041;
  assign n57369 = n53472 & n54897;
  assign n57343 = ~n57373;
  assign n57364 = ~n57378;
  assign n53437 = ~n53472;
  assign n57381 = ~n57395;
  assign n57321 = n367 ^ n57337;
  assign n57341 = ~n57353;
  assign n57326 = ~n57362;
  assign n57351 = ~n57363;
  assign n57345 = n57364 & n57365;
  assign n56068 = ~n57369;
  assign n57366 = n57381 & n57382;
  assign n55524 = n57318 ^ n57321;
  assign n57317 = ~n57321;
  assign n57335 = n57341 & n57342;
  assign n57333 = n57345 ^ n57346;
  assign n57299 = n57351 & n57352;
  assign n57344 = ~n57345;
  assign n57350 = n57366 ^ n54777;
  assign n57367 = ~n57366;
  assign n56906 = ~n55524;
  assign n57269 = n57317 & n57318;
  assign n57304 = n57332 ^ n57333;
  assign n57322 = ~n57335;
  assign n57336 = n57299 & n57339;
  assign n57340 = n57343 & n57344;
  assign n57338 = ~n57299;
  assign n53395 = n57349 ^ n57350;
  assign n57357 = n57367 & n57368;
  assign n57284 = ~n57269;
  assign n57307 = n57304 & n366;
  assign n57303 = n57322 & n57323;
  assign n57316 = ~n57304;
  assign n57310 = ~n57336;
  assign n57328 = n53395 & n56000;
  assign n57334 = n53395 & n54828;
  assign n57327 = n57338 & n57309;
  assign n53431 = ~n53395;
  assign n57325 = ~n57340;
  assign n57347 = ~n57357;
  assign n57289 = n57303 ^ n57304;
  assign n57274 = ~n57307;
  assign n57305 = n57316 & n4556;
  assign n57298 = ~n57303;
  assign n57308 = n57325 & n57326;
  assign n57302 = ~n57327;
  assign n57319 = ~n57328;
  assign n56014 = ~n57334;
  assign n57329 = n57347 & n57348;
  assign n57270 = n366 ^ n57289;
  assign n57297 = ~n57305;
  assign n57300 = n57308 ^ n57309;
  assign n57253 = n57319 & n57320;
  assign n57311 = ~n57308;
  assign n57313 = n57329 ^ n54708;
  assign n57330 = ~n57329;
  assign n55447 = n57269 ^ n57270;
  assign n57228 = n57270 & n57284;
  assign n57290 = n57297 & n57298;
  assign n57256 = n57299 ^ n57300;
  assign n57268 = ~n57253;
  assign n57306 = n57310 & n57311;
  assign n53386 = n57312 ^ n57313;
  assign n57324 = n57330 & n57331;
  assign n56859 = ~n55447;
  assign n57227 = ~n57228;
  assign n57280 = n57256 & n365;
  assign n57283 = ~n57256;
  assign n57273 = ~n57290;
  assign n57293 = n53386 & n54728;
  assign n57292 = n53386 & n55967;
  assign n57301 = ~n57306;
  assign n53347 = ~n53386;
  assign n57314 = ~n57324;
  assign n57255 = n57273 & n57274;
  assign n57243 = ~n57280;
  assign n57271 = n57283 & n4506;
  assign n57287 = ~n57292;
  assign n55981 = ~n57293;
  assign n57285 = n57301 & n57302;
  assign n57294 = n57314 & n57315;
  assign n57244 = n57255 ^ n57256;
  assign n57252 = ~n57255;
  assign n57251 = ~n57271;
  assign n57254 = n57285 ^ n57286;
  assign n57275 = n57285 & n57286;
  assign n57213 = n57287 & n57288;
  assign n57276 = ~n57285;
  assign n57281 = n57294 ^ n54631;
  assign n57295 = ~n57294;
  assign n57229 = n365 ^ n57244;
  assign n57250 = n57251 & n57252;
  assign n57220 = n57253 ^ n57254;
  assign n57266 = n57213 & n57231;
  assign n57264 = ~n57213;
  assign n57267 = ~n57275;
  assign n57272 = n57276 & n57277;
  assign n53308 = n57281 ^ n57282;
  assign n57291 = n57295 & n57296;
  assign n56827 = n57228 ^ n57229;
  assign n57226 = ~n57229;
  assign n57236 = n57220 & n4471;
  assign n57242 = ~n57250;
  assign n57237 = ~n57220;
  assign n57257 = n57264 & n57265;
  assign n57258 = n53308 & n55924;
  assign n57259 = n53308 & n54631;
  assign n57233 = ~n57266;
  assign n57263 = n57267 & n57268;
  assign n53350 = ~n53308;
  assign n57246 = ~n57272;
  assign n57278 = ~n57291;
  assign n56817 = ~n56827;
  assign n57192 = n57226 & n57227;
  assign n57224 = ~n57236;
  assign n57235 = n57237 & n364;
  assign n57219 = n57242 & n57243;
  assign n57212 = ~n57257;
  assign n57247 = ~n57258;
  assign n55940 = ~n57259;
  assign n57245 = ~n57263;
  assign n57262 = n57278 & n57279;
  assign n57184 = ~n57192;
  assign n57204 = n57219 ^ n57220;
  assign n57225 = ~n57219;
  assign n57209 = ~n57235;
  assign n57230 = n57245 & n57246;
  assign n57168 = n57247 & n57248;
  assign n57241 = n57262 ^ n54582;
  assign n57260 = ~n57262;
  assign n57193 = n364 ^ n57204;
  assign n57215 = n57224 & n57225;
  assign n57214 = n57230 ^ n57231;
  assign n57232 = ~n57230;
  assign n57182 = ~n57168;
  assign n53260 = n57240 ^ n57241;
  assign n57249 = n57260 & n57261;
  assign n55324 = n57192 ^ n57193;
  assign n57183 = ~n57193;
  assign n57191 = n57213 ^ n57214;
  assign n57208 = ~n57215;
  assign n57223 = n57232 & n57233;
  assign n53290 = ~n53260;
  assign n57238 = ~n57249;
  assign n56777 = ~n55324;
  assign n57146 = n57183 & n57184;
  assign n57194 = n57191 & n4427;
  assign n57195 = ~n57191;
  assign n57190 = n57208 & n57209;
  assign n57216 = n53290 & n55870;
  assign n57218 = n53290 & n54545;
  assign n57211 = ~n57223;
  assign n57234 = n57238 & n57239;
  assign n57165 = n57190 ^ n57191;
  assign n57176 = ~n57194;
  assign n57185 = n57195 & n363;
  assign n57177 = ~n57190;
  assign n57196 = n57211 & n57212;
  assign n57205 = ~n57216;
  assign n55891 = ~n57218;
  assign n57222 = n57234 & n54530;
  assign n57221 = ~n57234;
  assign n57147 = n363 ^ n57165;
  assign n57175 = n57176 & n57177;
  assign n57164 = ~n57185;
  assign n57169 = n57196 ^ n57197;
  assign n57200 = n57196 & n57197;
  assign n57201 = ~n57196;
  assign n57123 = n57205 & n57206;
  assign n57217 = n57221 & n54496;
  assign n57210 = ~n57222;
  assign n55209 = n57146 ^ n57147;
  assign n57148 = ~n57147;
  assign n57145 = n57168 ^ n57169;
  assign n57163 = ~n57175;
  assign n57181 = ~n57200;
  assign n57188 = n57123 & n57136;
  assign n57189 = n57201 & n57202;
  assign n57186 = ~n57123;
  assign n57207 = n57210 & n57179;
  assign n57199 = ~n57217;
  assign n56707 = ~n55209;
  assign n57095 = n57148 & n57146;
  assign n57151 = n57145 & n4376;
  assign n57144 = n57163 & n57164;
  assign n57152 = ~n57145;
  assign n57170 = n57181 & n57182;
  assign n57178 = n57186 & n57187;
  assign n57138 = ~n57188;
  assign n57162 = ~n57189;
  assign n57198 = ~n57207;
  assign n57203 = n57199 & n57210;
  assign n57108 = ~n57095;
  assign n57122 = n57144 ^ n57145;
  assign n57142 = ~n57144;
  assign n57143 = ~n57151;
  assign n57150 = n57152 & n362;
  assign n57161 = ~n57170;
  assign n57117 = ~n57178;
  assign n57171 = n57198 & n57199;
  assign n57180 = ~n57203;
  assign n57096 = n362 ^ n57122;
  assign n57127 = n57142 & n57143;
  assign n57121 = ~n57150;
  assign n57135 = n57161 & n57162;
  assign n57157 = n57171 ^ n57172;
  assign n53217 = n57179 ^ n57180;
  assign n57173 = ~n57171;
  assign n55123 = n57095 ^ n57096;
  assign n57063 = n57096 & n57108;
  assign n57120 = ~n57127;
  assign n57124 = n57135 ^ n57136;
  assign n53240 = n57157 ^ n54510;
  assign n57137 = ~n57135;
  assign n57160 = n53217 & n57166;
  assign n57159 = ~n57157;
  assign n53252 = ~n53217;
  assign n57167 = n57173 & n57174;
  assign n56653 = ~n55123;
  assign n57062 = ~n57063;
  assign n57097 = n57120 & n57121;
  assign n57098 = n57123 ^ n57124;
  assign n57128 = n57137 & n57138;
  assign n57129 = n53240 & n57139;
  assign n57130 = n53240 & n55754;
  assign n53155 = ~n53240;
  assign n57149 = n57159 & n54449;
  assign n55911 = ~n57160;
  assign n57153 = n53252 & n55894;
  assign n57154 = n53252 & n54530;
  assign n57158 = n53252 & n55818;
  assign n57155 = ~n57167;
  assign n57078 = n57097 ^ n57098;
  assign n57107 = n57098 & n4334;
  assign n57086 = ~n57097;
  assign n57099 = ~n57098;
  assign n57116 = ~n57128;
  assign n55883 = ~n57129;
  assign n57125 = n53155 & n55885;
  assign n57118 = ~n57130;
  assign n55829 = ~n57149;
  assign n55896 = ~n57153;
  assign n55867 = ~n57154;
  assign n57133 = n57155 & n57156;
  assign n57140 = ~n57158;
  assign n57064 = n361 ^ n57078;
  assign n57094 = n57099 & n361;
  assign n57085 = ~n57107;
  assign n57104 = n57116 & n57117;
  assign n57041 = n57118 & n57119;
  assign n55859 = ~n57125;
  assign n57112 = n57133 ^ n57134;
  assign n57075 = n57140 & n57141;
  assign n57131 = ~n57133;
  assign n55034 = n57063 ^ n57064;
  assign n57061 = ~n57064;
  assign n57074 = n57085 & n57086;
  assign n57067 = ~n57094;
  assign n57076 = n57104 ^ n57105;
  assign n57103 = n57041 & n57110;
  assign n57102 = n57104 & n57111;
  assign n57100 = ~n57041;
  assign n57106 = ~n57104;
  assign n53117 = n57112 ^ n54433;
  assign n57113 = ~n57112;
  assign n57126 = n57131 & n57132;
  assign n57082 = ~n57075;
  assign n56597 = ~n55034;
  assign n57004 = n57061 & n57062;
  assign n57066 = ~n57074;
  assign n57047 = n57075 ^ n57076;
  assign n57087 = n57100 & n57028;
  assign n57089 = n53117 & n57101;
  assign n57081 = ~n57102;
  assign n57026 = ~n57103;
  assign n57090 = n53117 & n55758;
  assign n57088 = n57106 & n57105;
  assign n53176 = ~n53117;
  assign n57109 = n57113 & n54433;
  assign n57114 = ~n57126;
  assign n57014 = ~n57004;
  assign n57046 = n57066 & n57067;
  assign n57057 = n57047 & n360;
  assign n57056 = ~n57047;
  assign n57077 = n57081 & n57082;
  assign n57048 = ~n57087;
  assign n57069 = ~n57088;
  assign n55821 = ~n57089;
  assign n57079 = ~n57090;
  assign n57083 = n53176 & n55840;
  assign n55786 = ~n57109;
  assign n57091 = n57114 & n57115;
  assign n57029 = n57046 ^ n57047;
  assign n57038 = ~n57046;
  assign n57050 = n57056 & n4295;
  assign n57024 = ~n57057;
  assign n57068 = ~n57077;
  assign n57007 = n57079 & n57080;
  assign n55843 = ~n57083;
  assign n57073 = n57091 ^ n54370;
  assign n57092 = ~n57091;
  assign n57005 = n360 ^ n57029;
  assign n57039 = ~n57050;
  assign n57040 = n57068 & n57069;
  assign n57065 = n57007 & n56994;
  assign n57058 = ~n57007;
  assign n53100 = n57072 ^ n57073;
  assign n57084 = n57092 & n57093;
  assign n54949 = n57004 ^ n57005;
  assign n57013 = ~n57005;
  assign n57030 = n57038 & n57039;
  assign n57027 = n57040 ^ n57041;
  assign n57049 = ~n57040;
  assign n57051 = n57058 & n57059;
  assign n57052 = n53100 & n57060;
  assign n57009 = ~n57065;
  assign n53102 = ~n53100;
  assign n57070 = ~n57084;
  assign n56519 = ~n54949;
  assign n56961 = n57013 & n57014;
  assign n56984 = n57027 ^ n57028;
  assign n57023 = ~n57030;
  assign n57037 = n57048 & n57049;
  assign n56990 = ~n57051;
  assign n55801 = ~n57052;
  assign n57043 = n53102 & n55780;
  assign n57044 = n53102 & n54370;
  assign n57042 = n53102 & n55665;
  assign n57053 = n57070 & n57071;
  assign n57012 = n56984 & n375;
  assign n56999 = n57023 & n57024;
  assign n57015 = ~n56984;
  assign n57025 = ~n57037;
  assign n57035 = ~n57042;
  assign n55773 = ~n57043;
  assign n55730 = ~n57044;
  assign n57032 = n57053 ^ n54327;
  assign n57054 = ~n57053;
  assign n56983 = n375 ^ n56999;
  assign n56965 = ~n57012;
  assign n57003 = n57015 & n4257;
  assign n56992 = ~n56999;
  assign n57006 = n57025 & n57026;
  assign n53038 = n57031 ^ n57032;
  assign n56946 = n57035 & n57036;
  assign n57045 = n57054 & n57055;
  assign n56962 = n56983 ^ n56984;
  assign n56991 = ~n57003;
  assign n56993 = n57006 ^ n57007;
  assign n57008 = ~n57006;
  assign n57019 = n53038 & n57022;
  assign n57016 = n53038 & n55601;
  assign n57017 = n53038 & n54373;
  assign n56956 = ~n56946;
  assign n53098 = ~n53038;
  assign n57033 = ~n57045;
  assign n54864 = n56961 ^ n56962;
  assign n56963 = ~n56962;
  assign n56985 = n56991 & n56992;
  assign n56945 = n56993 ^ n56994;
  assign n57000 = n57008 & n57009;
  assign n57001 = ~n57016;
  assign n57010 = n53098 & n55721;
  assign n55679 = ~n57017;
  assign n55720 = ~n57019;
  assign n57018 = n57033 & n57034;
  assign n56453 = ~n54864;
  assign n56907 = n56963 & n56961;
  assign n56966 = n56945 & n4218;
  assign n56964 = ~n56985;
  assign n56974 = ~n56945;
  assign n56989 = ~n57000;
  assign n56892 = n57001 & n57002;
  assign n55751 = ~n57010;
  assign n56997 = n57018 ^ n54290;
  assign n57020 = ~n57018;
  assign n56910 = ~n56907;
  assign n56944 = n56964 & n56965;
  assign n56949 = ~n56966;
  assign n56957 = n56974 & n374;
  assign n56986 = n56892 & n56917;
  assign n56967 = n56989 & n56990;
  assign n56987 = ~n56892;
  assign n52999 = n56997 ^ n56998;
  assign n57011 = n57020 & n57021;
  assign n56935 = n56944 ^ n56945;
  assign n56934 = ~n56957;
  assign n56950 = ~n56944;
  assign n56947 = n56967 ^ n56968;
  assign n56971 = n56967 & n56968;
  assign n56969 = ~n56967;
  assign n56919 = ~n56986;
  assign n56978 = n52999 & n55666;
  assign n56975 = n56987 & n56988;
  assign n56979 = n52999 & n54290;
  assign n56977 = n52999 & n55561;
  assign n53057 = ~n52999;
  assign n56995 = ~n57011;
  assign n56908 = n374 ^ n56935;
  assign n56912 = n56946 ^ n56947;
  assign n56943 = n56949 & n56950;
  assign n56960 = n56969 & n56970;
  assign n56955 = ~n56971;
  assign n56903 = ~n56975;
  assign n56972 = n53057 & n56976;
  assign n56958 = ~n56977;
  assign n55669 = ~n56978;
  assign n55605 = ~n56979;
  assign n56982 = n56995 & n56996;
  assign n54787 = n56907 ^ n56908;
  assign n56909 = ~n56908;
  assign n56927 = n56912 & n4169;
  assign n56933 = ~n56943;
  assign n56932 = ~n56912;
  assign n56948 = n56955 & n56956;
  assign n56852 = n56958 & n56959;
  assign n56937 = ~n56960;
  assign n55694 = ~n56972;
  assign n56952 = n56982 ^ n54259;
  assign n56980 = ~n56982;
  assign n56868 = n56909 & n56910;
  assign n56914 = ~n56927;
  assign n56926 = n56932 & n373;
  assign n56911 = n56933 & n56934;
  assign n56936 = ~n56948;
  assign n52957 = n56951 ^ n56952;
  assign n56865 = ~n56852;
  assign n56973 = n56980 & n56981;
  assign n56886 = n56911 ^ n56912;
  assign n56915 = ~n56911;
  assign n56888 = ~n56926;
  assign n56916 = n56936 & n56937;
  assign n56939 = n52957 & n55606;
  assign n53015 = ~n52957;
  assign n56953 = ~n56973;
  assign n56871 = n373 ^ n56886;
  assign n56905 = n56914 & n56915;
  assign n56893 = n56916 ^ n56917;
  assign n56918 = ~n56916;
  assign n56928 = n53015 & n56938;
  assign n55640 = ~n56939;
  assign n56929 = n53015 & n55483;
  assign n56930 = n53015 & n54257;
  assign n56940 = n56953 & n56954;
  assign n56849 = n56868 ^ n56871;
  assign n56867 = ~n56871;
  assign n56863 = n56892 ^ n56893;
  assign n56887 = ~n56905;
  assign n56913 = n56918 & n56919;
  assign n55609 = ~n56928;
  assign n56920 = ~n56929;
  assign n55535 = ~n56930;
  assign n56923 = n56940 ^ n54196;
  assign n56941 = ~n56940;
  assign n52680 = n56849 ^ n53849;
  assign n56741 = n56849 & n53849;
  assign n56850 = n56849 & n53846;
  assign n56830 = n56867 & n56868;
  assign n56872 = n56863 & n4120;
  assign n56883 = n56887 & n56888;
  assign n56877 = ~n56863;
  assign n56902 = ~n56913;
  assign n56799 = n56920 & n56921;
  assign n52971 = n56922 ^ n56923;
  assign n56931 = n56941 & n56942;
  assign n56832 = n52680 & n55803;
  assign n52678 = ~n52680;
  assign n55827 = ~n56850;
  assign n56866 = ~n56872;
  assign n56869 = n56877 & n372;
  assign n56862 = ~n56883;
  assign n56873 = n56902 & n56903;
  assign n56895 = n56799 & n56904;
  assign n56897 = n52971 & n55362;
  assign n56896 = n52971 & n56906;
  assign n56898 = n52971 & n54196;
  assign n52914 = ~n52971;
  assign n56894 = ~n56799;
  assign n56924 = ~n56931;
  assign n56813 = ~n56832;
  assign n56840 = n56862 ^ n56863;
  assign n56851 = n56866 & n56862;
  assign n56842 = ~n56869;
  assign n56853 = n56873 ^ n56874;
  assign n56882 = n56873 & n56874;
  assign n56880 = ~n56873;
  assign n56889 = n56894 & n56823;
  assign n56829 = ~n56895;
  assign n55527 = ~n56896;
  assign n56884 = ~n56897;
  assign n56890 = n52914 & n55524;
  assign n55463 = ~n56898;
  assign n56899 = n56924 & n56925;
  assign n56786 = n56813 & n56814;
  assign n56831 = n372 ^ n56840;
  assign n56841 = ~n56851;
  assign n56819 = n56852 ^ n56853;
  assign n56870 = n56880 & n56881;
  assign n56864 = ~n56882;
  assign n56745 = n56884 & n56885;
  assign n56794 = ~n56889;
  assign n55564 = ~n56890;
  assign n56879 = n56899 ^ n54159;
  assign n56900 = ~n56899;
  assign n56764 = n56786 ^ n56787;
  assign n56788 = ~n56786;
  assign n56802 = n56830 ^ n56831;
  assign n56768 = n56831 & n56830;
  assign n56818 = n56841 & n56842;
  assign n56834 = n56819 & n4067;
  assign n56835 = ~n56819;
  assign n56854 = n56864 & n56865;
  assign n56846 = ~n56870;
  assign n56754 = ~n56745;
  assign n52879 = n56878 ^ n56879;
  assign n56891 = n56900 & n56901;
  assign n54385 = n7 ^ n56764;
  assign n56497 = n56764 & n7;
  assign n56604 = n56788 & n56789;
  assign n56791 = n56802 & n53801;
  assign n56801 = ~n56802;
  assign n56792 = n56818 ^ n56819;
  assign n56821 = ~n56818;
  assign n56820 = ~n56834;
  assign n56833 = n56835 & n371;
  assign n56845 = ~n56854;
  assign n56855 = n52879 & n55447;
  assign n56856 = n52879 & n55339;
  assign n56857 = n52879 & n54159;
  assign n52930 = ~n52879;
  assign n56875 = ~n56891;
  assign n55652 = ~n54385;
  assign n56766 = ~n56791;
  assign n56774 = n371 ^ n56792;
  assign n56782 = n56801 & n53796;
  assign n56805 = n56820 & n56821;
  assign n56798 = ~n56833;
  assign n56822 = n56845 & n56846;
  assign n55449 = ~n56855;
  assign n56843 = ~n56856;
  assign n55385 = ~n56857;
  assign n56848 = n52930 & n56859;
  assign n56858 = n56875 & n56876;
  assign n56692 = n56768 ^ n56774;
  assign n56765 = n56766 & n56741;
  assign n56752 = ~n56782;
  assign n56767 = ~n56774;
  assign n56797 = ~n56805;
  assign n56800 = n56822 ^ n56823;
  assign n56828 = ~n56822;
  assign n56667 = n56843 & n56844;
  assign n55489 = ~n56848;
  assign n56837 = n56858 ^ n54099;
  assign n56860 = ~n56858;
  assign n56739 = n56692 & n53756;
  assign n56738 = ~n56692;
  assign n56751 = ~n56765;
  assign n56740 = n56766 & n56752;
  assign n56719 = n56767 & n56768;
  assign n56772 = n56797 & n56798;
  assign n56773 = n56799 ^ n56800;
  assign n56806 = n56828 & n56829;
  assign n56826 = n56667 & n56697;
  assign n52835 = n56836 ^ n56837;
  assign n56824 = ~n56667;
  assign n56847 = n56860 & n56861;
  assign n56732 = n56738 & n53778;
  assign n56695 = ~n56739;
  assign n52585 = n56740 ^ n56741;
  assign n56742 = n56751 & n56752;
  assign n56728 = ~n56719;
  assign n56750 = n56772 ^ n56773;
  assign n56769 = n56773 & n370;
  assign n56744 = ~n56772;
  assign n56779 = ~n56773;
  assign n56793 = ~n56806;
  assign n56807 = n56824 & n56825;
  assign n56699 = ~n56826;
  assign n56809 = n52835 & n56827;
  assign n56808 = n52835 & n55154;
  assign n56810 = n52835 & n54099;
  assign n52847 = ~n52835;
  assign n56838 = ~n56847;
  assign n56716 = n52585 & n53801;
  assign n56715 = n52585 & n55646;
  assign n56725 = ~n56732;
  assign n52594 = ~n52585;
  assign n56717 = ~n56742;
  assign n56720 = n370 ^ n56750;
  assign n56722 = ~n56769;
  assign n56762 = n56779 & n4032;
  assign n56775 = n56793 & n56794;
  assign n56671 = ~n56807;
  assign n56795 = ~n56808;
  assign n55366 = ~n56809;
  assign n55344 = ~n56810;
  assign n56804 = n52847 & n56817;
  assign n56811 = n56838 & n56839;
  assign n56702 = ~n56715;
  assign n55703 = ~n56716;
  assign n56693 = n56717 ^ n53756;
  assign n56623 = n56719 ^ n56720;
  assign n56704 = n56725 & n56717;
  assign n56727 = ~n56720;
  assign n56743 = ~n56762;
  assign n56746 = n56775 ^ n56776;
  assign n56778 = n56775 & n56776;
  assign n56770 = ~n56775;
  assign n56644 = n56795 & n56796;
  assign n55413 = ~n56804;
  assign n56783 = n56811 ^ n56812;
  assign n56815 = ~n56811;
  assign n52534 = n56692 ^ n56693;
  assign n56679 = n56702 & n56703;
  assign n56684 = n56623 & n53741;
  assign n56694 = ~n56704;
  assign n56683 = ~n56623;
  assign n56631 = n56727 & n56728;
  assign n56735 = n56743 & n56744;
  assign n56686 = n56745 ^ n56746;
  assign n56763 = n56770 & n56771;
  assign n56753 = ~n56778;
  assign n56616 = ~n56644;
  assign n52765 = n54056 ^ n56783;
  assign n56780 = n55366 & n55413;
  assign n56790 = ~n56783;
  assign n56803 = n56815 & n56816;
  assign n56664 = n52534 & n53778;
  assign n56656 = n52534 & n55613;
  assign n52522 = ~n52534;
  assign n56669 = n56679 & n56680;
  assign n56672 = ~n56679;
  assign n56675 = n56683 & n53729;
  assign n56626 = ~n56684;
  assign n56662 = n56694 & n56695;
  assign n56630 = ~n56631;
  assign n56724 = n56686 & n3990;
  assign n56726 = ~n56686;
  assign n56721 = ~n56735;
  assign n56747 = n56753 & n56754;
  assign n56730 = ~n56763;
  assign n56761 = n52765 & n55119;
  assign n56757 = n52765 & n56777;
  assign n55406 = ~n56780;
  assign n52850 = ~n52765;
  assign n56781 = n56790 & n54056;
  assign n56784 = ~n56803;
  assign n56647 = ~n56656;
  assign n56624 = n56662 ^ n53729;
  assign n55616 = ~n56664;
  assign n56635 = ~n56669;
  assign n56663 = n56672 & n56673;
  assign n56665 = ~n56662;
  assign n56666 = ~n56675;
  assign n56685 = n56721 & n56722;
  assign n56687 = ~n56724;
  assign n56705 = n56726 & n369;
  assign n56729 = ~n56747;
  assign n55288 = ~n56757;
  assign n56755 = n52850 & n55324;
  assign n56748 = ~n56761;
  assign n55217 = ~n56781;
  assign n56758 = n56784 & n56785;
  assign n52460 = n56623 ^ n56624;
  assign n56533 = n56647 & n56648;
  assign n56642 = n56635 & n56604;
  assign n56622 = ~n56663;
  assign n56649 = n56665 & n56666;
  assign n56657 = n56685 ^ n56686;
  assign n56688 = ~n56685;
  assign n56659 = ~n56705;
  assign n56696 = n56729 & n56730;
  assign n56520 = n56748 & n56749;
  assign n55326 = ~n56755;
  assign n56737 = n56758 ^ n54020;
  assign n56759 = ~n56758;
  assign n56600 = n52460 & n55502;
  assign n56598 = n52460 & n53729;
  assign n52476 = ~n52460;
  assign n56601 = n56533 & n56568;
  assign n56609 = ~n56533;
  assign n56603 = n56622 & n56635;
  assign n56621 = ~n56642;
  assign n56625 = ~n56649;
  assign n56632 = n369 ^ n56657;
  assign n56681 = n56687 & n56688;
  assign n56668 = n56696 ^ n56697;
  assign n56698 = ~n56696;
  assign n56718 = n56520 & n56731;
  assign n56723 = ~n56520;
  assign n52739 = n56736 ^ n56737;
  assign n56756 = n56759 & n56760;
  assign n55552 = ~n56598;
  assign n56574 = ~n56600;
  assign n56592 = ~n56601;
  assign n56579 = n56603 ^ n56604;
  assign n56593 = n56609 & n56610;
  assign n56608 = n56621 & n56622;
  assign n56594 = n56625 & n56626;
  assign n56556 = n56631 ^ n56632;
  assign n56629 = ~n56632;
  assign n56634 = n56667 ^ n56668;
  assign n56658 = ~n56681;
  assign n56689 = n56698 & n56699;
  assign n56714 = n52739 & n55104;
  assign n56548 = ~n56718;
  assign n56708 = n52739 & n55209;
  assign n56711 = n52739 & n54020;
  assign n56706 = n56723 & n56546;
  assign n52807 = ~n52739;
  assign n56733 = ~n56756;
  assign n56479 = n56574 & n56575;
  assign n56566 = n56579 & n6;
  assign n56554 = ~n56593;
  assign n56557 = n56594 ^ n53705;
  assign n56565 = ~n56579;
  assign n56595 = n56556 & n53692;
  assign n56567 = ~n56608;
  assign n56599 = ~n56556;
  assign n56570 = ~n56594;
  assign n56562 = n56629 & n56630;
  assign n56636 = n56634 & n3965;
  assign n56633 = n56658 & n56659;
  assign n56643 = ~n56634;
  assign n56670 = ~n56689;
  assign n56518 = ~n56706;
  assign n56700 = n52807 & n56707;
  assign n55202 = ~n56708;
  assign n55143 = ~n56711;
  assign n56690 = ~n56714;
  assign n56709 = n56733 & n56734;
  assign n56532 = n56479 & n56555;
  assign n52411 = n56556 ^ n56557;
  assign n56539 = ~n56479;
  assign n56558 = n56565 & n21721;
  assign n56499 = ~n56566;
  assign n56534 = n56567 ^ n56568;
  assign n56578 = n56592 & n56567;
  assign n56569 = ~n56595;
  assign n56580 = n56599 & n53705;
  assign n56571 = ~n56562;
  assign n56596 = n56633 ^ n56634;
  assign n56611 = ~n56636;
  assign n56627 = n56643 & n368;
  assign n56612 = ~n56633;
  assign n56645 = n56670 & n56671;
  assign n56446 = n56690 & n56691;
  assign n55253 = ~n56700;
  assign n56682 = n56709 ^ n56710;
  assign n56712 = ~n56709;
  assign n56515 = ~n56532;
  assign n56525 = n52411 & n55459;
  assign n56450 = n56533 ^ n56534;
  assign n56524 = n56539 & n56523;
  assign n56526 = n52411 & n53692;
  assign n52417 = ~n52411;
  assign n56540 = ~n56558;
  assign n56559 = n56569 & n56570;
  assign n56553 = ~n56578;
  assign n56536 = ~n56580;
  assign n56563 = n368 ^ n56596;
  assign n56602 = n56611 & n56612;
  assign n56582 = ~n56627;
  assign n56606 = n56644 ^ n56645;
  assign n56646 = n56645 & n56607;
  assign n56637 = ~n56645;
  assign n56661 = n56446 & n56674;
  assign n56660 = ~n56446;
  assign n52693 = n56682 ^ n54042;
  assign n56676 = n56682 & n54042;
  assign n56701 = n56712 & n56713;
  assign n56491 = n56450 & n5;
  assign n56484 = ~n56524;
  assign n56494 = ~n56525;
  assign n55491 = ~n56526;
  assign n56503 = ~n56450;
  assign n56527 = n56540 & n56497;
  assign n56496 = n56540 & n56499;
  assign n56522 = n56553 & n56554;
  assign n56535 = ~n56559;
  assign n56462 = n56562 ^ n56563;
  assign n56467 = n56563 & n56571;
  assign n56581 = ~n56602;
  assign n56506 = n56606 ^ n56607;
  assign n56628 = n56637 & n56638;
  assign n56615 = ~n56646;
  assign n56650 = n56660 & n56471;
  assign n56482 = ~n56661;
  assign n56651 = n52693 & n55123;
  assign n52755 = ~n52693;
  assign n55029 = ~n56676;
  assign n56677 = ~n56701;
  assign n56424 = ~n56491;
  assign n56409 = n56494 & n56495;
  assign n54316 = n56496 ^ n56497;
  assign n56488 = n56503 & n21670;
  assign n56480 = n56522 ^ n56523;
  assign n56498 = ~n56527;
  assign n56516 = ~n56522;
  assign n56492 = n56535 & n56536;
  assign n56529 = n56462 & n53646;
  assign n56528 = ~n56462;
  assign n56542 = n56581 & n56582;
  assign n56572 = n56506 & n3911;
  assign n56577 = ~n56506;
  assign n56605 = n56615 & n56616;
  assign n56591 = ~n56628;
  assign n56444 = ~n56650;
  assign n56639 = n52755 & n54992;
  assign n55159 = ~n56651;
  assign n56640 = n52755 & n56653;
  assign n56652 = n56677 & n56678;
  assign n56387 = n56479 ^ n56480;
  assign n56458 = n56409 & n56440;
  assign n56456 = ~n56409;
  assign n54348 = ~n54316;
  assign n56461 = ~n56488;
  assign n56463 = n56492 ^ n53643;
  assign n56489 = n56498 & n56499;
  assign n56490 = n56515 & n56516;
  assign n56504 = n56528 & n53643;
  assign n56502 = ~n56529;
  assign n56501 = ~n56492;
  assign n56505 = n383 ^ n56542;
  assign n56543 = ~n56542;
  assign n56544 = ~n56572;
  assign n56564 = n56577 & n383;
  assign n56590 = ~n56605;
  assign n56617 = ~n56639;
  assign n55126 = ~n56640;
  assign n56619 = n56652 ^ n53944;
  assign n56654 = ~n56652;
  assign n56445 = n56387 & n4;
  assign n56438 = ~n56387;
  assign n56448 = n56456 & n56457;
  assign n56442 = ~n56458;
  assign n52355 = n56462 ^ n56463;
  assign n56449 = ~n56489;
  assign n56483 = ~n56490;
  assign n56485 = n56501 & n56502;
  assign n56465 = ~n56504;
  assign n56468 = n56505 ^ n56506;
  assign n56541 = n56543 & n56544;
  assign n56508 = ~n56564;
  assign n56545 = n56590 & n56591;
  assign n56369 = n56617 & n56618;
  assign n52721 = n56619 ^ n56620;
  assign n56641 = n56654 & n56655;
  assign n56418 = n56438 & n21468;
  assign n56422 = n52355 & n55312;
  assign n56420 = n52355 & n53646;
  assign n56361 = ~n56445;
  assign n56412 = ~n56448;
  assign n52362 = ~n52355;
  assign n56413 = n56449 ^ n56450;
  assign n56455 = n56461 & n56449;
  assign n56380 = n56467 ^ n56468;
  assign n56439 = n56483 & n56484;
  assign n56464 = ~n56485;
  assign n56395 = n56468 & n56467;
  assign n56507 = ~n56541;
  assign n56521 = n56545 ^ n56546;
  assign n56547 = ~n56545;
  assign n56585 = n52721 & n56597;
  assign n56583 = n52721 & n53944;
  assign n56584 = n52721 & n54861;
  assign n56383 = ~n56369;
  assign n52640 = ~n52721;
  assign n56613 = ~n56641;
  assign n56378 = n5 ^ n56413;
  assign n56391 = ~n56418;
  assign n55374 = ~n56420;
  assign n56407 = ~n56422;
  assign n56410 = n56439 ^ n56440;
  assign n56423 = ~n56455;
  assign n56428 = n56380 & n53621;
  assign n56441 = ~n56439;
  assign n56451 = n56464 & n56465;
  assign n56427 = ~n56380;
  assign n56414 = ~n56395;
  assign n56474 = n56507 & n56508;
  assign n56475 = n56520 ^ n56521;
  assign n56537 = n56547 & n56548;
  assign n54965 = ~n56583;
  assign n56560 = ~n56584;
  assign n55031 = ~n56585;
  assign n56576 = n52640 & n55034;
  assign n56586 = n56613 & n56614;
  assign n54296 = n56378 ^ n54316;
  assign n56334 = n56378 & n54316;
  assign n56345 = n56407 & n56408;
  assign n56327 = n56409 ^ n56410;
  assign n56386 = n56423 & n56424;
  assign n56421 = n56427 & n53585;
  assign n56375 = ~n56428;
  assign n56419 = n56441 & n56442;
  assign n56393 = ~n56451;
  assign n56429 = n56474 ^ n56475;
  assign n56469 = n56475 & n382;
  assign n56431 = ~n56474;
  assign n56478 = ~n56475;
  assign n56517 = ~n56537;
  assign n56294 = n56560 & n56561;
  assign n55079 = ~n56576;
  assign n56549 = n56586 ^ n56587;
  assign n56588 = ~n56586;
  assign n55494 = ~n54296;
  assign n56342 = ~n56334;
  assign n56362 = n56327 & n21407;
  assign n56366 = n56345 & n56365;
  assign n56357 = n56386 ^ n56387;
  assign n56376 = ~n56345;
  assign n56363 = ~n56327;
  assign n56381 = n56393 ^ n53621;
  assign n56392 = ~n56386;
  assign n56411 = ~n56419;
  assign n56394 = ~n56421;
  assign n56396 = n382 ^ n56429;
  assign n56403 = ~n56469;
  assign n56459 = n56478 & n3849;
  assign n56470 = n56517 & n56518;
  assign n56530 = n56294 & n56538;
  assign n56531 = ~n56294;
  assign n52590 = n53915 ^ n56549;
  assign n56550 = n56549 & n53959;
  assign n56573 = n56588 & n56589;
  assign n56335 = n4 ^ n56357;
  assign n56332 = ~n56362;
  assign n56356 = n56363 & n3;
  assign n56350 = ~n56366;
  assign n56358 = n56376 & n56377;
  assign n52316 = n56380 ^ n56381;
  assign n56379 = n56391 & n56392;
  assign n56390 = n56393 & n56394;
  assign n56315 = n56395 ^ n56396;
  assign n56364 = n56411 & n56412;
  assign n56313 = n56396 & n56414;
  assign n56430 = ~n56459;
  assign n56447 = n56470 ^ n56471;
  assign n56481 = ~n56470;
  assign n56321 = ~n56530;
  assign n56511 = n52590 & n54949;
  assign n56510 = n52590 & n54834;
  assign n56509 = n56531 & n56323;
  assign n52671 = ~n52590;
  assign n54880 = ~n56550;
  assign n56551 = ~n56573;
  assign n54252 = n56334 ^ n56335;
  assign n56274 = n56335 & n56342;
  assign n56299 = ~n56356;
  assign n56325 = ~n56358;
  assign n56348 = n52316 & n55195;
  assign n56349 = n52316 & n53585;
  assign n56346 = n56364 ^ n56365;
  assign n52320 = ~n52316;
  assign n56360 = ~n56379;
  assign n56351 = ~n56364;
  assign n56374 = ~n56390;
  assign n56426 = n56430 & n56431;
  assign n56368 = n56446 ^ n56447;
  assign n56460 = n56481 & n56482;
  assign n56293 = ~n56509;
  assign n56486 = ~n56510;
  assign n54951 = ~n56511;
  assign n56493 = n52671 & n56519;
  assign n56512 = n56551 & n56552;
  assign n55403 = ~n54252;
  assign n56288 = ~n56274;
  assign n56280 = n56345 ^ n56346;
  assign n56330 = ~n56348;
  assign n55283 = ~n56349;
  assign n56336 = n56350 & n56351;
  assign n56326 = n56360 & n56361;
  assign n56337 = n56374 & n56375;
  assign n56398 = n56368 & n381;
  assign n56397 = ~n56368;
  assign n56402 = ~n56426;
  assign n56443 = ~n56460;
  assign n56229 = n56486 & n56487;
  assign n54996 = ~n56493;
  assign n56472 = n56512 ^ n53890;
  assign n56513 = ~n56512;
  assign n56317 = n56280 & n21353;
  assign n56303 = n56326 ^ n56327;
  assign n56305 = ~n56280;
  assign n56269 = n56330 & n56331;
  assign n56324 = ~n56336;
  assign n56316 = n56337 ^ n53555;
  assign n56333 = ~n56326;
  assign n56347 = n56337 & n53587;
  assign n56344 = ~n56337;
  assign n56388 = n56397 & n3787;
  assign n56341 = ~n56398;
  assign n56367 = n56402 & n56403;
  assign n56399 = n56443 & n56444;
  assign n56454 = n56229 & n56466;
  assign n56452 = ~n56229;
  assign n52613 = n56472 ^ n56473;
  assign n56500 = n56513 & n56514;
  assign n56275 = n3 ^ n56303;
  assign n56300 = n56305 & n2;
  assign n56301 = n56269 & n56306;
  assign n52272 = n56315 ^ n56316;
  assign n56276 = ~n56317;
  assign n56302 = ~n56269;
  assign n56296 = n56324 & n56325;
  assign n56319 = n56332 & n56333;
  assign n56328 = n56344 & n53555;
  assign n56318 = ~n56347;
  assign n56343 = n56367 ^ n56368;
  assign n56373 = ~n56388;
  assign n56372 = ~n56367;
  assign n56370 = n56399 ^ n56400;
  assign n56401 = n56399 & n56415;
  assign n56406 = ~n56399;
  assign n56432 = n56452 & n56262;
  assign n56433 = n52613 & n56453;
  assign n56264 = ~n56454;
  assign n56434 = n52613 & n54719;
  assign n56435 = n52613 & n53890;
  assign n52547 = ~n52613;
  assign n56476 = ~n56500;
  assign n55372 = n56274 ^ n56275;
  assign n56214 = n56275 & n56288;
  assign n56270 = n56296 ^ n56297;
  assign n56243 = ~n56300;
  assign n56283 = ~n56301;
  assign n52274 = ~n52272;
  assign n56289 = n56302 & n56297;
  assign n56282 = ~n56296;
  assign n56307 = n56318 & n56315;
  assign n56298 = ~n56319;
  assign n56291 = ~n56328;
  assign n56314 = n381 ^ n56343;
  assign n56309 = n56369 ^ n56370;
  assign n56359 = n56372 & n56373;
  assign n56382 = ~n56401;
  assign n56389 = n56406 & n56400;
  assign n56236 = ~n56432;
  assign n54867 = ~n56433;
  assign n56416 = ~n56434;
  assign n54800 = ~n56435;
  assign n56425 = n52547 & n54864;
  assign n56436 = n56476 & n56477;
  assign n55383 = ~n55372;
  assign n56198 = n56269 ^ n56270;
  assign n56220 = ~n56214;
  assign n56271 = n56282 & n56283;
  assign n56278 = n52274 & n55140;
  assign n56272 = n52274 & n53587;
  assign n56247 = ~n56289;
  assign n56279 = n56298 & n56299;
  assign n56290 = ~n56307;
  assign n56238 = n56313 ^ n56314;
  assign n56249 = n56314 & n56313;
  assign n56339 = n56309 & n380;
  assign n56340 = ~n56359;
  assign n56338 = ~n56309;
  assign n56371 = n56382 & n56383;
  assign n56355 = ~n56389;
  assign n56172 = n56416 & n56417;
  assign n54910 = ~n56425;
  assign n52598 = n56436 ^ n56437;
  assign n56228 = n56198 & n1;
  assign n56231 = ~n56198;
  assign n56246 = ~n56271;
  assign n55223 = ~n56272;
  assign n56255 = ~n56278;
  assign n56245 = n56279 ^ n56280;
  assign n56259 = n56290 & n56291;
  assign n56287 = n56238 & n53553;
  assign n56277 = ~n56279;
  assign n56281 = ~n56238;
  assign n56252 = ~n56249;
  assign n56329 = n56338 & n3736;
  assign n56285 = ~n56339;
  assign n56308 = n56340 & n56341;
  assign n56354 = ~n56371;
  assign n56182 = ~n56172;
  assign n56405 = n52598 & n53909;
  assign n56404 = n52598 & n54686;
  assign n53935 = ~n52598;
  assign n56176 = ~n56228;
  assign n56221 = n56231 & n21237;
  assign n56215 = n2 ^ n56245;
  assign n56244 = n56246 & n56247;
  assign n56185 = n56255 & n56256;
  assign n56239 = n56259 ^ n53520;
  assign n56265 = n56276 & n56277;
  assign n56267 = ~n56259;
  assign n56273 = n56281 & n53520;
  assign n56266 = ~n56287;
  assign n56286 = n56308 ^ n56309;
  assign n56311 = ~n56308;
  assign n56310 = ~n56329;
  assign n56322 = n56354 & n56355;
  assign n56384 = ~n56404;
  assign n54726 = ~n56405;
  assign n54189 = n56214 ^ n56215;
  assign n56213 = ~n56221;
  assign n56219 = ~n56215;
  assign n56227 = n56185 & n56237;
  assign n52226 = n56238 ^ n56239;
  assign n56226 = ~n56185;
  assign n56199 = ~n56244;
  assign n56242 = ~n56265;
  assign n56248 = n56266 & n56267;
  assign n56234 = ~n56273;
  assign n56250 = n380 ^ n56286;
  assign n56304 = n56310 & n56311;
  assign n56295 = n56322 ^ n56323;
  assign n56320 = ~n56322;
  assign n56352 = n56384 & n56385;
  assign n55261 = ~n54189;
  assign n56201 = n52226 & n55099;
  assign n56202 = n52226 & n53553;
  assign n56186 = n56199 ^ n56216;
  assign n56150 = n56219 & n56220;
  assign n52265 = ~n52226;
  assign n56217 = n56226 & n56216;
  assign n56200 = ~n56227;
  assign n56232 = n56242 & n56243;
  assign n56233 = ~n56248;
  assign n56171 = n56249 ^ n56250;
  assign n56251 = ~n56250;
  assign n56258 = n56294 ^ n56295;
  assign n56284 = ~n56304;
  assign n56312 = n56320 & n56321;
  assign n56101 = n56352 ^ n56353;
  assign n56140 = n56185 ^ n56186;
  assign n56157 = ~n56150;
  assign n56195 = n56199 & n56200;
  assign n56183 = ~n56201;
  assign n55131 = ~n56202;
  assign n56169 = ~n56217;
  assign n56197 = ~n56232;
  assign n56203 = n56233 & n56234;
  assign n56222 = n56171 & n53477;
  assign n56225 = ~n56171;
  assign n56190 = n56251 & n56252;
  assign n56268 = n56258 & n379;
  assign n56260 = ~n56258;
  assign n56257 = n56284 & n56285;
  assign n56292 = ~n56312;
  assign n56152 = n56140 & n21168;
  assign n56159 = ~n56140;
  assign n56108 = n56183 & n56184;
  assign n56168 = ~n56195;
  assign n56167 = n56197 ^ n56198;
  assign n56170 = n56203 ^ n53516;
  assign n56196 = n56213 & n56197;
  assign n56188 = ~n56203;
  assign n56165 = ~n56222;
  assign n56218 = n56225 & n53516;
  assign n56224 = n56257 ^ n56258;
  assign n56253 = n56260 & n3634;
  assign n56209 = ~n56268;
  assign n56241 = ~n56257;
  assign n56261 = n56292 & n56293;
  assign n56130 = ~n56152;
  assign n56141 = n56159 & n0;
  assign n56154 = n56108 & n56160;
  assign n56151 = n1 ^ n56167;
  assign n56153 = ~n56108;
  assign n56161 = n56168 & n56169;
  assign n52194 = n56170 ^ n56171;
  assign n56175 = ~n56196;
  assign n56189 = ~n56218;
  assign n56191 = n379 ^ n56224;
  assign n56240 = ~n56253;
  assign n56230 = n56261 ^ n56262;
  assign n56263 = ~n56261;
  assign n56111 = ~n56141;
  assign n54150 = n56150 ^ n56151;
  assign n56148 = n56153 & n56136;
  assign n56134 = ~n56154;
  assign n56143 = n52194 & n53516;
  assign n56088 = n56151 & n56157;
  assign n56142 = n52194 & n54976;
  assign n56135 = ~n56161;
  assign n52197 = ~n52194;
  assign n56139 = n56175 & n56176;
  assign n56187 = n56188 & n56189;
  assign n56112 = n56190 ^ n56191;
  assign n56194 = ~n56191;
  assign n56178 = n56229 ^ n56230;
  assign n56223 = n56240 & n56241;
  assign n56254 = n56263 & n56264;
  assign n55183 = ~n54150;
  assign n56128 = n56134 & n56135;
  assign n56109 = n56135 ^ n56136;
  assign n56116 = n56139 ^ n56140;
  assign n56123 = ~n56142;
  assign n55022 = ~n56143;
  assign n56091 = ~n56088;
  assign n56106 = ~n56148;
  assign n56131 = ~n56139;
  assign n56162 = n56112 & n53437;
  assign n56166 = ~n56112;
  assign n56164 = ~n56187;
  assign n56119 = n56194 & n56190;
  assign n56205 = n56178 & n378;
  assign n56208 = ~n56223;
  assign n56204 = ~n56178;
  assign n56235 = ~n56254;
  assign n56075 = n56108 ^ n56109;
  assign n56089 = n0 ^ n56116;
  assign n56060 = n56123 & n56124;
  assign n56105 = ~n56128;
  assign n56129 = n56130 & n56131;
  assign n56133 = ~n56162;
  assign n56138 = n56164 & n56165;
  assign n56158 = n56166 & n53472;
  assign n56126 = ~n56119;
  assign n56192 = n56204 & n3578;
  assign n56146 = ~n56205;
  assign n56177 = n56208 & n56209;
  assign n56206 = n56235 & n56236;
  assign n55102 = n56088 ^ n56089;
  assign n56087 = n56075 & n21044;
  assign n56086 = ~n56075;
  assign n56090 = ~n56089;
  assign n56079 = n56105 & n56106;
  assign n56104 = n56060 & n56080;
  assign n56098 = ~n56060;
  assign n56110 = ~n56129;
  assign n56113 = n56138 ^ n53472;
  assign n56132 = ~n56138;
  assign n56115 = ~n56158;
  assign n56144 = n56177 ^ n56178;
  assign n56180 = ~n56177;
  assign n56179 = ~n56192;
  assign n56173 = n56206 ^ n56207;
  assign n56210 = n56206 & n56207;
  assign n56211 = ~n56206;
  assign n56061 = n56079 ^ n56080;
  assign n56076 = n56086 & n15;
  assign n56066 = ~n56087;
  assign n54091 = ~n55102;
  assign n56036 = n56090 & n56091;
  assign n56092 = n56098 & n56099;
  assign n56085 = ~n56079;
  assign n56084 = ~n56104;
  assign n56102 = n56110 & n56111;
  assign n52142 = n56112 ^ n56113;
  assign n56125 = n56132 & n56133;
  assign n56120 = n378 ^ n56144;
  assign n56122 = n56172 ^ n56173;
  assign n56163 = n56179 & n56180;
  assign n56181 = ~n56210;
  assign n56193 = n56211 & n56212;
  assign n56020 = n56060 ^ n56061;
  assign n56051 = ~n56076;
  assign n56078 = n56084 & n56085;
  assign n56063 = ~n56092;
  assign n56081 = n52142 & n54872;
  assign n56082 = n52142 & n53437;
  assign n52192 = ~n52142;
  assign n56065 = ~n56102;
  assign n56057 = n56119 ^ n56120;
  assign n56114 = ~n56125;
  assign n56073 = n56120 & n56126;
  assign n56147 = n56122 & n3502;
  assign n56145 = ~n56163;
  assign n56149 = ~n56122;
  assign n56174 = n56181 & n56182;
  assign n56156 = ~n56193;
  assign n56038 = n56020 & n20935;
  assign n56043 = ~n56020;
  assign n56064 = n56065 & n56066;
  assign n56055 = n56065 ^ n56075;
  assign n56062 = ~n56078;
  assign n56067 = ~n56081;
  assign n54938 = ~n56082;
  assign n56097 = n56057 & n53395;
  assign n56093 = ~n56057;
  assign n56103 = n56114 & n56115;
  assign n56077 = ~n56073;
  assign n56121 = n56145 & n56146;
  assign n56118 = ~n56147;
  assign n56137 = n56149 & n377;
  assign n56155 = ~n56174;
  assign n56027 = ~n56038;
  assign n56033 = n56043 & n14;
  assign n56037 = n15 ^ n56055;
  assign n56040 = n56062 & n56063;
  assign n56050 = ~n56064;
  assign n56017 = n56067 & n56068;
  assign n56083 = n56093 & n53431;
  assign n56047 = ~n56097;
  assign n56070 = ~n56103;
  assign n56094 = n56121 ^ n56122;
  assign n56117 = ~n56121;
  assign n56096 = ~n56137;
  assign n56127 = n56155 & n56156;
  assign n56012 = ~n56033;
  assign n54048 = n56036 ^ n56037;
  assign n55986 = n56037 & n56036;
  assign n56018 = n56040 ^ n56041;
  assign n56044 = n56050 & n56051;
  assign n56045 = n56017 & n56058;
  assign n56034 = ~n56040;
  assign n56049 = ~n56017;
  assign n56056 = n56070 ^ n53431;
  assign n56069 = ~n56083;
  assign n56074 = n377 ^ n56094;
  assign n56107 = n56117 & n56118;
  assign n56100 = n376 ^ n56127;
  assign n55997 = n56017 ^ n56018;
  assign n55007 = ~n54048;
  assign n56019 = ~n56044;
  assign n56035 = ~n56045;
  assign n56039 = n56049 & n56041;
  assign n52110 = n56056 ^ n56057;
  assign n56059 = n56069 & n56070;
  assign n56007 = n56073 ^ n56074;
  assign n56052 = n56074 & n56077;
  assign n56072 = n56100 ^ n56101;
  assign n56095 = ~n56107;
  assign n56004 = n55997 & n13;
  assign n56006 = ~n55997;
  assign n56003 = n56019 ^ n56020;
  assign n56023 = n56027 & n56019;
  assign n56032 = n56034 & n56035;
  assign n56016 = ~n56039;
  assign n52152 = ~n52110;
  assign n56054 = n56007 & n53347;
  assign n56046 = ~n56059;
  assign n56048 = ~n56007;
  assign n56071 = n56095 & n56096;
  assign n55987 = n14 ^ n56003;
  assign n55971 = ~n56004;
  assign n55998 = n56006 & n20920;
  assign n56011 = ~n56023;
  assign n56015 = ~n56032;
  assign n56024 = n52152 & n54777;
  assign n56031 = n52152 & n53431;
  assign n56025 = n56046 & n56047;
  assign n56042 = n56048 & n53386;
  assign n56030 = ~n56054;
  assign n56053 = n56071 ^ n56072;
  assign n54907 = n55986 ^ n55987;
  assign n55955 = n55987 & n55986;
  assign n55988 = ~n55998;
  assign n55996 = n56011 & n56012;
  assign n56002 = n56015 & n56016;
  assign n56013 = ~n56024;
  assign n56008 = n56025 ^ n53386;
  assign n54844 = ~n56031;
  assign n56029 = ~n56025;
  assign n56010 = ~n56042;
  assign n55973 = n56052 ^ n56053;
  assign n54010 = ~n54907;
  assign n55972 = n55996 ^ n55997;
  assign n55978 = n56002 ^ n56000;
  assign n55989 = ~n55996;
  assign n55983 = ~n56002;
  assign n52120 = n56007 ^ n56008;
  assign n55977 = n56013 & n56014;
  assign n56021 = n56029 & n56030;
  assign n56026 = n55973 & n53308;
  assign n56028 = ~n55973;
  assign n55956 = n13 ^ n55972;
  assign n55950 = n55977 ^ n55978;
  assign n55982 = n55988 & n55989;
  assign n55990 = n52120 & n54708;
  assign n55991 = n52120 & n53347;
  assign n52072 = ~n52120;
  assign n56001 = n55977 & n56005;
  assign n55999 = ~n55977;
  assign n56009 = ~n56021;
  assign n55976 = ~n56026;
  assign n56022 = n56028 & n53350;
  assign n53965 = n55955 ^ n55956;
  assign n54734 = n55956 & n55955;
  assign n55962 = n55950 & n12;
  assign n55961 = ~n55950;
  assign n55970 = ~n55982;
  assign n55980 = ~n55990;
  assign n54771 = ~n55991;
  assign n55992 = n55999 & n56000;
  assign n55984 = ~n56001;
  assign n55993 = n56009 & n56010;
  assign n55995 = ~n56022;
  assign n54835 = ~n53965;
  assign n55919 = ~n54734;
  assign n55957 = n55961 & n20836;
  assign n55931 = ~n55962;
  assign n55949 = n55970 & n55971;
  assign n55927 = n55980 & n55981;
  assign n55979 = n55983 & n55984;
  assign n55969 = ~n55992;
  assign n55974 = n55993 ^ n53308;
  assign n55994 = ~n55993;
  assign n55934 = n55949 ^ n55950;
  assign n55944 = ~n55957;
  assign n55943 = ~n55949;
  assign n55963 = n55927 & n55947;
  assign n55966 = ~n55927;
  assign n52031 = n55973 ^ n55974;
  assign n55968 = ~n55979;
  assign n55985 = n55994 & n55995;
  assign n54700 = n12 ^ n55934;
  assign n55942 = n55943 & n55944;
  assign n55954 = ~n55963;
  assign n55958 = n55966 & n55967;
  assign n52076 = ~n52031;
  assign n55964 = n55968 & n55969;
  assign n55975 = ~n55985;
  assign n55918 = ~n54700;
  assign n55930 = ~n55942;
  assign n55937 = ~n55958;
  assign n55952 = n52076 & n53350;
  assign n55951 = n52076 & n54625;
  assign n55946 = ~n55964;
  assign n55965 = n55975 & n55976;
  assign n55875 = n55918 & n55919;
  assign n55916 = n55930 & n55931;
  assign n55928 = n55946 ^ n55947;
  assign n55939 = ~n55951;
  assign n54682 = ~n55952;
  assign n55945 = n55954 & n55946;
  assign n55959 = n55965 & n53260;
  assign n55960 = ~n55965;
  assign n55897 = ~n55916;
  assign n55917 = n55927 ^ n55928;
  assign n55904 = n55939 & n55940;
  assign n55936 = ~n55945;
  assign n55941 = ~n55959;
  assign n55953 = n55960 & n53290;
  assign n55901 = n55916 ^ n55917;
  assign n55915 = n55917 & n11;
  assign n55912 = ~n55917;
  assign n55926 = n55904 & n55929;
  assign n55925 = ~n55904;
  assign n55923 = n55936 & n55937;
  assign n55938 = n55941 & n55948;
  assign n55933 = ~n55953;
  assign n55887 = n11 ^ n55901;
  assign n55908 = n55912 & n20775;
  assign n55877 = ~n55915;
  assign n55905 = n55923 ^ n55924;
  assign n55922 = n55925 & n55924;
  assign n55913 = ~n55926;
  assign n55914 = ~n55923;
  assign n55932 = ~n55938;
  assign n55935 = n55933 & n55941;
  assign n55857 = n55875 ^ n55887;
  assign n55874 = ~n55887;
  assign n55849 = n55904 ^ n55905;
  assign n55898 = ~n55908;
  assign n55906 = n55913 & n55914;
  assign n55900 = ~n55922;
  assign n55909 = n55932 & n55933;
  assign n55921 = ~n55935;
  assign n51616 = n52680 ^ n55857;
  assign n55862 = ~n55857;
  assign n55812 = n55874 & n55875;
  assign n55889 = n55849 & n10;
  assign n55888 = ~n55849;
  assign n55892 = n55897 & n55898;
  assign n55899 = ~n55906;
  assign n55893 = n55909 ^ n53217;
  assign n51987 = n55920 ^ n55921;
  assign n55910 = ~n55909;
  assign n51614 = ~n51616;
  assign n55853 = n55862 & n52678;
  assign n55737 = n55862 & n52680;
  assign n55886 = n55888 & n20683;
  assign n55845 = ~n55889;
  assign n55876 = ~n55892;
  assign n51953 = n55893 ^ n55894;
  assign n55878 = n55899 & n55900;
  assign n55902 = n51987 & n54582;
  assign n55903 = n51987 & n53260;
  assign n52050 = ~n51987;
  assign n55907 = n55910 & n55911;
  assign n55833 = n51614 & n53849;
  assign n53860 = ~n55853;
  assign n55873 = n55876 & n55877;
  assign n55864 = n55878 ^ n55879;
  assign n55865 = ~n55886;
  assign n55880 = n51953 & n54496;
  assign n55881 = n51953 & n53217;
  assign n55861 = ~n55878;
  assign n52006 = ~n51953;
  assign n55890 = ~n55902;
  assign n54610 = ~n55903;
  assign n55895 = ~n55907;
  assign n55826 = ~n55833;
  assign n55848 = ~n55873;
  assign n55866 = ~n55880;
  assign n54549 = ~n55881;
  assign n55863 = n55890 & n55891;
  assign n55884 = n55895 & n55896;
  assign n55802 = n55826 & n55827;
  assign n55830 = n55848 ^ n55849;
  assign n55825 = n55863 ^ n55864;
  assign n55854 = n55865 & n55848;
  assign n55793 = n55866 & n55867;
  assign n55855 = n55884 ^ n55885;
  assign n55871 = n55863 & n55879;
  assign n55869 = ~n55863;
  assign n55882 = ~n55884;
  assign n55764 = n55802 ^ n55803;
  assign n55804 = ~n55802;
  assign n55813 = n10 ^ n55830;
  assign n55834 = n55825 & n20607;
  assign n55835 = ~n55825;
  assign n55847 = n55793 & n55850;
  assign n55844 = ~n55854;
  assign n51911 = n55855 ^ n53240;
  assign n55846 = ~n55793;
  assign n55868 = n55869 & n55870;
  assign n55860 = ~n55871;
  assign n55856 = ~n55855;
  assign n55872 = n55882 & n55883;
  assign n53695 = n167 ^ n55764;
  assign n55765 = ~n55764;
  assign n55677 = n55804 & n55803;
  assign n55806 = n55812 ^ n55813;
  assign n55775 = n55813 & n55812;
  assign n55822 = ~n55834;
  assign n55832 = n55835 & n9;
  assign n55824 = n55844 & n55845;
  assign n55836 = n55846 & n55818;
  assign n55814 = ~n55847;
  assign n55841 = n51911 & n54510;
  assign n51921 = ~n51911;
  assign n55852 = n55856 & n53240;
  assign n55851 = n55860 & n55861;
  assign n55838 = ~n55868;
  assign n55858 = ~n55872;
  assign n55533 = ~n53695;
  assign n55589 = n55765 & n167;
  assign n55777 = n55677 & n55646;
  assign n55783 = ~n55677;
  assign n55789 = n55806 & n52585;
  assign n55790 = ~n55806;
  assign n55767 = ~n55775;
  assign n55805 = n55824 ^ n55825;
  assign n55823 = ~n55824;
  assign n55792 = ~n55832;
  assign n55796 = ~n55836;
  assign n55828 = ~n55841;
  assign n55837 = ~n55851;
  assign n54537 = ~n55852;
  assign n55839 = n55858 & n55859;
  assign n55747 = n55589 & n166;
  assign n55746 = ~n55589;
  assign n55644 = ~n55777;
  assign n55763 = n55783 & n55784;
  assign n55735 = ~n55789;
  assign n55787 = n55790 & n52594;
  assign n55776 = n9 ^ n55805;
  assign n55809 = n55822 & n55823;
  assign n55769 = n55828 & n55829;
  assign n55817 = n55837 & n55838;
  assign n55816 = n55839 ^ n55840;
  assign n55842 = ~n55839;
  assign n55731 = n55746 & n17578;
  assign n55578 = ~n55747;
  assign n55671 = ~n55763;
  assign n55755 = n55775 ^ n55776;
  assign n55760 = ~n55787;
  assign n55766 = ~n55776;
  assign n55791 = ~n55809;
  assign n55807 = n55769 & n55810;
  assign n55808 = ~n55769;
  assign n51842 = n53117 ^ n55816;
  assign n55794 = n55817 ^ n55818;
  assign n55819 = n55816 & n53176;
  assign n55815 = ~n55817;
  assign n55831 = n55842 & n55843;
  assign n55592 = ~n55731;
  assign n55739 = n55755 & n52522;
  assign n55683 = ~n55755;
  assign n55756 = n55760 & n55737;
  assign n55736 = n55760 & n55735;
  assign n55715 = n55766 & n55767;
  assign n55778 = n55791 & n55792;
  assign n55779 = n55793 ^ n55794;
  assign n55770 = ~n55807;
  assign n55798 = n51842 & n54420;
  assign n55797 = n55808 & n55754;
  assign n51932 = ~n51842;
  assign n55811 = n55814 & n55815;
  assign n54470 = ~n55819;
  assign n55820 = ~n55831;
  assign n51514 = n55736 ^ n55737;
  assign n55738 = n55683 & n52534;
  assign n55707 = ~n55739;
  assign n55734 = ~n55756;
  assign n55740 = n55778 ^ n55779;
  assign n55774 = n55779 & n8;
  assign n55782 = ~n55779;
  assign n55749 = ~n55778;
  assign n55742 = ~n55797;
  assign n55785 = ~n55798;
  assign n55795 = ~n55811;
  assign n55799 = n55820 & n55821;
  assign n55709 = n51514 & n53796;
  assign n55714 = n51514 & n52594;
  assign n51523 = ~n51514;
  assign n55712 = n55734 & n55735;
  assign n55686 = ~n55738;
  assign n55716 = n8 ^ n55740;
  assign n55725 = ~n55774;
  assign n55761 = n55782 & n20542;
  assign n55697 = n55785 & n55786;
  assign n55768 = n55795 & n55796;
  assign n55781 = n55799 ^ n53100;
  assign n55800 = ~n55799;
  assign n55702 = ~n55709;
  assign n55684 = n55712 ^ n52534;
  assign n53807 = ~n55714;
  assign n55623 = n55715 ^ n55716;
  assign n55626 = n55716 & n55715;
  assign n55708 = ~n55712;
  assign n55748 = ~n55761;
  assign n55759 = n55697 & n55718;
  assign n55753 = n55768 ^ n55769;
  assign n55757 = ~n55697;
  assign n51883 = n55780 ^ n55781;
  assign n55771 = ~n55768;
  assign n55788 = n55800 & n55801;
  assign n51414 = n55683 ^ n55684;
  assign n55676 = n55702 & n55703;
  assign n55688 = n55623 & n52476;
  assign n55706 = n55707 & n55708;
  assign n55687 = ~n55623;
  assign n55629 = ~n55626;
  assign n55732 = n55748 & n55749;
  assign n55673 = n55753 ^ n55754;
  assign n55752 = n55757 & n55758;
  assign n55726 = ~n55759;
  assign n55743 = n51883 & n54411;
  assign n55744 = n51883 & n53100;
  assign n51823 = ~n51883;
  assign n55762 = n55770 & n55771;
  assign n55772 = ~n55788;
  assign n55645 = n55676 ^ n55677;
  assign n51449 = ~n51414;
  assign n55670 = ~n55676;
  assign n55682 = n55687 & n52460;
  assign n55658 = ~n55688;
  assign n55685 = ~n55706;
  assign n55723 = n55673 & n23;
  assign n55728 = ~n55673;
  assign n55724 = ~n55732;
  assign n55729 = ~n55743;
  assign n54432 = ~n55744;
  assign n55701 = ~n55752;
  assign n55741 = ~n55762;
  assign n55745 = n55772 & n55773;
  assign n55590 = n55645 ^ n55646;
  assign n55647 = n51449 & n53756;
  assign n55648 = n51449 & n52522;
  assign n55654 = n55670 & n55671;
  assign n55618 = ~n55682;
  assign n55653 = n55685 & n55686;
  assign n55661 = ~n55723;
  assign n55689 = n55724 & n55725;
  assign n55710 = n55728 & n20485;
  assign n55634 = n55729 & n55730;
  assign n55717 = n55741 & n55742;
  assign n55722 = n55745 ^ n53038;
  assign n55750 = ~n55745;
  assign n55565 = n55589 ^ n55590;
  assign n55591 = ~n55590;
  assign n55615 = ~n55647;
  assign n53786 = ~n55648;
  assign n55624 = n55653 ^ n52460;
  assign n55643 = ~n55654;
  assign n55659 = ~n55653;
  assign n55672 = n23 ^ n55689;
  assign n55695 = ~n55710;
  assign n55704 = n55634 & n55713;
  assign n55696 = ~n55689;
  assign n55698 = n55717 ^ n55718;
  assign n55705 = ~n55634;
  assign n51846 = n55721 ^ n55722;
  assign n55727 = ~n55717;
  assign n55733 = n55750 & n55751;
  assign n55531 = n166 ^ n55565;
  assign n55587 = n55591 & n55592;
  assign n55575 = n55615 & n55616;
  assign n51342 = n55623 ^ n55624;
  assign n55610 = n55643 & n55644;
  assign n55649 = n55658 & n55659;
  assign n55627 = n55672 ^ n55673;
  assign n55680 = n55695 & n55696;
  assign n55631 = n55697 ^ n55698;
  assign n55675 = ~n55704;
  assign n55690 = n55705 & n55665;
  assign n55699 = n51846 & n54327;
  assign n55691 = n51846 & n53098;
  assign n51781 = ~n51846;
  assign n55711 = n55726 & n55727;
  assign n55719 = ~n55733;
  assign n53670 = n55531 ^ n53695;
  assign n55532 = ~n55531;
  assign n55577 = ~n55587;
  assign n55576 = n55610 ^ n55611;
  assign n55581 = n51342 & n53741;
  assign n55582 = n51342 & n52476;
  assign n51384 = ~n51342;
  assign n55593 = n55610 & n55611;
  assign n55580 = ~n55575;
  assign n55612 = ~n55610;
  assign n55544 = n55626 ^ n55627;
  assign n55617 = ~n55649;
  assign n55628 = ~n55627;
  assign n55662 = n55631 & n20442;
  assign n55660 = ~n55680;
  assign n55663 = ~n55631;
  assign n55642 = ~n55690;
  assign n54384 = ~n55691;
  assign n55678 = ~n55699;
  assign n55700 = ~n55711;
  assign n55692 = n55719 & n55720;
  assign n55347 = ~n53670;
  assign n55450 = n55532 & n55533;
  assign n55539 = n55575 ^ n55576;
  assign n55538 = n55577 & n55578;
  assign n55551 = ~n55581;
  assign n53753 = ~n55582;
  assign n55579 = ~n55593;
  assign n55588 = n55612 & n55613;
  assign n55594 = n55544 & n52411;
  assign n55583 = n55617 & n55618;
  assign n55595 = ~n55544;
  assign n55568 = n55628 & n55629;
  assign n55630 = n55660 & n55661;
  assign n55632 = ~n55662;
  assign n55655 = n55663 & n22;
  assign n55570 = n55678 & n55679;
  assign n55667 = n55692 ^ n52999;
  assign n55664 = n55700 & n55701;
  assign n55693 = ~n55692;
  assign n55453 = ~n55450;
  assign n55500 = n55538 ^ n55539;
  assign n55528 = n55539 & n17487;
  assign n55505 = ~n55538;
  assign n55515 = ~n55539;
  assign n55460 = n55551 & n55552;
  assign n55553 = n55579 & n55580;
  assign n55543 = n55583 ^ n52417;
  assign n55542 = ~n55588;
  assign n55530 = ~n55594;
  assign n55584 = n55595 & n52417;
  assign n55554 = ~n55583;
  assign n55574 = ~n55568;
  assign n55596 = n55630 ^ n55631;
  assign n55633 = ~n55630;
  assign n55598 = ~n55655;
  assign n55650 = n55570 & n55656;
  assign n55635 = n55664 ^ n55665;
  assign n55651 = ~n55570;
  assign n51738 = n55666 ^ n55667;
  assign n55674 = ~n55664;
  assign n55681 = n55693 & n55694;
  assign n55451 = n165 ^ n55500;
  assign n55507 = n55515 & n165;
  assign n55504 = ~n55528;
  assign n55467 = ~n55460;
  assign n51292 = n55543 ^ n55544;
  assign n55541 = ~n55553;
  assign n55555 = ~n55584;
  assign n55569 = n22 ^ n55596;
  assign n55625 = n55632 & n55633;
  assign n55557 = n55634 ^ n55635;
  assign n55603 = ~n55650;
  assign n55638 = n55651 & n55601;
  assign n55636 = n51738 & n55652;
  assign n51795 = ~n51738;
  assign n55657 = n55674 & n55675;
  assign n55668 = ~n55681;
  assign n55237 = n55450 ^ n55451;
  assign n55452 = ~n55451;
  assign n55475 = n55504 & n55505;
  assign n55466 = ~n55507;
  assign n55514 = n51292 & n53705;
  assign n55513 = n51292 & n52417;
  assign n51264 = ~n51292;
  assign n55506 = n55541 & n55542;
  assign n55550 = n55554 & n55555;
  assign n55540 = n55568 ^ n55569;
  assign n55573 = ~n55569;
  assign n55599 = n55557 & n21;
  assign n55614 = ~n55557;
  assign n55597 = ~n55625;
  assign n54408 = ~n55636;
  assign n55559 = ~n55638;
  assign n55619 = n51795 & n53057;
  assign n55622 = n51795 & n54329;
  assign n55621 = n51795 & n54385;
  assign n55641 = ~n55657;
  assign n55637 = n55668 & n55669;
  assign n53634 = ~n55237;
  assign n55336 = n55452 & n55453;
  assign n55465 = ~n55475;
  assign n55461 = n55506 ^ n55502;
  assign n55503 = n55506 & n55508;
  assign n53723 = ~n55513;
  assign n55490 = ~n55514;
  assign n55501 = ~n55506;
  assign n55516 = n55540 & n52362;
  assign n55433 = ~n55540;
  assign n55529 = ~n55550;
  assign n55492 = n55573 & n55574;
  assign n55556 = n55597 & n55598;
  assign n55537 = ~n55599;
  assign n55585 = n55614 & n20379;
  assign n54343 = ~n55619;
  assign n54381 = ~n55621;
  assign n55604 = ~n55622;
  assign n55607 = n55637 ^ n52957;
  assign n55600 = n55641 & n55642;
  assign n55639 = ~n55637;
  assign n55425 = n55460 ^ n55461;
  assign n55424 = n55465 & n55466;
  assign n55341 = n55490 & n55491;
  assign n55477 = n55501 & n55502;
  assign n55468 = ~n55503;
  assign n55476 = ~n55516;
  assign n55509 = n55433 & n52355;
  assign n55510 = n55529 & n55530;
  assign n55517 = n55556 ^ n55557;
  assign n55567 = ~n55556;
  assign n55566 = ~n55585;
  assign n55571 = n55600 ^ n55601;
  assign n55480 = n55604 & n55605;
  assign n51695 = n55606 ^ n55607;
  assign n55602 = ~n55600;
  assign n55620 = n55639 & n55640;
  assign n55379 = n55424 ^ n55425;
  assign n55420 = n55425 & n164;
  assign n55387 = ~n55424;
  assign n55426 = ~n55425;
  assign n55436 = n55341 & n55382;
  assign n55464 = n55467 & n55468;
  assign n55458 = ~n55341;
  assign n55429 = ~n55477;
  assign n55438 = ~n55509;
  assign n55469 = ~n55510;
  assign n55493 = n21 ^ n55517;
  assign n55545 = n55566 & n55567;
  assign n55499 = n55570 ^ n55571;
  assign n55572 = n55480 & n55521;
  assign n55560 = ~n55480;
  assign n51767 = ~n51695;
  assign n55586 = n55602 & n55603;
  assign n55608 = ~n55620;
  assign n55337 = n164 ^ n55379;
  assign n55346 = ~n55420;
  assign n55395 = n55426 & n17421;
  assign n55388 = ~n55436;
  assign n55427 = n55458 & n55459;
  assign n55428 = ~n55464;
  assign n55434 = n55469 ^ n52355;
  assign n55474 = n55476 & n55469;
  assign n55376 = n55492 ^ n55493;
  assign n55414 = n55493 & n55492;
  assign n55519 = n55499 & n20;
  assign n55536 = ~n55545;
  assign n55518 = ~n55499;
  assign n55546 = n55560 & n55561;
  assign n55547 = n51767 & n54259;
  assign n55548 = n51767 & n52957;
  assign n55523 = ~n55572;
  assign n55558 = ~n55586;
  assign n55562 = n55608 & n55609;
  assign n55172 = n55336 ^ n55337;
  assign n55224 = n55337 & n55336;
  assign n55386 = ~n55395;
  assign n55354 = ~n55427;
  assign n55421 = n55428 & n55429;
  assign n51192 = n55433 ^ n55434;
  assign n55454 = n55376 & n52320;
  assign n55439 = ~n55376;
  assign n55437 = ~n55474;
  assign n55397 = ~n55414;
  assign n55511 = n55518 & n20341;
  assign n55456 = ~n55519;
  assign n55498 = n55536 & n55537;
  assign n55497 = ~n55546;
  assign n55534 = ~n55547;
  assign n54286 = ~n55548;
  assign n55520 = n55558 & n55559;
  assign n55525 = n55562 ^ n52971;
  assign n55563 = ~n55562;
  assign n53590 = ~n55172;
  assign n55355 = n55386 & n55387;
  assign n55389 = n51192 & n53643;
  assign n55390 = n51192 & n52362;
  assign n55381 = ~n55421;
  assign n51226 = ~n51192;
  assign n55419 = n55437 & n55438;
  assign n55430 = n55439 & n52316;
  assign n55407 = ~n55454;
  assign n55440 = n55498 ^ n55499;
  assign n55478 = ~n55511;
  assign n55479 = ~n55498;
  assign n55481 = n55520 ^ n55521;
  assign n51651 = n55524 ^ n55525;
  assign n55409 = n55534 & n55535;
  assign n55522 = ~n55520;
  assign n55549 = n55563 & n55564;
  assign n55345 = ~n55355;
  assign n55342 = n55381 ^ n55382;
  assign n55380 = n55388 & n55381;
  assign n55373 = ~n55389;
  assign n53660 = ~n55390;
  assign n55375 = n55419 ^ n52320;
  assign n55378 = ~n55430;
  assign n55408 = ~n55419;
  assign n55415 = n20 ^ n55440;
  assign n55470 = n55478 & n55479;
  assign n55399 = n55480 ^ n55481;
  assign n55485 = n55409 & n55443;
  assign n55486 = n51651 & n52914;
  assign n55484 = n51651 & n54232;
  assign n55495 = n51651 & n54296;
  assign n55482 = ~n55409;
  assign n51725 = ~n51651;
  assign n55512 = n55522 & n55523;
  assign n55526 = ~n55549;
  assign n55297 = n55341 ^ n55342;
  assign n55296 = n55345 & n55346;
  assign n55268 = n55373 & n55374;
  assign n51132 = n55375 ^ n55376;
  assign n55353 = ~n55380;
  assign n55394 = n55407 & n55408;
  assign n55292 = n55414 ^ n55415;
  assign n55396 = ~n55415;
  assign n55441 = n55399 & n20295;
  assign n55455 = ~n55470;
  assign n55457 = ~n55399;
  assign n55471 = n55482 & n55483;
  assign n55462 = ~n55484;
  assign n55445 = ~n55485;
  assign n54251 = ~n55486;
  assign n55472 = n51725 & n55494;
  assign n54292 = ~n55495;
  assign n55496 = ~n55512;
  assign n55487 = n55526 & n55527;
  assign n55267 = n55296 ^ n55297;
  assign n55301 = n55297 & n163;
  assign n55298 = ~n55297;
  assign n55265 = ~n55296;
  assign n55313 = n51132 & n55347;
  assign n55335 = n55268 & n55348;
  assign n51151 = ~n51132;
  assign n55333 = ~n55268;
  assign n55311 = n55353 & n55354;
  assign n55356 = n55292 & n52274;
  assign n55370 = ~n55292;
  assign n55377 = ~n55394;
  assign n55327 = n55396 & n55397;
  assign n55416 = ~n55441;
  assign n55398 = n55455 & n55456;
  assign n55431 = n55457 & n19;
  assign n55318 = n55462 & n55463;
  assign n55401 = ~n55471;
  assign n54310 = ~n55472;
  assign n55446 = n55487 ^ n52930;
  assign n55442 = n55496 & n55497;
  assign n55488 = ~n55487;
  assign n55225 = n163 ^ n55267;
  assign n55272 = n55298 & n17333;
  assign n55221 = ~n55301;
  assign n55269 = n55311 ^ n55312;
  assign n53688 = ~n55313;
  assign n55303 = n51151 & n52320;
  assign n55309 = n51151 & n53621;
  assign n55304 = n55333 & n55312;
  assign n55302 = n51151 & n53670;
  assign n55300 = ~n55335;
  assign n55299 = ~n55311;
  assign n55286 = ~n55356;
  assign n55349 = n55370 & n52272;
  assign n55334 = n55377 & n55378;
  assign n55315 = ~n55327;
  assign n55371 = n55398 ^ n55399;
  assign n55417 = ~n55398;
  assign n55358 = ~n55431;
  assign n55423 = n55318 & n55435;
  assign n55410 = n55442 ^ n55443;
  assign n55422 = ~n55318;
  assign n51674 = n55446 ^ n55447;
  assign n55444 = ~n55442;
  assign n55473 = n55488 & n55489;
  assign n53556 = n55224 ^ n55225;
  assign n55094 = n55225 & n55224;
  assign n55178 = n55268 ^ n55269;
  assign n55264 = ~n55272;
  assign n55284 = n55299 & n55300;
  assign n53672 = ~n55302;
  assign n53641 = ~n55303;
  assign n55263 = ~n55304;
  assign n55282 = ~n55309;
  assign n55293 = n55334 ^ n52272;
  assign n55330 = ~n55349;
  assign n55329 = ~n55334;
  assign n55328 = n19 ^ n55371;
  assign n55332 = n55409 ^ n55410;
  assign n55391 = n55416 & n55417;
  assign n55402 = n55422 & n55362;
  assign n55369 = ~n55423;
  assign n55411 = n51674 & n54252;
  assign n55418 = n51674 & n52930;
  assign n55404 = n51674 & n54186;
  assign n51602 = ~n51674;
  assign n55432 = n55444 & n55445;
  assign n55448 = ~n55473;
  assign n55065 = ~n53556;
  assign n55097 = ~n55094;
  assign n55232 = n55178 & n162;
  assign n55260 = n55264 & n55265;
  assign n55233 = ~n55178;
  assign n55163 = n55282 & n55283;
  assign n55262 = ~n55284;
  assign n51073 = n55292 ^ n55293;
  assign n55203 = n55327 ^ n55328;
  assign n55305 = n55329 & n55330;
  assign n55314 = ~n55328;
  assign n55359 = n55332 & n20271;
  assign n55360 = ~n55332;
  assign n55357 = ~n55391;
  assign n55321 = ~n55402;
  assign n55392 = n51602 & n55403;
  assign n55384 = ~n55404;
  assign n54255 = ~n55411;
  assign n54210 = ~n55418;
  assign n55400 = ~n55432;
  assign n55405 = n55448 & n55449;
  assign n55135 = ~n55232;
  assign n55214 = n55233 & n17249;
  assign n55220 = ~n55260;
  assign n55236 = n51073 & n53634;
  assign n55259 = n51073 & n52272;
  assign n55258 = n55262 & n55263;
  assign n55234 = n55163 & n55266;
  assign n55235 = n51073 & n53555;
  assign n51081 = ~n51073;
  assign n55254 = ~n55163;
  assign n55285 = ~n55305;
  assign n55219 = ~n55203;
  assign n55240 = n55314 & n55315;
  assign n55331 = n55357 & n55358;
  assign n55317 = ~n55359;
  assign n55352 = n55360 & n18;
  assign n55245 = n55384 & n55385;
  assign n54277 = ~n55392;
  assign n55361 = n55400 & n55401;
  assign n51547 = n55405 ^ n55406;
  assign n55412 = ~n55405;
  assign n55175 = ~n55214;
  assign n55177 = n55220 & n55221;
  assign n55215 = ~n55234;
  assign n55222 = ~n55235;
  assign n53636 = ~n55236;
  assign n55227 = n51081 & n55237;
  assign n55226 = n55254 & n55195;
  assign n55194 = ~n55258;
  assign n53602 = ~n55259;
  assign n55255 = n55285 & n55286;
  assign n55273 = n55331 ^ n55332;
  assign n55340 = n55245 & n55276;
  assign n55316 = ~n55331;
  assign n55290 = ~n55352;
  assign n55319 = n55361 ^ n55362;
  assign n55338 = ~n55245;
  assign n55363 = n51547 & n55383;
  assign n55364 = n51547 & n54174;
  assign n55367 = n51547 & n52847;
  assign n55368 = ~n55361;
  assign n51552 = ~n51547;
  assign n55393 = n55412 & n55413;
  assign n55136 = n55177 ^ n55178;
  assign n55164 = n55194 ^ n55195;
  assign n55176 = ~n55177;
  assign n55193 = n55215 & n55194;
  assign n55084 = n55222 & n55223;
  assign n55180 = ~n55226;
  assign n53651 = ~n55227;
  assign n55204 = n55255 ^ n52226;
  assign n55239 = n55255 & n52265;
  assign n55238 = ~n55255;
  assign n55241 = n18 ^ n55273;
  assign n55306 = n55316 & n55317;
  assign n55257 = n55318 ^ n55319;
  assign n55322 = n55338 & n55339;
  assign n55278 = ~n55340;
  assign n54213 = ~n55363;
  assign n55343 = ~n55364;
  assign n54198 = ~n55367;
  assign n55350 = n55368 & n55369;
  assign n55351 = n51552 & n55372;
  assign n55365 = ~n55393;
  assign n55095 = n162 ^ n55136;
  assign n55087 = n55163 ^ n55164;
  assign n55171 = n55175 & n55176;
  assign n55181 = n55084 & n55191;
  assign n55179 = ~n55193;
  assign n51000 = n55203 ^ n55204;
  assign n55187 = ~n55084;
  assign n55228 = n55238 & n52226;
  assign n55218 = ~n55239;
  assign n55106 = n55240 ^ n55241;
  assign n55242 = ~n55241;
  assign n55274 = n55257 & n17;
  assign n55289 = ~n55306;
  assign n55291 = ~n55257;
  assign n55248 = ~n55322;
  assign n55200 = n55343 & n55344;
  assign n55320 = ~n55350;
  assign n54235 = ~n55351;
  assign n55323 = n55365 & n55366;
  assign n53527 = n55094 ^ n55095;
  assign n55096 = ~n55095;
  assign n55127 = n55087 & n17182;
  assign n55122 = ~n55087;
  assign n55134 = ~n55171;
  assign n55139 = n55179 & n55180;
  assign n55132 = ~n55181;
  assign n55149 = n51000 & n53520;
  assign n55150 = n51000 & n53590;
  assign n55165 = n51000 & n52265;
  assign n55148 = n55187 & n55140;
  assign n51008 = ~n51000;
  assign n55213 = n55106 & n52194;
  assign n55196 = n55218 & n55219;
  assign n55186 = ~n55228;
  assign n55205 = ~n55106;
  assign n55151 = n55242 & n55240;
  assign n55207 = ~n55274;
  assign n55256 = n55289 & n55290;
  assign n55270 = n55291 & n20212;
  assign n55295 = n55200 & n55310;
  assign n55275 = n55320 & n55321;
  assign n55294 = ~n55200;
  assign n55279 = n55323 ^ n55324;
  assign n55307 = n54235 & n54213;
  assign n55325 = ~n55323;
  assign n54971 = ~n53527;
  assign n55001 = n55096 & n55097;
  assign n55107 = n55122 & n161;
  assign n55093 = ~n55127;
  assign n55086 = n55134 & n55135;
  assign n55085 = n55139 ^ n55140;
  assign n55101 = ~n55148;
  assign n55130 = ~n55149;
  assign n53600 = ~n55150;
  assign n53565 = ~n55165;
  assign n55133 = ~n55139;
  assign n55144 = n51008 & n55172;
  assign n55185 = ~n55196;
  assign n55188 = n55205 & n52197;
  assign n55090 = ~n55213;
  assign n55170 = ~n55151;
  assign n55197 = n55256 ^ n55257;
  assign n55244 = ~n55256;
  assign n55243 = ~n55270;
  assign n55246 = n55275 ^ n55276;
  assign n51418 = n52765 ^ n55279;
  assign n55280 = n55294 & n55154;
  assign n55281 = n55279 & n52850;
  assign n55211 = ~n55295;
  assign n55277 = ~n55275;
  assign n54237 = ~n55307;
  assign n55308 = n55325 & n55326;
  assign n55017 = ~n55001;
  assign n55006 = n55084 ^ n55085;
  assign n55044 = n55086 ^ n55087;
  assign n55055 = ~n55107;
  assign n55092 = ~n55086;
  assign n55003 = n55130 & n55131;
  assign n55111 = n55132 & n55133;
  assign n53610 = ~n55144;
  assign n55141 = n55185 & n55186;
  assign n55138 = ~n55188;
  assign n55152 = n17 ^ n55197;
  assign n55229 = n55243 & n55244;
  assign n55167 = n55245 ^ n55246;
  assign n55249 = n51418 & n55261;
  assign n55250 = n51418 & n54080;
  assign n51582 = ~n51418;
  assign n55271 = n55277 & n55278;
  assign n55174 = ~n55280;
  assign n54137 = ~n55281;
  assign n55287 = ~n55308;
  assign n55002 = n161 ^ n55044;
  assign n55059 = n55006 & n160;
  assign n55053 = ~n55006;
  assign n55083 = n55092 & n55093;
  assign n55088 = n55003 & n55046;
  assign n55100 = ~n55111;
  assign n55098 = ~n55003;
  assign n55105 = n55141 ^ n52197;
  assign n55015 = n55151 ^ n55152;
  assign n55137 = ~n55141;
  assign n55169 = ~n55152;
  assign n55198 = n55167 & n20204;
  assign n55206 = ~n55229;
  assign n55212 = ~n55167;
  assign n54166 = ~n55249;
  assign n55231 = n51582 & n54189;
  assign n55216 = ~n55250;
  assign n55247 = ~n55271;
  assign n55251 = n55287 & n55288;
  assign n53482 = n55001 ^ n55002;
  assign n55016 = ~n55002;
  assign n55041 = n55053 & n17111;
  assign n54970 = ~n55059;
  assign n55054 = ~n55083;
  assign n55058 = ~n55088;
  assign n55082 = n55098 & n55099;
  assign n55045 = n55100 & n55101;
  assign n50940 = n55105 ^ n55106;
  assign n55114 = n55015 & n52142;
  assign n55112 = n55137 & n55138;
  assign n55113 = ~n55015;
  assign n55066 = n55169 & n55170;
  assign n55162 = ~n55198;
  assign n55166 = n55206 & n55207;
  assign n55189 = n55212 & n16;
  assign n55071 = n55216 & n55217;
  assign n54194 = ~n55231;
  assign n55199 = n55247 & n55248;
  assign n55208 = n55251 ^ n52807;
  assign n55252 = ~n55251;
  assign n54891 = ~n53482;
  assign n54919 = n55016 & n55017;
  assign n55008 = ~n55041;
  assign n55004 = n55045 ^ n55046;
  assign n55005 = n55054 & n55055;
  assign n55047 = n50940 & n53477;
  assign n55049 = n50940 & n52197;
  assign n55048 = n50940 & n55065;
  assign n50975 = ~n50940;
  assign n55057 = ~n55045;
  assign n55013 = ~n55082;
  assign n55089 = ~n55112;
  assign n55108 = n55113 & n52192;
  assign n55011 = ~n55114;
  assign n55069 = ~n55066;
  assign n55115 = n55166 ^ n55167;
  assign n55161 = ~n55166;
  assign n55121 = ~n55189;
  assign n55182 = n55071 & n55192;
  assign n55153 = n55199 ^ n55200;
  assign n55184 = ~n55071;
  assign n51518 = n55208 ^ n55209;
  assign n55210 = ~n55199;
  assign n55230 = n55252 & n55253;
  assign n54922 = ~n54919;
  assign n54924 = n55003 ^ n55004;
  assign n54958 = n55005 ^ n55006;
  assign n55009 = ~n55005;
  assign n55021 = ~n55047;
  assign n55023 = n50975 & n53556;
  assign n53563 = ~n55048;
  assign n53530 = ~n55049;
  assign n55043 = n55057 & n55058;
  assign n55056 = n55089 & n55090;
  assign n55051 = ~n55108;
  assign n55067 = n16 ^ n55115;
  assign n55025 = n55153 ^ n55154;
  assign n55145 = n55161 & n55162;
  assign n55129 = ~n55182;
  assign n55156 = n51518 & n52807;
  assign n55168 = n51518 & n54085;
  assign n55160 = n51518 & n55183;
  assign n55155 = n55184 & n55119;
  assign n51389 = ~n51518;
  assign n55190 = n55210 & n55211;
  assign n55201 = ~n55230;
  assign n54920 = n160 ^ n54958;
  assign n54959 = n54924 & n17044;
  assign n54972 = ~n54924;
  assign n54980 = n55008 & n55009;
  assign n54893 = n55021 & n55022;
  assign n53580 = ~n55023;
  assign n55012 = ~n55043;
  assign n55014 = n55056 ^ n52192;
  assign n55050 = ~n55056;
  assign n55052 = n55066 ^ n55067;
  assign n55068 = ~n55067;
  assign n55117 = n55025 & n31;
  assign n55120 = ~n55145;
  assign n55116 = ~n55025;
  assign n55076 = ~n55155;
  assign n54097 = ~n55156;
  assign n54129 = ~n55160;
  assign n55146 = n51389 & n54150;
  assign n55142 = ~n55168;
  assign n55173 = ~n55190;
  assign n55157 = n55201 & n55202;
  assign n53439 = n54919 ^ n54920;
  assign n54921 = ~n54920;
  assign n54925 = ~n54959;
  assign n54939 = n54972 & n175;
  assign n54969 = ~n54980;
  assign n54978 = n54893 & n54957;
  assign n54981 = n55012 & n55013;
  assign n50904 = n55014 ^ n55015;
  assign n54975 = ~n54893;
  assign n55036 = n55050 & n55051;
  assign n55042 = n55052 & n52110;
  assign n54930 = ~n55052;
  assign n54989 = n55068 & n55069;
  assign n55109 = n55116 & n20137;
  assign n55027 = ~n55117;
  assign n55070 = n55120 & n55121;
  assign n55039 = n55142 & n55143;
  assign n54152 = ~n55146;
  assign n55124 = n55157 ^ n52693;
  assign n55118 = n55173 & n55174;
  assign n55158 = ~n55157;
  assign n54798 = ~n53439;
  assign n54840 = n54921 & n54922;
  assign n54886 = ~n54939;
  assign n54923 = n54969 & n54970;
  assign n54960 = n54975 & n54976;
  assign n54966 = n50904 & n53527;
  assign n54952 = ~n54978;
  assign n54961 = n50904 & n53472;
  assign n54962 = n50904 & n52192;
  assign n54953 = ~n54981;
  assign n50911 = ~n50904;
  assign n55018 = n54930 & n52152;
  assign n55010 = ~n55036;
  assign n54968 = ~n55042;
  assign n55024 = n31 ^ n55070;
  assign n55081 = ~n55109;
  assign n55091 = n55039 & n54985;
  assign n55080 = ~n55070;
  assign n55072 = n55118 ^ n55119;
  assign n55103 = ~n55039;
  assign n51310 = n55123 ^ n55124;
  assign n55128 = ~n55118;
  assign n55147 = n55158 & n55159;
  assign n54884 = n54923 ^ n54924;
  assign n54926 = ~n54923;
  assign n54933 = n54952 & n54953;
  assign n54894 = n54953 ^ n54957;
  assign n54896 = ~n54960;
  assign n54937 = ~n54961;
  assign n53491 = ~n54962;
  assign n53524 = ~n54966;
  assign n54940 = n50911 & n54971;
  assign n54963 = n55010 & n55011;
  assign n54929 = ~n55018;
  assign n54990 = n55024 ^ n55025;
  assign n54983 = n55071 ^ n55072;
  assign n55064 = n55080 & n55081;
  assign n55033 = ~n55091;
  assign n55073 = n51310 & n55102;
  assign n55077 = n55103 & n55104;
  assign n51442 = ~n51310;
  assign n55110 = n55128 & n55129;
  assign n55125 = ~n55147;
  assign n54841 = n175 ^ n54884;
  assign n54839 = n54893 ^ n54894;
  assign n54913 = n54925 & n54926;
  assign n54895 = ~n54933;
  assign n54809 = n54937 & n54938;
  assign n53540 = ~n54940;
  assign n54931 = n54963 ^ n52110;
  assign n54967 = ~n54963;
  assign n54878 = n54989 ^ n54990;
  assign n54917 = n54990 & n54989;
  assign n55037 = n54983 & n30;
  assign n55040 = ~n54983;
  assign n55026 = ~n55064;
  assign n55060 = n51442 & n53980;
  assign n54115 = ~n55073;
  assign n55061 = n51442 & n54091;
  assign n55062 = n51442 & n52693;
  assign n54998 = ~n55077;
  assign n55075 = ~n55110;
  assign n55074 = n55125 & n55126;
  assign n53398 = n54840 ^ n54841;
  assign n54757 = n54841 & n54840;
  assign n54851 = n54839 & n174;
  assign n54873 = ~n54839;
  assign n54871 = n54895 & n54896;
  assign n54889 = n54809 & n54897;
  assign n54885 = ~n54913;
  assign n54892 = ~n54809;
  assign n50861 = n54930 ^ n54931;
  assign n54941 = n54967 & n54968;
  assign n54850 = ~n54878;
  assign n54899 = ~n54917;
  assign n54982 = n55026 & n55027;
  assign n54955 = ~n55037;
  assign n55019 = n55040 & n20098;
  assign n55028 = ~n55060;
  assign n54090 = ~n55061;
  assign n54053 = ~n55062;
  assign n55035 = n55074 ^ n52721;
  assign n55038 = n55075 & n55076;
  assign n55078 = ~n55074;
  assign n54705 = ~n53398;
  assign n54775 = ~n54851;
  assign n54810 = n54871 ^ n54872;
  assign n54842 = n54873 & n17004;
  assign n54838 = n54885 & n54886;
  assign n54876 = n50861 & n52110;
  assign n54854 = ~n54889;
  assign n54853 = ~n54871;
  assign n54875 = n50861 & n53395;
  assign n54874 = n50861 & n54891;
  assign n54883 = n54892 & n54872;
  assign n50870 = ~n50861;
  assign n54928 = ~n54941;
  assign n54956 = n54982 ^ n54983;
  assign n54994 = ~n55019;
  assign n54993 = ~n54982;
  assign n54911 = n55028 & n55029;
  assign n51230 = n55034 ^ n55035;
  assign n54984 = n55038 ^ n55039;
  assign n55032 = ~n55038;
  assign n55063 = n55078 & n55079;
  assign n54730 = n54809 ^ n54810;
  assign n54795 = n54838 ^ n54839;
  assign n54821 = ~n54842;
  assign n54848 = n54853 & n54854;
  assign n54822 = ~n54838;
  assign n54852 = n50870 & n53482;
  assign n53485 = ~n54874;
  assign n54843 = ~n54875;
  assign n53446 = ~n54876;
  assign n54830 = ~n54883;
  assign n54877 = n54928 & n54929;
  assign n54918 = n30 ^ n54956;
  assign n54901 = n54984 ^ n54985;
  assign n54977 = n54993 & n54994;
  assign n54986 = n51230 & n53997;
  assign n54987 = n51230 & n55007;
  assign n54999 = n54911 & n54945;
  assign n55000 = n51230 & n52640;
  assign n54991 = ~n54911;
  assign n51379 = ~n51230;
  assign n55020 = n55032 & n55033;
  assign n55030 = ~n55063;
  assign n54758 = n174 ^ n54795;
  assign n54773 = n54730 & n173;
  assign n54789 = ~n54730;
  assign n54805 = n54821 & n54822;
  assign n54755 = n54843 & n54844;
  assign n54829 = ~n54848;
  assign n53499 = ~n54852;
  assign n54831 = n54877 ^ n54878;
  assign n54881 = n54877 & n52072;
  assign n54882 = ~n54877;
  assign n54731 = n54917 ^ n54918;
  assign n54898 = ~n54918;
  assign n54942 = n54901 & n20052;
  assign n54943 = ~n54901;
  assign n54954 = ~n54977;
  assign n54964 = ~n54986;
  assign n54050 = ~n54987;
  assign n54974 = n51379 & n54048;
  assign n54973 = n54991 & n54992;
  assign n54947 = ~n54999;
  assign n54012 = ~n55000;
  assign n54997 = ~n55020;
  assign n54988 = n55030 & n55031;
  assign n53378 = n54757 ^ n54758;
  assign n54724 = ~n54773;
  assign n54762 = n54789 & n16960;
  assign n54759 = ~n54758;
  assign n54774 = ~n54805;
  assign n54802 = n54755 & n54828;
  assign n54776 = n54829 & n54830;
  assign n50819 = n52120 ^ n54831;
  assign n54804 = ~n54755;
  assign n54832 = n54831 & n52072;
  assign n54849 = ~n54881;
  assign n54855 = n54882 & n52120;
  assign n54856 = n54731 & n52076;
  assign n54857 = ~n54731;
  assign n54823 = n54898 & n54899;
  assign n54903 = ~n54942;
  assign n54934 = n54943 & n29;
  assign n54900 = n54954 & n54955;
  assign n54813 = n54964 & n54965;
  assign n54915 = ~n54973;
  assign n54074 = ~n54974;
  assign n54948 = n54988 ^ n52671;
  assign n54944 = n54997 & n54998;
  assign n54995 = ~n54988;
  assign n54641 = ~n53378;
  assign n54661 = n54759 & n54757;
  assign n54751 = ~n54762;
  assign n54772 = n54774 & n54775;
  assign n54756 = n54776 ^ n54777;
  assign n54778 = ~n54776;
  assign n54779 = ~n54802;
  assign n54797 = n50819 & n53386;
  assign n54796 = n50819 & n53439;
  assign n54801 = n54804 & n54777;
  assign n50859 = ~n50819;
  assign n53402 = ~n54832;
  assign n54836 = n54849 & n54850;
  assign n54807 = ~n54855;
  assign n54736 = ~n54856;
  assign n54845 = n54857 & n52031;
  assign n54858 = n54900 ^ n54901;
  assign n54869 = ~n54934;
  assign n54927 = n54813 & n54935;
  assign n54902 = ~n54900;
  assign n54912 = n54944 ^ n54945;
  assign n51167 = n54948 ^ n54949;
  assign n54932 = ~n54813;
  assign n54946 = ~n54944;
  assign n54979 = n54995 & n54996;
  assign n54640 = n54755 ^ n54756;
  assign n54729 = ~n54772;
  assign n54763 = n54778 & n54779;
  assign n53441 = ~n54796;
  assign n54770 = ~n54797;
  assign n54791 = n50859 & n54798;
  assign n54739 = ~n54801;
  assign n54806 = ~n54836;
  assign n54766 = ~n54845;
  assign n54824 = n29 ^ n54858;
  assign n54890 = n54902 & n54903;
  assign n54812 = n54911 ^ n54912;
  assign n54863 = ~n54927;
  assign n54916 = n51167 & n53915;
  assign n54905 = n51167 & n52671;
  assign n54906 = n51167 & n54010;
  assign n54904 = n54932 & n54861;
  assign n51299 = ~n51167;
  assign n54936 = n54946 & n54947;
  assign n54950 = ~n54979;
  assign n54720 = n54640 & n172;
  assign n54706 = ~n54640;
  assign n54702 = n54729 ^ n54730;
  assign n54737 = n54751 & n54729;
  assign n54738 = ~n54763;
  assign n54667 = n54770 & n54771;
  assign n53466 = ~n54791;
  assign n54764 = n54806 & n54807;
  assign n54657 = n54823 ^ n54824;
  assign n54740 = n54824 & n54823;
  assign n54859 = n54812 & n20006;
  assign n54870 = ~n54812;
  assign n54868 = ~n54890;
  assign n54816 = ~n54904;
  assign n53975 = ~n54905;
  assign n54008 = ~n54906;
  assign n54887 = n51299 & n54907;
  assign n54879 = ~n54916;
  assign n54914 = ~n54936;
  assign n54908 = n54950 & n54951;
  assign n54662 = n173 ^ n54702;
  assign n54691 = n54706 & n16911;
  assign n54649 = ~n54720;
  assign n54723 = ~n54737;
  assign n54707 = n54738 & n54739;
  assign n54688 = ~n54667;
  assign n54732 = n54764 ^ n52031;
  assign n54765 = ~n54764;
  assign n54781 = n54657 & n51987;
  assign n54780 = ~n54657;
  assign n54743 = ~n54740;
  assign n54827 = ~n54859;
  assign n54811 = n54868 & n54869;
  assign n54846 = n54870 & n28;
  assign n54748 = n54879 & n54880;
  assign n54034 = ~n54887;
  assign n54865 = n54908 ^ n52613;
  assign n54860 = n54914 & n54915;
  assign n54909 = ~n54908;
  assign n53314 = n54661 ^ n54662;
  assign n54607 = n54662 & n54661;
  assign n54666 = ~n54691;
  assign n54668 = n54707 ^ n54708;
  assign n54664 = n54723 & n54724;
  assign n54709 = n54707 & n54728;
  assign n54722 = ~n54707;
  assign n50785 = n54731 ^ n54732;
  assign n54761 = n54765 & n54766;
  assign n54767 = n54780 & n52050;
  assign n54659 = ~n54781;
  assign n54782 = n54811 ^ n54812;
  assign n54784 = ~n54846;
  assign n54837 = n54748 & n54786;
  assign n54826 = ~n54811;
  assign n54814 = n54860 ^ n54861;
  assign n54833 = ~n54748;
  assign n51106 = n54864 ^ n54865;
  assign n54862 = ~n54860;
  assign n54888 = n54909 & n54910;
  assign n54580 = ~n53314;
  assign n54639 = n172 ^ n54664;
  assign n54590 = n54667 ^ n54668;
  assign n54665 = ~n54664;
  assign n54692 = n50785 & n53398;
  assign n54694 = n50785 & n53308;
  assign n54687 = ~n54709;
  assign n54695 = n50785 & n52031;
  assign n54693 = n54722 & n54708;
  assign n50822 = ~n50785;
  assign n54735 = ~n54761;
  assign n54697 = ~n54767;
  assign n54741 = n28 ^ n54782;
  assign n54745 = n54813 ^ n54814;
  assign n54808 = n54826 & n54827;
  assign n54817 = n54833 & n54834;
  assign n54825 = n51106 & n54835;
  assign n54818 = n51106 & n53884;
  assign n54819 = n51106 & n52547;
  assign n54794 = ~n54837;
  assign n51233 = ~n51106;
  assign n54847 = n54862 & n54863;
  assign n54866 = ~n54888;
  assign n54608 = n54639 ^ n54640;
  assign n54663 = n54665 & n54666;
  assign n54669 = n54687 & n54688;
  assign n53400 = ~n54692;
  assign n54652 = ~n54693;
  assign n54681 = ~n54694;
  assign n53366 = ~n54695;
  assign n54683 = n50822 & n54705;
  assign n54703 = n54735 & n54736;
  assign n54598 = n54740 ^ n54741;
  assign n54742 = ~n54741;
  assign n54790 = n54745 & n27;
  assign n54792 = ~n54745;
  assign n54783 = ~n54808;
  assign n54754 = ~n54817;
  assign n54799 = ~n54818;
  assign n53939 = ~n54819;
  assign n54803 = n51233 & n53965;
  assign n53970 = ~n54825;
  assign n54815 = ~n54847;
  assign n54820 = n54866 & n54867;
  assign n54554 = n54607 ^ n54608;
  assign n54619 = ~n54608;
  assign n54648 = ~n54663;
  assign n54651 = ~n54669;
  assign n54591 = n54681 & n54682;
  assign n53422 = ~n54683;
  assign n54656 = n54703 ^ n52050;
  assign n54696 = ~n54703;
  assign n54710 = n54598 & n52006;
  assign n54717 = ~n54598;
  assign n54670 = n54742 & n54743;
  assign n54744 = n54783 & n54784;
  assign n54713 = ~n54790;
  assign n54769 = n54792 & n19971;
  assign n54674 = n54799 & n54800;
  assign n53995 = ~n54803;
  assign n54785 = n54815 & n54816;
  assign n54788 = n54820 ^ n52598;
  assign n54563 = ~n54554;
  assign n54557 = n54619 & n54607;
  assign n54622 = n54648 & n54649;
  assign n54624 = n54651 & n54652;
  assign n50752 = n54656 ^ n54657;
  assign n54606 = ~n54591;
  assign n54684 = n54696 & n54697;
  assign n54636 = ~n54710;
  assign n54704 = n54717 & n51953;
  assign n54678 = ~n54670;
  assign n54711 = n54744 ^ n54745;
  assign n54746 = ~n54744;
  assign n54747 = ~n54769;
  assign n54749 = n54785 ^ n54786;
  assign n54690 = ~n54674;
  assign n51201 = n54787 ^ n54788;
  assign n54793 = ~n54785;
  assign n54556 = ~n54557;
  assign n54621 = n54622 & n16887;
  assign n54592 = n54624 ^ n54625;
  assign n54604 = ~n54622;
  assign n54629 = n54624 & n54631;
  assign n54630 = n50752 & n54641;
  assign n54633 = n50752 & n52050;
  assign n54626 = ~n54624;
  assign n54632 = n50752 & n53290;
  assign n50761 = ~n50752;
  assign n54658 = ~n54684;
  assign n54602 = ~n54704;
  assign n54671 = n27 ^ n54711;
  assign n54733 = n54746 & n54747;
  assign n54680 = n54748 ^ n54749;
  assign n54752 = n51201 & n52598;
  assign n54750 = n51201 & n54760;
  assign n52652 = ~n51201;
  assign n54768 = n54793 & n54794;
  assign n54529 = n54591 ^ n54592;
  assign n54570 = n54604 ^ n54590;
  assign n54603 = n54604 & n171;
  assign n54589 = ~n54621;
  assign n54620 = n54626 & n54625;
  assign n54605 = ~n54629;
  assign n53357 = ~n54630;
  assign n54609 = ~n54632;
  assign n53313 = ~n54633;
  assign n54623 = n50761 & n53378;
  assign n54634 = n54658 & n54659;
  assign n54653 = n54670 ^ n54671;
  assign n54677 = ~n54671;
  assign n54714 = n54680 & n19943;
  assign n54712 = ~n54733;
  assign n54715 = ~n54680;
  assign n54699 = n54734 ^ n52652;
  assign n54725 = ~n54750;
  assign n53922 = ~n54752;
  assign n54753 = ~n54768;
  assign n54558 = n171 ^ n54570;
  assign n54587 = n54589 & n54590;
  assign n54565 = ~n54603;
  assign n54593 = n54605 & n54606;
  assign n54526 = n54609 & n54610;
  assign n54572 = ~n54620;
  assign n53380 = ~n54623;
  assign n54597 = n54634 ^ n52006;
  assign n54642 = n54653 & n51911;
  assign n54635 = ~n54634;
  assign n54650 = ~n54653;
  assign n54611 = n54677 & n54678;
  assign n53952 = n54699 ^ n54700;
  assign n54679 = n54712 & n54713;
  assign n54673 = ~n54714;
  assign n54698 = n54715 & n26;
  assign n54685 = n54725 & n54726;
  assign n54721 = n54753 & n54754;
  assign n53244 = n54557 ^ n54558;
  assign n54555 = ~n54558;
  assign n54564 = ~n54587;
  assign n54571 = ~n54593;
  assign n54588 = n54526 & n54545;
  assign n54581 = ~n54526;
  assign n50705 = n54597 ^ n54598;
  assign n54627 = n54635 & n54636;
  assign n54553 = ~n54642;
  assign n54638 = n54650 & n51921;
  assign n54614 = ~n54611;
  assign n54643 = n54679 ^ n54680;
  assign n54596 = n54685 ^ n54686;
  assign n54645 = ~n54698;
  assign n54672 = ~n54679;
  assign n54675 = n54721 ^ n54719;
  assign n54716 = n54721 & n54727;
  assign n54718 = ~n54721;
  assign n54490 = ~n53244;
  assign n54488 = n54555 & n54556;
  assign n54543 = n54564 & n54565;
  assign n54544 = n54571 & n54572;
  assign n54579 = n50705 & n54580;
  assign n54573 = n54581 & n54582;
  assign n54547 = ~n54588;
  assign n50741 = ~n50705;
  assign n54601 = ~n54627;
  assign n54575 = ~n54638;
  assign n54612 = n26 ^ n54643;
  assign n54660 = n54672 & n54673;
  assign n54616 = n54674 ^ n54675;
  assign n54689 = ~n54716;
  assign n54701 = n54718 & n54719;
  assign n54493 = ~n54488;
  assign n54541 = n54543 & n16859;
  assign n54527 = n54544 ^ n54545;
  assign n54535 = ~n54543;
  assign n54546 = ~n54544;
  assign n54566 = n50741 & n53314;
  assign n54519 = ~n54573;
  assign n54568 = n50741 & n52006;
  assign n53337 = ~n54579;
  assign n54567 = n50741 & n53252;
  assign n54577 = n54601 & n54602;
  assign n54594 = n54611 ^ n54612;
  assign n54599 = n54575 & n54553;
  assign n54613 = ~n54612;
  assign n54647 = n54616 & n25;
  assign n54644 = ~n54660;
  assign n54646 = ~n54616;
  assign n54676 = n54689 & n54690;
  assign n54655 = ~n54701;
  assign n54475 = n54526 ^ n54527;
  assign n54508 = n54535 ^ n54529;
  assign n54538 = n54535 & n170;
  assign n54528 = ~n54541;
  assign n54540 = n54546 & n54547;
  assign n53317 = ~n54566;
  assign n54548 = ~n54567;
  assign n53278 = ~n54568;
  assign n54574 = ~n54577;
  assign n54583 = n54594 & n51932;
  assign n54578 = ~n54599;
  assign n54500 = ~n54594;
  assign n54561 = n54613 & n54614;
  assign n54615 = n54644 & n54645;
  assign n54637 = n54646 & n19881;
  assign n54586 = ~n54647;
  assign n54654 = ~n54676;
  assign n54489 = n170 ^ n54508;
  assign n54494 = n54475 & n16793;
  assign n54505 = ~n54475;
  assign n54514 = n54528 & n54529;
  assign n54507 = ~n54538;
  assign n54518 = ~n54540;
  assign n54478 = n54548 & n54549;
  assign n54569 = n54574 & n54575;
  assign n50641 = n54577 ^ n54578;
  assign n54525 = ~n54583;
  assign n54576 = n54500 & n51842;
  assign n54584 = n54615 ^ n54616;
  assign n54617 = ~n54615;
  assign n54618 = ~n54637;
  assign n54628 = n54654 & n54655;
  assign n53205 = n54488 ^ n54489;
  assign n54437 = n54489 & n54493;
  assign n54477 = ~n54494;
  assign n54492 = n54505 & n169;
  assign n54506 = ~n54514;
  assign n54495 = n54518 & n54519;
  assign n54521 = n54478 & n54530;
  assign n54520 = ~n54478;
  assign n54550 = n50641 & n53155;
  assign n54551 = n50641 & n51921;
  assign n54542 = n50641 & n54563;
  assign n50708 = ~n50641;
  assign n54552 = ~n54569;
  assign n54503 = ~n54576;
  assign n54562 = n25 ^ n54584;
  assign n54600 = n54617 & n54618;
  assign n54595 = n24 ^ n54628;
  assign n54453 = ~n53205;
  assign n54468 = ~n54492;
  assign n54479 = n54495 ^ n54496;
  assign n54474 = n54506 & n54507;
  assign n54497 = ~n54495;
  assign n54515 = n54520 & n54496;
  assign n54498 = ~n54521;
  assign n53266 = ~n54542;
  assign n54536 = ~n54550;
  assign n53255 = ~n54551;
  assign n54522 = n54552 & n54553;
  assign n54539 = n50708 & n54554;
  assign n54458 = n54561 ^ n54562;
  assign n54533 = n54562 & n54561;
  assign n54560 = n54595 ^ n54596;
  assign n54585 = ~n54600;
  assign n54462 = n54474 ^ n54475;
  assign n54440 = n54478 ^ n54479;
  assign n54476 = ~n54474;
  assign n54491 = n54497 & n54498;
  assign n54486 = ~n54515;
  assign n54499 = n54522 ^ n51932;
  assign n54457 = n54536 & n54537;
  assign n53299 = ~n54539;
  assign n54532 = n54458 & n51823;
  assign n54524 = ~n54522;
  assign n54531 = ~n54458;
  assign n54559 = n54585 & n54586;
  assign n54438 = n169 ^ n54462;
  assign n54466 = n54440 & n168;
  assign n54465 = ~n54440;
  assign n54473 = n54476 & n54477;
  assign n54485 = ~n54491;
  assign n50620 = n54499 ^ n54500;
  assign n54513 = n54457 & n54449;
  assign n54509 = ~n54457;
  assign n54517 = n53266 & n53299;
  assign n54516 = n54524 & n54525;
  assign n54523 = n54531 & n51883;
  assign n54483 = ~n54532;
  assign n54534 = n54559 ^ n54560;
  assign n53142 = n54437 ^ n54438;
  assign n54403 = n54438 & n54437;
  assign n54454 = n54465 & n16739;
  assign n54428 = ~n54466;
  assign n54467 = ~n54473;
  assign n54456 = n54485 & n54486;
  assign n54487 = n50620 & n54490;
  assign n54480 = n50620 & n53117;
  assign n54484 = n50620 & n51932;
  assign n50672 = ~n50620;
  assign n54501 = n54509 & n54510;
  assign n54464 = ~n54513;
  assign n54502 = ~n54516;
  assign n53297 = ~n54517;
  assign n54461 = ~n54523;
  assign n54423 = n54533 ^ n54534;
  assign n54415 = ~n53142;
  assign n54451 = ~n54454;
  assign n54448 = n54456 ^ n54457;
  assign n54439 = n54467 & n54468;
  assign n54463 = ~n54456;
  assign n54471 = n50672 & n53244;
  assign n54469 = ~n54480;
  assign n53195 = ~n54484;
  assign n53225 = ~n54487;
  assign n54442 = ~n54501;
  assign n54481 = n54502 & n54503;
  assign n54511 = n54423 & n51846;
  assign n54512 = ~n54423;
  assign n54430 = n54439 ^ n54440;
  assign n54378 = n54448 ^ n54449;
  assign n54450 = ~n54439;
  assign n54455 = n54463 & n54464;
  assign n54405 = n54469 & n54470;
  assign n53246 = ~n54471;
  assign n54459 = n54481 ^ n51883;
  assign n54482 = ~n54481;
  assign n54426 = ~n54511;
  assign n54504 = n54512 & n51781;
  assign n54404 = n168 ^ n54430;
  assign n54418 = n54378 & n16715;
  assign n54429 = ~n54378;
  assign n54435 = n54450 & n54451;
  assign n54441 = ~n54455;
  assign n54414 = ~n54405;
  assign n50534 = n54458 ^ n54459;
  assign n54472 = n54482 & n54483;
  assign n54446 = ~n54504;
  assign n53126 = n54403 ^ n54404;
  assign n54409 = ~n54404;
  assign n54398 = ~n54418;
  assign n54416 = n54429 & n183;
  assign n54427 = ~n54435;
  assign n54419 = n54441 & n54442;
  assign n54443 = n50534 & n53102;
  assign n54444 = n50534 & n51823;
  assign n54447 = n50534 & n54453;
  assign n50623 = ~n50534;
  assign n54460 = ~n54472;
  assign n54375 = ~n53126;
  assign n54353 = n54409 & n54403;
  assign n54388 = ~n54416;
  assign n54406 = n54419 ^ n54420;
  assign n54397 = n54427 & n54428;
  assign n54422 = n54419 & n54433;
  assign n54421 = ~n54419;
  assign n54431 = ~n54443;
  assign n53153 = ~n54444;
  assign n54434 = n50623 & n53205;
  assign n53185 = ~n54447;
  assign n54452 = n54460 & n54461;
  assign n54368 = ~n54353;
  assign n54377 = n183 ^ n54397;
  assign n54357 = n54405 ^ n54406;
  assign n54399 = ~n54397;
  assign n54417 = n54421 & n54420;
  assign n54413 = ~n54422;
  assign n54344 = n54431 & n54432;
  assign n53207 = ~n54434;
  assign n54424 = n54452 ^ n51846;
  assign n54445 = ~n54452;
  assign n54354 = n54377 ^ n54378;
  assign n54379 = n54357 & n182;
  assign n54382 = ~n54357;
  assign n54392 = n54398 & n54399;
  assign n54400 = n54413 & n54414;
  assign n54390 = ~n54417;
  assign n54412 = n54344 & n54370;
  assign n54410 = ~n54344;
  assign n50510 = n54423 ^ n54424;
  assign n54436 = n54445 & n54446;
  assign n54299 = n54353 ^ n54354;
  assign n54367 = ~n54354;
  assign n54341 = ~n54379;
  assign n54376 = n54382 & n16633;
  assign n54387 = ~n54392;
  assign n54389 = ~n54400;
  assign n54401 = n54410 & n54411;
  assign n54372 = ~n54412;
  assign n54396 = n50510 & n54415;
  assign n50571 = ~n50510;
  assign n54425 = ~n54436;
  assign n53062 = ~n54299;
  assign n54321 = n54367 & n54368;
  assign n54365 = ~n54376;
  assign n54356 = n54387 & n54388;
  assign n54369 = n54389 & n54390;
  assign n53165 = ~n54396;
  assign n54347 = ~n54401;
  assign n54395 = n50571 & n53038;
  assign n54393 = n50571 & n51781;
  assign n54391 = n50571 & n53142;
  assign n54402 = n54425 & n54426;
  assign n54338 = n54356 ^ n54357;
  assign n54345 = n54369 ^ n54370;
  assign n54364 = ~n54356;
  assign n54371 = ~n54369;
  assign n53145 = ~n54391;
  assign n53115 = ~n54393;
  assign n54383 = ~n54395;
  assign n54386 = n54402 ^ n51738;
  assign n54407 = ~n54402;
  assign n54322 = n182 ^ n54338;
  assign n54315 = n54344 ^ n54345;
  assign n54350 = n54364 & n54365;
  assign n54358 = n54371 & n54372;
  assign n54311 = n54383 & n54384;
  assign n50490 = n54385 ^ n54386;
  assign n54394 = n54407 & n54408;
  assign n54282 = n54321 ^ n54322;
  assign n54280 = n54322 & n54321;
  assign n54324 = n54315 & n16558;
  assign n54325 = ~n54315;
  assign n54340 = ~n54350;
  assign n54346 = ~n54358;
  assign n54359 = n50490 & n52999;
  assign n54360 = n54311 & n54373;
  assign n54361 = n50490 & n51738;
  assign n54355 = n50490 & n54375;
  assign n54366 = ~n54311;
  assign n50441 = ~n50490;
  assign n54380 = ~n54394;
  assign n53022 = ~n54282;
  assign n54318 = ~n54324;
  assign n54323 = n54325 & n181;
  assign n54335 = n54340 & n54341;
  assign n54326 = n54346 & n54347;
  assign n54349 = n50441 & n53126;
  assign n53108 = ~n54355;
  assign n54342 = ~n54359;
  assign n54332 = ~n54360;
  assign n53073 = ~n54361;
  assign n54351 = n54366 & n54327;
  assign n54374 = n54380 & n54381;
  assign n54303 = ~n54323;
  assign n54312 = n54326 ^ n54327;
  assign n54314 = ~n54335;
  assign n54331 = ~n54326;
  assign n54274 = n54342 & n54343;
  assign n53128 = ~n54349;
  assign n54307 = ~n54351;
  assign n54363 = n54374 & n51695;
  assign n54362 = ~n54374;
  assign n54279 = n54311 ^ n54312;
  assign n54298 = n54314 ^ n54315;
  assign n54313 = n54318 & n54314;
  assign n54319 = n54331 & n54332;
  assign n54330 = n54274 & n54290;
  assign n54328 = ~n54274;
  assign n54352 = n54362 & n51767;
  assign n54339 = ~n54363;
  assign n54281 = n181 ^ n54298;
  assign n54287 = n54279 & n180;
  assign n54297 = ~n54279;
  assign n54302 = ~n54313;
  assign n54306 = ~n54319;
  assign n54320 = n54328 & n54329;
  assign n54294 = ~n54330;
  assign n54337 = n54339 & n54348;
  assign n54334 = ~n54352;
  assign n54240 = n54280 ^ n54281;
  assign n54241 = n54281 & n54280;
  assign n54261 = ~n54287;
  assign n54283 = n54297 & n16510;
  assign n54278 = n54302 & n54303;
  assign n54289 = n54306 & n54307;
  assign n54270 = ~n54320;
  assign n54333 = ~n54337;
  assign n54336 = n54334 & n54339;
  assign n52980 = ~n54240;
  assign n54262 = n54278 ^ n54279;
  assign n54272 = ~n54283;
  assign n54273 = ~n54278;
  assign n54275 = n54289 ^ n54290;
  assign n54293 = ~n54289;
  assign n54308 = n54333 & n54334;
  assign n54317 = ~n54336;
  assign n54242 = n180 ^ n54262;
  assign n54264 = n54272 & n54273;
  assign n54227 = n54274 ^ n54275;
  assign n54284 = n54293 & n54294;
  assign n54295 = n54308 ^ n51651;
  assign n50369 = n54316 ^ n54317;
  assign n54309 = ~n54308;
  assign n54215 = n54241 ^ n54242;
  assign n54181 = n54242 & n54241;
  assign n54247 = n54227 & n16437;
  assign n54260 = ~n54264;
  assign n54248 = ~n54227;
  assign n54269 = ~n54284;
  assign n50288 = n54295 ^ n54296;
  assign n54304 = n50369 & n53062;
  assign n54300 = n50369 & n53015;
  assign n54301 = n50369 & n51695;
  assign n54305 = n54309 & n54310;
  assign n50451 = ~n50369;
  assign n52966 = ~n54215;
  assign n54199 = ~n54181;
  assign n54239 = ~n54247;
  assign n54245 = n54248 & n179;
  assign n54226 = n54260 & n54261;
  assign n54256 = n54269 & n54270;
  assign n54268 = n50288 & n54282;
  assign n50373 = ~n50288;
  assign n54288 = n50451 & n54299;
  assign n54285 = ~n54300;
  assign n53033 = ~n54301;
  assign n53064 = ~n54304;
  assign n54291 = ~n54305;
  assign n54216 = n54226 ^ n54227;
  assign n54206 = ~n54245;
  assign n54238 = ~n54226;
  assign n54229 = n54256 ^ n54257;
  assign n54249 = n54256 & n54257;
  assign n54258 = ~n54256;
  assign n53047 = ~n54268;
  assign n54265 = n50373 & n52971;
  assign n54266 = n50373 & n51725;
  assign n54263 = n50373 & n53022;
  assign n54228 = n54285 & n54286;
  assign n53087 = ~n54288;
  assign n54271 = n54291 & n54292;
  assign n54182 = n179 ^ n54216;
  assign n54184 = n54228 ^ n54229;
  assign n54219 = n54238 & n54239;
  assign n54243 = ~n54249;
  assign n54246 = n54258 & n54259;
  assign n53025 = ~n54263;
  assign n54250 = ~n54265;
  assign n52991 = ~n54266;
  assign n54253 = n54271 ^ n51674;
  assign n54244 = ~n54228;
  assign n54276 = ~n54271;
  assign n52923 = n54181 ^ n54182;
  assign n54153 = n54182 & n54199;
  assign n54207 = n54184 & n16378;
  assign n54205 = ~n54219;
  assign n54208 = ~n54184;
  assign n54230 = n54243 & n54244;
  assign n54218 = ~n54246;
  assign n54176 = n54250 & n54251;
  assign n50213 = n54252 ^ n54253;
  assign n54267 = n54276 & n54277;
  assign n54155 = ~n52923;
  assign n54144 = ~n54153;
  assign n54183 = n54205 & n54206;
  assign n54191 = ~n54207;
  assign n54204 = n54208 & n178;
  assign n54217 = ~n54230;
  assign n54225 = n50213 & n54240;
  assign n54233 = n54176 & n54196;
  assign n54231 = ~n54176;
  assign n50292 = ~n50213;
  assign n54254 = ~n54267;
  assign n54167 = n54183 ^ n54184;
  assign n54169 = ~n54204;
  assign n54192 = ~n54183;
  assign n54195 = n54217 & n54218;
  assign n54223 = n50292 & n52980;
  assign n53009 = ~n54225;
  assign n54220 = n54231 & n54232;
  assign n54221 = n50292 & n52879;
  assign n54222 = n50292 & n51602;
  assign n54201 = ~n54233;
  assign n54236 = n54254 & n54255;
  assign n54154 = n178 ^ n54167;
  assign n54178 = n54191 & n54192;
  assign n54177 = n54195 ^ n54196;
  assign n54200 = ~n54195;
  assign n54172 = ~n54220;
  assign n54209 = ~n54221;
  assign n52947 = ~n54222;
  assign n52983 = ~n54223;
  assign n50126 = n54236 ^ n54237;
  assign n54234 = ~n54236;
  assign n52861 = n54153 ^ n54154;
  assign n54143 = ~n54154;
  assign n54140 = n54176 ^ n54177;
  assign n54168 = ~n54178;
  assign n54190 = n54200 & n54201;
  assign n54132 = n54209 & n54210;
  assign n54211 = n50126 & n52835;
  assign n54214 = n50126 & n52966;
  assign n50140 = ~n50126;
  assign n54224 = n54234 & n54235;
  assign n54121 = ~n52861;
  assign n54108 = n54143 & n54144;
  assign n54156 = n54140 & n16277;
  assign n54157 = ~n54140;
  assign n54162 = n54168 & n54169;
  assign n54171 = ~n54190;
  assign n54187 = n54132 & n54159;
  assign n54185 = ~n54132;
  assign n54197 = ~n54211;
  assign n54203 = n50140 & n51552;
  assign n52941 = ~n54214;
  assign n54202 = n50140 & n54215;
  assign n54212 = ~n54224;
  assign n54107 = ~n54108;
  assign n54142 = ~n54156;
  assign n54146 = n54157 & n177;
  assign n54139 = ~n54162;
  assign n54158 = n54171 & n54172;
  assign n54179 = n54185 & n54186;
  assign n54161 = ~n54187;
  assign n54120 = n54197 & n54198;
  assign n52968 = ~n54202;
  assign n52903 = ~n54203;
  assign n54188 = n54212 & n54213;
  assign n54126 = n54139 ^ n54140;
  assign n54131 = n54142 & n54139;
  assign n54125 = ~n54146;
  assign n54133 = n54158 ^ n54159;
  assign n54160 = ~n54158;
  assign n54135 = ~n54179;
  assign n54175 = n54120 & n54099;
  assign n54173 = ~n54120;
  assign n54170 = n54188 ^ n54189;
  assign n54193 = ~n54188;
  assign n54109 = n177 ^ n54126;
  assign n54124 = ~n54131;
  assign n54102 = n54132 ^ n54133;
  assign n54147 = n54160 & n54161;
  assign n49964 = n51418 ^ n54170;
  assign n54163 = n54173 & n54174;
  assign n54123 = ~n54175;
  assign n54164 = n54170 & n51582;
  assign n54180 = n54193 & n54194;
  assign n52819 = n54108 ^ n54109;
  assign n54106 = ~n54109;
  assign n54101 = n54124 & n54125;
  assign n54117 = n54102 & n16229;
  assign n54118 = ~n54102;
  assign n54134 = ~n54147;
  assign n54145 = n49964 & n54155;
  assign n54148 = n49964 & n52765;
  assign n50141 = ~n49964;
  assign n54095 = ~n54163;
  assign n52866 = ~n54164;
  assign n54165 = ~n54180;
  assign n54067 = ~n52819;
  assign n54088 = n54101 ^ n54102;
  assign n54059 = n54106 & n54107;
  assign n54104 = ~n54101;
  assign n54105 = ~n54117;
  assign n54116 = n54118 & n176;
  assign n54119 = n54134 & n54135;
  assign n54138 = n50141 & n52923;
  assign n52901 = ~n54145;
  assign n54136 = ~n54148;
  assign n54149 = n54165 & n54166;
  assign n54060 = n176 ^ n54088;
  assign n54093 = n54104 & n54105;
  assign n54087 = ~n54116;
  assign n54098 = n54119 ^ n54120;
  assign n54122 = ~n54119;
  assign n54077 = n54136 & n54137;
  assign n52925 = ~n54138;
  assign n54127 = n54149 ^ n54150;
  assign n54151 = ~n54149;
  assign n52779 = n54059 ^ n54060;
  assign n54015 = n54060 & n54059;
  assign n54086 = ~n54093;
  assign n54044 = n54098 ^ n54099;
  assign n54111 = n54122 & n54123;
  assign n54062 = ~n54077;
  assign n49917 = n51518 ^ n54127;
  assign n54130 = n54127 & n51389;
  assign n54141 = n54151 & n54152;
  assign n54038 = ~n52779;
  assign n54065 = n54086 & n54087;
  assign n54076 = n54044 & n16084;
  assign n54083 = ~n54044;
  assign n54094 = ~n54111;
  assign n54112 = n49917 & n52739;
  assign n54110 = n49917 & n54121;
  assign n50041 = ~n49917;
  assign n52824 = ~n54130;
  assign n54128 = ~n54141;
  assign n54043 = n191 ^ n54065;
  assign n54063 = ~n54065;
  assign n54064 = ~n54076;
  assign n54068 = n54083 & n191;
  assign n54078 = n54094 & n54095;
  assign n54100 = n50041 & n52861;
  assign n52864 = ~n54110;
  assign n54096 = ~n54112;
  assign n54113 = n54128 & n54129;
  assign n54016 = n54043 ^ n54044;
  assign n54051 = n54063 & n54064;
  assign n54041 = ~n54068;
  assign n54055 = n54077 ^ n54078;
  assign n54081 = n54078 & n54056;
  assign n54079 = ~n54078;
  assign n54005 = n54096 & n54097;
  assign n52884 = ~n54100;
  assign n54092 = n54113 ^ n51310;
  assign n54114 = ~n54113;
  assign n52732 = n54015 ^ n54016;
  assign n53985 = n54016 & n54015;
  assign n54040 = ~n54051;
  assign n54018 = n54055 ^ n54056;
  assign n54069 = n54079 & n54080;
  assign n54061 = ~n54081;
  assign n54082 = n54005 & n54020;
  assign n54084 = ~n54005;
  assign n49836 = n54091 ^ n54092;
  assign n54103 = n54114 & n54115;
  assign n53989 = ~n52732;
  assign n53977 = ~n53985;
  assign n54035 = n54018 & n16051;
  assign n54017 = n54040 & n54041;
  assign n54036 = ~n54018;
  assign n54054 = n54061 & n54062;
  assign n54046 = ~n54069;
  assign n54066 = n49836 & n52819;
  assign n54026 = ~n54082;
  assign n54075 = n54084 & n54085;
  assign n54071 = n49836 & n51310;
  assign n54070 = n49836 & n52755;
  assign n49967 = ~n49836;
  assign n54089 = ~n54103;
  assign n54000 = n54017 ^ n54018;
  assign n54027 = ~n54017;
  assign n54028 = ~n54035;
  assign n54030 = n54036 & n190;
  assign n54045 = ~n54054;
  assign n52822 = ~n54066;
  assign n54057 = n49967 & n54067;
  assign n54052 = ~n54070;
  assign n52777 = ~n54071;
  assign n54004 = ~n54075;
  assign n54072 = n54089 & n54090;
  assign n53986 = n190 ^ n54000;
  assign n54013 = n54027 & n54028;
  assign n54002 = ~n54030;
  assign n54019 = n54045 & n54046;
  assign n53961 = n54052 & n54053;
  assign n52843 = ~n54057;
  assign n54047 = n54072 ^ n51379;
  assign n54073 = ~n54072;
  assign n53947 = n53985 ^ n53986;
  assign n53976 = ~n53986;
  assign n54001 = ~n54013;
  assign n54006 = n54019 ^ n54020;
  assign n54025 = ~n54019;
  assign n54037 = n53961 & n54042;
  assign n54039 = ~n53961;
  assign n49753 = n54047 ^ n54048;
  assign n54058 = n54073 & n54074;
  assign n52688 = ~n53947;
  assign n53936 = n53976 & n53977;
  assign n53999 = n54001 & n54002;
  assign n53971 = n54005 ^ n54006;
  assign n54014 = n54025 & n54026;
  assign n53983 = ~n54037;
  assign n54029 = n49753 & n54038;
  assign n54031 = n54039 & n53980;
  assign n49865 = ~n49753;
  assign n54049 = ~n54058;
  assign n53988 = n53971 & n15951;
  assign n53968 = ~n53999;
  assign n53987 = ~n53971;
  assign n54003 = ~n54014;
  assign n52801 = ~n54029;
  assign n53964 = ~n54031;
  assign n54024 = n49865 & n52779;
  assign n54021 = n49865 & n52721;
  assign n54022 = n49865 & n51379;
  assign n54032 = n54049 & n54050;
  assign n53956 = n53968 ^ n53971;
  assign n53972 = n53987 & n189;
  assign n53967 = ~n53988;
  assign n53979 = n54003 & n54004;
  assign n54011 = ~n54021;
  assign n52741 = ~n54022;
  assign n52782 = ~n54024;
  assign n54009 = n54032 ^ n51299;
  assign n54033 = ~n54032;
  assign n53937 = n189 ^ n53956;
  assign n53960 = n53967 & n53968;
  assign n53954 = ~n53972;
  assign n53962 = n53979 ^ n53980;
  assign n53982 = ~n53979;
  assign n49781 = n54009 ^ n54010;
  assign n53927 = n54011 & n54012;
  assign n54023 = n54033 & n54034;
  assign n53919 = n53936 ^ n53937;
  assign n53902 = n53937 & n53936;
  assign n53953 = ~n53960;
  assign n53930 = n53961 ^ n53962;
  assign n53973 = n53982 & n53983;
  assign n53998 = n49781 & n52732;
  assign n53991 = n49781 & n52590;
  assign n53990 = n53927 & n53944;
  assign n53992 = n49781 & n51299;
  assign n53996 = ~n53927;
  assign n49675 = ~n49781;
  assign n54007 = ~n54023;
  assign n53905 = ~n53902;
  assign n53942 = n53930 & n188;
  assign n53929 = n53953 & n53954;
  assign n53941 = ~n53930;
  assign n53963 = ~n53973;
  assign n53978 = n49675 & n53989;
  assign n53946 = ~n53990;
  assign n53974 = ~n53991;
  assign n52687 = ~n53992;
  assign n53984 = n53996 & n53997;
  assign n52735 = ~n53998;
  assign n53993 = n54007 & n54008;
  assign n53918 = n53929 ^ n53930;
  assign n53933 = n53941 & n15860;
  assign n53911 = ~n53942;
  assign n53924 = ~n53929;
  assign n53943 = n53963 & n53964;
  assign n53898 = n53974 & n53975;
  assign n52763 = ~n53978;
  assign n53926 = ~n53984;
  assign n53966 = n53993 ^ n51106;
  assign n53994 = ~n53993;
  assign n53903 = n188 ^ n53918;
  assign n53923 = ~n53933;
  assign n53928 = n53943 ^ n53944;
  assign n53945 = ~n53943;
  assign n53957 = n53898 & n53959;
  assign n53958 = ~n53898;
  assign n49605 = n53965 ^ n53966;
  assign n53981 = n53994 & n53995;
  assign n53892 = n53902 ^ n53903;
  assign n53904 = ~n53903;
  assign n53920 = n53923 & n53924;
  assign n53895 = n53927 ^ n53928;
  assign n53934 = n53945 & n53946;
  assign n53955 = n49605 & n52688;
  assign n53917 = ~n53957;
  assign n53950 = n49605 & n51233;
  assign n53949 = n49605 & n52613;
  assign n53948 = n53958 & n53915;
  assign n49702 = ~n49605;
  assign n53969 = ~n53981;
  assign n50634 = n53892 ^ n51616;
  assign n53823 = n53892 & n51614;
  assign n53891 = n53892 & n51616;
  assign n53875 = n53904 & n53905;
  assign n53912 = n53895 & n15777;
  assign n53910 = ~n53920;
  assign n53913 = ~n53895;
  assign n53925 = ~n53934;
  assign n53940 = n49702 & n53947;
  assign n53901 = ~n53948;
  assign n53938 = ~n53949;
  assign n52634 = ~n53950;
  assign n52723 = ~n53955;
  assign n53951 = n53969 & n53970;
  assign n50636 = ~n50634;
  assign n52706 = ~n53891;
  assign n53874 = ~n53875;
  assign n53894 = n53910 & n53911;
  assign n53896 = ~n53912;
  assign n53906 = n53913 & n187;
  assign n53914 = n53925 & n53926;
  assign n53870 = n53938 & n53939;
  assign n52697 = ~n53940;
  assign n49647 = n53951 ^ n53952;
  assign n53865 = n50636 & n52680;
  assign n53881 = n53894 ^ n53895;
  assign n53889 = ~n53906;
  assign n53897 = ~n53894;
  assign n53899 = n53914 ^ n53915;
  assign n53916 = ~n53914;
  assign n53878 = ~n53870;
  assign n53932 = n49647 & n51201;
  assign n53931 = n49647 & n53935;
  assign n51273 = ~n49647;
  assign n53859 = ~n53865;
  assign n53876 = n187 ^ n53881;
  assign n53893 = n53896 & n53897;
  assign n53867 = n53898 ^ n53899;
  assign n53907 = n53916 & n53917;
  assign n52674 = n53919 ^ n51273;
  assign n53921 = ~n53931;
  assign n52625 = ~n53932;
  assign n53845 = n53859 & n53860;
  assign n53861 = n53875 ^ n53876;
  assign n53873 = ~n53876;
  assign n53882 = n53867 & n186;
  assign n53888 = ~n53893;
  assign n53887 = ~n53867;
  assign n53900 = ~n53907;
  assign n53908 = n53921 & n53922;
  assign n53829 = n53845 ^ n53846;
  assign n53848 = ~n53845;
  assign n53852 = n53861 & n51523;
  assign n53853 = ~n53861;
  assign n53837 = n53873 & n53874;
  assign n53856 = ~n53882;
  assign n53879 = n53887 & n15671;
  assign n53866 = n53888 & n53889;
  assign n53883 = n53900 & n53901;
  assign n53833 = n53908 ^ n53909;
  assign n52258 = n327 ^ n53829;
  assign n53721 = n53829 & n327;
  assign n53770 = n53848 & n53849;
  assign n53836 = ~n53852;
  assign n53850 = n53853 & n51514;
  assign n53840 = ~n53837;
  assign n53854 = n53866 ^ n53867;
  assign n53868 = ~n53866;
  assign n53869 = ~n53879;
  assign n53871 = n53883 ^ n53884;
  assign n53886 = n53883 & n53890;
  assign n53885 = ~n53883;
  assign n52285 = ~n52258;
  assign n53835 = n53836 & n53823;
  assign n53831 = ~n53850;
  assign n53838 = n186 ^ n53854;
  assign n53864 = n53868 & n53869;
  assign n53842 = n53870 ^ n53871;
  assign n53880 = n53885 & n53884;
  assign n53877 = ~n53886;
  assign n53830 = ~n53835;
  assign n53822 = n53831 & n53836;
  assign n53810 = n53837 ^ n53838;
  assign n53839 = ~n53838;
  assign n53858 = n53842 & n185;
  assign n53855 = ~n53864;
  assign n53857 = ~n53842;
  assign n53872 = n53877 & n53878;
  assign n53863 = ~n53880;
  assign n50516 = n53822 ^ n53823;
  assign n53819 = n53830 & n53831;
  assign n53825 = n53810 & n51449;
  assign n53824 = ~n53810;
  assign n53815 = n53839 & n53840;
  assign n53841 = n53855 & n53856;
  assign n53851 = n53857 & n15638;
  assign n53828 = ~n53858;
  assign n53862 = ~n53872;
  assign n53813 = n50516 & n52585;
  assign n53814 = n50516 & n51523;
  assign n53811 = n53819 ^ n51414;
  assign n50522 = ~n50516;
  assign n53817 = ~n53819;
  assign n53821 = n53824 & n51414;
  assign n53803 = ~n53825;
  assign n53820 = ~n53815;
  assign n53826 = n53841 ^ n53842;
  assign n53844 = ~n53851;
  assign n53843 = ~n53841;
  assign n53847 = n53862 & n53863;
  assign n50419 = n53810 ^ n53811;
  assign n53806 = ~n53813;
  assign n52616 = ~n53814;
  assign n53818 = ~n53821;
  assign n53816 = n185 ^ n53826;
  assign n53834 = n53843 & n53844;
  assign n53832 = n184 ^ n53847;
  assign n53793 = n50419 & n51414;
  assign n53792 = n50419 & n52534;
  assign n50463 = ~n50419;
  assign n53800 = n53806 & n53807;
  assign n53776 = n53815 ^ n53816;
  assign n53812 = n53817 & n53818;
  assign n53809 = n53816 & n53820;
  assign n53798 = n53832 ^ n53833;
  assign n53827 = ~n53834;
  assign n53785 = ~n53792;
  assign n52556 = ~n53793;
  assign n53794 = n53800 & n53801;
  assign n53795 = ~n53800;
  assign n53804 = n53776 & n51342;
  assign n53802 = ~n53812;
  assign n53805 = ~n53776;
  assign n53808 = n53827 & n53828;
  assign n53742 = n53785 & n53786;
  assign n53784 = ~n53794;
  assign n53788 = n53795 & n53796;
  assign n53789 = n53802 & n53803;
  assign n53780 = ~n53804;
  assign n53799 = n53805 & n51384;
  assign n53797 = n53808 ^ n53809;
  assign n53772 = n53742 & n53778;
  assign n53771 = ~n53742;
  assign n53781 = n53784 & n53770;
  assign n53774 = ~n53788;
  assign n53775 = n53789 ^ n51384;
  assign n53748 = n53797 ^ n53798;
  assign n53790 = ~n53789;
  assign n53791 = ~n53799;
  assign n53767 = n53771 & n53756;
  assign n53761 = ~n53772;
  assign n50382 = n53775 ^ n53776;
  assign n53773 = ~n53781;
  assign n53769 = n53774 & n53784;
  assign n53783 = n53748 & n51264;
  assign n53782 = ~n53748;
  assign n53787 = n53790 & n53791;
  assign n53746 = ~n53767;
  assign n53762 = n50382 & n52460;
  assign n53759 = n53769 ^ n53770;
  assign n53763 = n50382 & n51384;
  assign n50339 = ~n50382;
  assign n53768 = n53773 & n53774;
  assign n53777 = n53782 & n51292;
  assign n53765 = ~n53783;
  assign n53779 = ~n53787;
  assign n53757 = n53759 & n326;
  assign n53752 = ~n53762;
  assign n52486 = ~n53763;
  assign n53754 = ~n53759;
  assign n53755 = ~n53768;
  assign n53751 = ~n53777;
  assign n53766 = n53779 & n53780;
  assign n53709 = n53752 & n53753;
  assign n53747 = n53754 & n13593;
  assign n53743 = n53755 ^ n53756;
  assign n53719 = ~n53757;
  assign n53758 = n53761 & n53755;
  assign n53749 = n53766 ^ n51292;
  assign n53764 = ~n53766;
  assign n53699 = n53742 ^ n53743;
  assign n53739 = n53709 & n53729;
  assign n53744 = ~n53747;
  assign n50251 = n53748 ^ n53749;
  assign n53740 = ~n53709;
  assign n53745 = ~n53758;
  assign n53760 = n53764 & n53765;
  assign n53724 = n53699 & n13543;
  assign n53725 = ~n53699;
  assign n53731 = ~n53739;
  assign n53735 = n53740 & n53741;
  assign n53734 = n53744 & n53721;
  assign n53720 = n53744 & n53719;
  assign n53736 = n50251 & n52411;
  assign n53737 = n50251 & n51264;
  assign n50295 = ~n50251;
  assign n53728 = n53745 & n53746;
  assign n53750 = ~n53760;
  assign n53701 = n53720 ^ n53721;
  assign n53702 = ~n53724;
  assign n53716 = n53725 & n325;
  assign n53710 = n53728 ^ n53729;
  assign n53718 = ~n53734;
  assign n53712 = ~n53735;
  assign n53722 = ~n53736;
  assign n52436 = ~n53737;
  assign n53730 = ~n53728;
  assign n53738 = n53750 & n53751;
  assign n52233 = n53701 ^ n52258;
  assign n53662 = n53709 ^ n53710;
  assign n53683 = ~n53716;
  assign n53703 = ~n53701;
  assign n53714 = n53718 & n53719;
  assign n53677 = n53722 & n53723;
  assign n53726 = n53730 & n53731;
  assign n53733 = n53738 & n51226;
  assign n53732 = ~n53738;
  assign n53689 = n53662 & n13481;
  assign n53506 = ~n52233;
  assign n53690 = ~n53662;
  assign n53664 = n53703 & n52285;
  assign n53706 = n53677 & n53692;
  assign n53698 = ~n53714;
  assign n53704 = ~n53677;
  assign n53711 = ~n53726;
  assign n53727 = n53732 & n51192;
  assign n53715 = ~n53733;
  assign n53668 = ~n53689;
  assign n53684 = n53690 & n324;
  assign n53667 = ~n53664;
  assign n53679 = n53698 ^ n53699;
  assign n53697 = n53702 & n53698;
  assign n53700 = n53704 & n53705;
  assign n53694 = ~n53706;
  assign n53691 = n53711 & n53712;
  assign n53717 = n53715 & n53695;
  assign n53708 = ~n53727;
  assign n53665 = n325 ^ n53679;
  assign n53649 = ~n53684;
  assign n53678 = n53691 ^ n53692;
  assign n53682 = ~n53697;
  assign n53676 = ~n53700;
  assign n53693 = ~n53691;
  assign n53713 = n53708 & n53715;
  assign n53707 = ~n53717;
  assign n52199 = n53664 ^ n53665;
  assign n53630 = n53677 ^ n53678;
  assign n53666 = ~n53665;
  assign n53680 = n53682 & n53683;
  assign n53685 = n53693 & n53694;
  assign n53686 = n53707 & n53708;
  assign n53696 = ~n53713;
  assign n53462 = ~n52199;
  assign n53656 = n53630 & n13439;
  assign n53624 = n53666 & n53667;
  assign n53657 = ~n53630;
  assign n53661 = ~n53680;
  assign n53675 = ~n53685;
  assign n53669 = n53686 ^ n51132;
  assign n50173 = n53695 ^ n53696;
  assign n53687 = ~n53686;
  assign n53631 = ~n53656;
  assign n53652 = n53657 & n323;
  assign n53645 = n53661 ^ n53662;
  assign n53663 = n53668 & n53661;
  assign n50084 = n53669 ^ n53670;
  assign n53658 = n53675 & n53676;
  assign n53681 = n53687 & n53688;
  assign n50195 = ~n50173;
  assign n53627 = n324 ^ n53645;
  assign n53612 = ~n53652;
  assign n53654 = n50084 & n51132;
  assign n53653 = n50084 & n52316;
  assign n53639 = n53658 ^ n53643;
  assign n50138 = ~n50084;
  assign n53648 = ~n53663;
  assign n53626 = ~n53658;
  assign n53673 = n50195 & n52355;
  assign n53674 = n50195 & n51226;
  assign n53671 = ~n53681;
  assign n52182 = n53624 ^ n53627;
  assign n53623 = ~n53627;
  assign n53629 = n53648 & n53649;
  assign n53640 = ~n53653;
  assign n52349 = ~n53654;
  assign n53655 = n53671 & n53672;
  assign n53659 = ~n53673;
  assign n52388 = ~n53674;
  assign n53424 = ~n52182;
  assign n53595 = n53623 & n53624;
  assign n53608 = n53629 ^ n53630;
  assign n53566 = n53640 & n53641;
  assign n53632 = ~n53629;
  assign n53633 = n53655 ^ n51081;
  assign n53638 = n53659 & n53660;
  assign n53650 = ~n53655;
  assign n53596 = n323 ^ n53608;
  assign n53598 = ~n53595;
  assign n53618 = n53566 & n53585;
  assign n53628 = n53631 & n53632;
  assign n53620 = ~n53566;
  assign n49999 = n53633 ^ n53634;
  assign n53592 = n53638 ^ n53639;
  assign n53644 = n53638 & n53646;
  assign n53647 = n53650 & n53651;
  assign n53642 = ~n53638;
  assign n52129 = n53595 ^ n53596;
  assign n53597 = ~n53596;
  assign n53586 = ~n53618;
  assign n53614 = n53620 & n53621;
  assign n53615 = n49999 & n52274;
  assign n53616 = n49999 & n51081;
  assign n53619 = n53592 & n322;
  assign n53611 = ~n53628;
  assign n50052 = ~n49999;
  assign n53617 = ~n53592;
  assign n53637 = n53642 & n53643;
  assign n53625 = ~n53644;
  assign n53635 = ~n53647;
  assign n53388 = ~n52129;
  assign n53560 = n53597 & n53598;
  assign n53591 = n53611 & n53612;
  assign n53569 = ~n53614;
  assign n53601 = ~n53615;
  assign n52314 = ~n53616;
  assign n53613 = n53617 & n13411;
  assign n53575 = ~n53619;
  assign n53622 = n53625 & n53626;
  assign n53607 = n53635 & n53636;
  assign n53605 = ~n53637;
  assign n53559 = ~n53560;
  assign n53576 = n53591 ^ n53592;
  assign n53533 = n53601 & n53602;
  assign n53593 = ~n53591;
  assign n53589 = n53607 ^ n51008;
  assign n53594 = ~n53613;
  assign n53604 = ~n53622;
  assign n53609 = ~n53607;
  assign n53561 = n322 ^ n53576;
  assign n53582 = n53533 & n53587;
  assign n49910 = n53589 ^ n53590;
  assign n53588 = n53593 & n53594;
  assign n53581 = ~n53533;
  assign n53603 = n53604 & n53605;
  assign n53606 = n53609 & n53610;
  assign n52094 = n53560 ^ n53561;
  assign n53558 = ~n53561;
  assign n53577 = n49910 & n51008;
  assign n53573 = n53581 & n53555;
  assign n53572 = n49910 & n52226;
  assign n53552 = ~n53582;
  assign n53574 = ~n53588;
  assign n49962 = ~n49910;
  assign n53584 = ~n53603;
  assign n53599 = ~n53606;
  assign n53344 = ~n52094;
  assign n53507 = n53558 & n53559;
  assign n53564 = ~n53572;
  assign n53536 = ~n53573;
  assign n53570 = n53574 & n53575;
  assign n52279 = ~n53577;
  assign n53567 = n53584 ^ n53585;
  assign n53583 = n53586 & n53584;
  assign n53578 = n53599 & n53600;
  assign n53513 = ~n53507;
  assign n53495 = n53564 & n53565;
  assign n53545 = n53566 ^ n53567;
  assign n53532 = ~n53570;
  assign n53557 = n53578 ^ n50940;
  assign n53568 = ~n53583;
  assign n53579 = ~n53578;
  assign n53528 = n53532 ^ n53545;
  assign n53548 = n53495 & n53553;
  assign n53549 = n53545 & n321;
  assign n49826 = n53556 ^ n53557;
  assign n53546 = ~n53495;
  assign n53547 = ~n53545;
  assign n53554 = n53568 & n53569;
  assign n53571 = n53579 & n53580;
  assign n53508 = n321 ^ n53528;
  assign n53542 = n53546 & n53520;
  assign n53541 = n53547 & n13365;
  assign n53522 = ~n53548;
  assign n53538 = n49826 & n52194;
  assign n53511 = ~n53549;
  assign n53543 = n49826 & n50975;
  assign n53534 = n53554 ^ n53555;
  assign n49878 = ~n49826;
  assign n53551 = ~n53554;
  assign n53562 = ~n53571;
  assign n53293 = n53507 ^ n53508;
  assign n53512 = ~n53508;
  assign n53489 = n53533 ^ n53534;
  assign n53529 = ~n53538;
  assign n53531 = ~n53541;
  assign n53493 = ~n53542;
  assign n52230 = ~n53543;
  assign n53550 = n53551 & n53552;
  assign n53544 = n53562 & n53563;
  assign n52056 = ~n53293;
  assign n53447 = n53512 & n53513;
  assign n53518 = n53489 & n320;
  assign n53517 = ~n53489;
  assign n53453 = n53529 & n53530;
  assign n53525 = n53531 & n53532;
  assign n53526 = n53544 ^ n50911;
  assign n53535 = ~n53550;
  assign n53539 = ~n53544;
  assign n53450 = ~n53447;
  assign n53509 = n53453 & n53516;
  assign n53505 = n53517 & n13319;
  assign n53468 = ~n53518;
  assign n53514 = ~n53453;
  assign n53510 = ~n53525;
  assign n49761 = n53526 ^ n53527;
  assign n53519 = n53535 & n53536;
  assign n53537 = n53539 & n53540;
  assign n53486 = ~n53505;
  assign n53501 = n49761 & n52142;
  assign n53503 = n49761 & n53506;
  assign n53479 = ~n53509;
  assign n53488 = n53510 & n53511;
  assign n53500 = n53514 & n53477;
  assign n53502 = n49761 & n50911;
  assign n53496 = n53519 ^ n53520;
  assign n49747 = ~n49761;
  assign n53521 = ~n53519;
  assign n53523 = ~n53537;
  assign n53469 = n53488 ^ n53489;
  assign n53444 = n53495 ^ n53496;
  assign n53494 = n49747 & n52233;
  assign n53487 = ~n53488;
  assign n53456 = ~n53500;
  assign n53490 = ~n53501;
  assign n52207 = ~n53502;
  assign n52235 = ~n53503;
  assign n53515 = n53521 & n53522;
  assign n53504 = n53523 & n53524;
  assign n53448 = n320 ^ n53469;
  assign n53475 = n53444 & n335;
  assign n53481 = n53486 & n53487;
  assign n53480 = ~n53444;
  assign n53410 = n53490 & n53491;
  assign n52250 = ~n53494;
  assign n53483 = n53504 ^ n50861;
  assign n53492 = ~n53515;
  assign n53498 = ~n53504;
  assign n53279 = n53447 ^ n53448;
  assign n53449 = ~n53448;
  assign n53473 = n53410 & n53437;
  assign n53427 = ~n53475;
  assign n53470 = n53480 & n13293;
  assign n53467 = ~n53481;
  assign n53471 = ~n53410;
  assign n49652 = n53482 ^ n53483;
  assign n53476 = n53492 & n53493;
  assign n53497 = n53498 & n53499;
  assign n53270 = ~n53279;
  assign n53403 = n53449 & n53450;
  assign n53443 = n53467 & n53468;
  assign n53451 = ~n53470;
  assign n53459 = n53471 & n53472;
  assign n53460 = n49652 & n52152;
  assign n53433 = ~n53473;
  assign n53461 = n49652 & n52199;
  assign n53463 = n49652 & n50870;
  assign n49711 = ~n49652;
  assign n53454 = n53476 ^ n53477;
  assign n53478 = ~n53476;
  assign n53484 = ~n53497;
  assign n53423 = n53443 ^ n53444;
  assign n53407 = n53453 ^ n53454;
  assign n53413 = ~n53459;
  assign n53452 = ~n53443;
  assign n53445 = ~n53460;
  assign n52201 = ~n53461;
  assign n53457 = n49711 & n53462;
  assign n52167 = ~n53463;
  assign n53474 = n53478 & n53479;
  assign n53464 = n53484 & n53485;
  assign n53404 = n335 ^ n53423;
  assign n53435 = n53407 & n334;
  assign n53369 = n53445 & n53446;
  assign n53442 = n53451 & n53452;
  assign n53434 = ~n53407;
  assign n52219 = ~n53457;
  assign n53438 = n53464 ^ n50859;
  assign n53455 = ~n53474;
  assign n53465 = ~n53464;
  assign n51992 = n53403 ^ n53404;
  assign n53405 = ~n53404;
  assign n53429 = n53369 & n53431;
  assign n53425 = n53434 & n13253;
  assign n53383 = ~n53435;
  assign n53428 = ~n53369;
  assign n49577 = n53438 ^ n53439;
  assign n53426 = ~n53442;
  assign n53436 = n53455 & n53456;
  assign n53458 = n53465 & n53466;
  assign n53212 = ~n51992;
  assign n53359 = n53405 & n53403;
  assign n53419 = n49577 & n53424;
  assign n53408 = ~n53425;
  assign n53406 = n53426 & n53427;
  assign n53417 = n53428 & n53395;
  assign n53391 = ~n53429;
  assign n53418 = n49577 & n52120;
  assign n53420 = n49577 & n50859;
  assign n53411 = n53436 ^ n53437;
  assign n49608 = ~n49577;
  assign n53432 = ~n53436;
  assign n53440 = ~n53458;
  assign n53381 = n53406 ^ n53407;
  assign n53362 = n53410 ^ n53411;
  assign n53409 = ~n53406;
  assign n53368 = ~n53417;
  assign n53401 = ~n53418;
  assign n52165 = ~n53419;
  assign n53414 = n49608 & n52182;
  assign n52135 = ~n53420;
  assign n53430 = n53432 & n53433;
  assign n53416 = n53440 & n53441;
  assign n53360 = n334 ^ n53381;
  assign n53392 = n53362 & n13222;
  assign n53326 = n53401 & n53402;
  assign n53396 = n53408 & n53409;
  assign n53393 = ~n53362;
  assign n52184 = ~n53414;
  assign n53397 = n53416 ^ n50822;
  assign n53412 = ~n53430;
  assign n53421 = ~n53416;
  assign n51959 = n53359 ^ n53360;
  assign n53358 = ~n53360;
  assign n53364 = ~n53392;
  assign n53384 = n53393 & n333;
  assign n53387 = n53326 & n53347;
  assign n53385 = ~n53326;
  assign n53382 = ~n53396;
  assign n49514 = n53397 ^ n53398;
  assign n53394 = n53412 & n53413;
  assign n53415 = n53421 & n53422;
  assign n53171 = ~n51959;
  assign n53318 = n53358 & n53359;
  assign n53376 = n49514 & n50822;
  assign n53361 = n53382 & n53383;
  assign n53341 = ~n53384;
  assign n53373 = n53385 & n53386;
  assign n53374 = n49514 & n52076;
  assign n53352 = ~n53387;
  assign n53375 = n49514 & n53388;
  assign n53370 = n53394 ^ n53395;
  assign n49546 = ~n49514;
  assign n53390 = ~n53394;
  assign n53399 = ~n53415;
  assign n53321 = ~n53318;
  assign n53338 = n53361 ^ n53362;
  assign n53323 = n53369 ^ n53370;
  assign n53371 = n49546 & n52129;
  assign n53363 = ~n53361;
  assign n53329 = ~n53373;
  assign n53365 = ~n53374;
  assign n52131 = ~n53375;
  assign n52091 = ~n53376;
  assign n53389 = n53390 & n53391;
  assign n53377 = n53399 & n53400;
  assign n53319 = n333 ^ n53338;
  assign n53349 = n53323 & n332;
  assign n53353 = n53363 & n53364;
  assign n53348 = ~n53323;
  assign n53282 = n53365 & n53366;
  assign n52149 = ~n53371;
  assign n53354 = n53377 ^ n53378;
  assign n53367 = ~n53389;
  assign n53379 = ~n53377;
  assign n51894 = n53318 ^ n53319;
  assign n53320 = ~n53319;
  assign n53339 = n53348 & n13196;
  assign n53302 = ~n53349;
  assign n53343 = n53282 & n53350;
  assign n53340 = ~n53353;
  assign n53342 = ~n53282;
  assign n49458 = n53354 ^ n50761;
  assign n53355 = n53354 & n50761;
  assign n53346 = n53367 & n53368;
  assign n53372 = n53379 & n53380;
  assign n53131 = ~n51894;
  assign n53271 = n53320 & n53321;
  assign n53325 = ~n53339;
  assign n53322 = n53340 & n53341;
  assign n53333 = n53342 & n53308;
  assign n53310 = ~n53343;
  assign n53334 = n49458 & n53344;
  assign n53327 = n53346 ^ n53347;
  assign n49468 = ~n49458;
  assign n52062 = ~n53355;
  assign n53351 = ~n53346;
  assign n53356 = ~n53372;
  assign n53281 = ~n53271;
  assign n53300 = n53322 ^ n53323;
  assign n53274 = n53326 ^ n53327;
  assign n53330 = n49468 & n51987;
  assign n53324 = ~n53322;
  assign n53285 = ~n53333;
  assign n53331 = n49468 & n52094;
  assign n52116 = ~n53334;
  assign n53345 = n53351 & n53352;
  assign n53335 = n53356 & n53357;
  assign n53272 = n332 ^ n53300;
  assign n53305 = n53274 & n13171;
  assign n53311 = n53324 & n53325;
  assign n53306 = ~n53274;
  assign n53312 = ~n53330;
  assign n52097 = ~n53331;
  assign n53315 = n53335 ^ n50705;
  assign n53328 = ~n53345;
  assign n53336 = ~n53335;
  assign n51855 = n53271 ^ n53272;
  assign n53280 = ~n53272;
  assign n53276 = ~n53305;
  assign n53303 = n53306 & n331;
  assign n53301 = ~n53311;
  assign n53236 = n53312 & n53313;
  assign n49400 = n53314 ^ n53315;
  assign n53307 = n53328 & n53329;
  assign n53332 = n53336 & n53337;
  assign n53082 = ~n51855;
  assign n53226 = n53280 & n53281;
  assign n53273 = n53301 & n53302;
  assign n53249 = ~n53303;
  assign n53291 = n49400 & n51953;
  assign n53292 = n53236 & n53260;
  assign n53294 = n49400 & n52056;
  assign n53295 = n49400 & n50705;
  assign n53283 = n53307 ^ n53308;
  assign n53289 = ~n53236;
  assign n49435 = ~n49400;
  assign n53309 = ~n53307;
  assign n53316 = ~n53332;
  assign n53229 = ~n53226;
  assign n53247 = n53273 ^ n53274;
  assign n53231 = n53282 ^ n53283;
  assign n53275 = ~n53273;
  assign n53286 = n53289 & n53290;
  assign n53277 = ~n53291;
  assign n53261 = ~n53292;
  assign n53287 = n49435 & n53293;
  assign n52058 = ~n53294;
  assign n52020 = ~n53295;
  assign n53304 = n53309 & n53310;
  assign n53296 = n53316 & n53317;
  assign n53227 = n331 ^ n53247;
  assign n53258 = n53231 & n330;
  assign n53267 = n53275 & n53276;
  assign n53257 = ~n53231;
  assign n53196 = n53277 & n53278;
  assign n53239 = ~n53286;
  assign n52082 = ~n53287;
  assign n49337 = n53296 ^ n53297;
  assign n53284 = ~n53304;
  assign n53298 = ~n53296;
  assign n51816 = n53226 ^ n53227;
  assign n53228 = ~n53227;
  assign n53250 = n53257 & n13098;
  assign n53210 = ~n53258;
  assign n53253 = n53196 & n53217;
  assign n53248 = ~n53267;
  assign n53251 = ~n53196;
  assign n53268 = n49337 & n51911;
  assign n53269 = n49337 & n53279;
  assign n53259 = n53284 & n53285;
  assign n49389 = ~n49337;
  assign n53288 = n53298 & n53299;
  assign n53054 = ~n51816;
  assign n53186 = n53228 & n53229;
  assign n53230 = n53248 & n53249;
  assign n53233 = ~n53250;
  assign n53242 = n53251 & n53252;
  assign n53219 = ~n53253;
  assign n53237 = n53259 ^ n53260;
  assign n53254 = ~n53268;
  assign n52018 = ~n53269;
  assign n53263 = n49389 & n53270;
  assign n53264 = n49389 & n50708;
  assign n53262 = ~n53259;
  assign n53265 = ~n53288;
  assign n53189 = ~n53186;
  assign n53208 = n53230 ^ n53231;
  assign n53191 = n53236 ^ n53237;
  assign n53232 = ~n53230;
  assign n53199 = ~n53242;
  assign n53178 = n53254 & n53255;
  assign n53256 = n53261 & n53262;
  assign n52042 = ~n53263;
  assign n51999 = ~n53264;
  assign n53243 = n53265 & n53266;
  assign n53187 = n330 ^ n53208;
  assign n53214 = n53191 & n13075;
  assign n53220 = n53232 & n53233;
  assign n53215 = ~n53191;
  assign n53235 = n53178 & n53240;
  assign n53234 = ~n53178;
  assign n52039 = n52018 & n52042;
  assign n53221 = n53243 ^ n53244;
  assign n53238 = ~n53256;
  assign n53245 = ~n53243;
  assign n51775 = n53186 ^ n53187;
  assign n53188 = ~n53187;
  assign n53193 = ~n53214;
  assign n53211 = n53215 & n329;
  assign n53209 = ~n53220;
  assign n49319 = n50620 ^ n53221;
  assign n53222 = n53234 & n53155;
  assign n53223 = n53221 & n50672;
  assign n53180 = ~n53235;
  assign n53216 = n53238 & n53239;
  assign n53241 = n53245 & n53246;
  assign n53003 = ~n51775;
  assign n53146 = n53188 & n53189;
  assign n53190 = n53209 & n53210;
  assign n53168 = ~n53211;
  assign n53202 = n49319 & n53212;
  assign n53203 = n49319 & n51842;
  assign n53197 = n53216 ^ n53217;
  assign n49348 = ~n49319;
  assign n53157 = ~n53222;
  assign n51942 = ~n53223;
  assign n53218 = ~n53216;
  assign n53224 = ~n53241;
  assign n53166 = n53190 ^ n53191;
  assign n53149 = n53196 ^ n53197;
  assign n53192 = ~n53190;
  assign n51977 = ~n53202;
  assign n53200 = n49348 & n51992;
  assign n53194 = ~n53203;
  assign n53213 = n53218 & n53219;
  assign n53204 = n53224 & n53225;
  assign n53147 = n329 ^ n53166;
  assign n53174 = n53149 & n13017;
  assign n53181 = n53192 & n53193;
  assign n53175 = ~n53149;
  assign n53138 = n53194 & n53195;
  assign n51994 = ~n53200;
  assign n53182 = n53204 ^ n53205;
  assign n53198 = ~n53213;
  assign n53206 = ~n53204;
  assign n51732 = n53146 ^ n53147;
  assign n53109 = n53147 & n53146;
  assign n53150 = ~n53174;
  assign n53169 = n53175 & n328;
  assign n53172 = n53138 & n53176;
  assign n53167 = ~n53181;
  assign n53170 = ~n53138;
  assign n49291 = n50534 ^ n53182;
  assign n53183 = n53182 & n50623;
  assign n53177 = n53198 & n53199;
  assign n53201 = n53206 & n53207;
  assign n52963 = ~n51732;
  assign n53148 = n53167 & n53168;
  assign n53134 = ~n53169;
  assign n53160 = n53170 & n53117;
  assign n53161 = n49291 & n51883;
  assign n53162 = n49291 & n53171;
  assign n53139 = ~n53172;
  assign n53154 = n53177 ^ n53178;
  assign n49280 = ~n49291;
  assign n51899 = ~n53183;
  assign n53179 = ~n53177;
  assign n53184 = ~n53201;
  assign n53129 = n53148 ^ n53149;
  assign n53089 = n53154 ^ n53155;
  assign n53151 = ~n53148;
  assign n53119 = ~n53160;
  assign n53152 = ~n53161;
  assign n51940 = ~n53162;
  assign n53158 = n49280 & n51959;
  assign n53173 = n53179 & n53180;
  assign n53163 = n53184 & n53185;
  assign n53110 = n328 ^ n53129;
  assign n53136 = n53089 & n343;
  assign n53141 = n53150 & n53151;
  assign n53135 = ~n53089;
  assign n53074 = n53152 & n53153;
  assign n51961 = ~n53158;
  assign n53143 = n53163 ^ n50510;
  assign n53156 = ~n53173;
  assign n53164 = ~n53163;
  assign n52920 = n53109 ^ n53110;
  assign n53065 = n53110 & n53109;
  assign n53130 = n53135 & n12996;
  assign n53091 = ~n53136;
  assign n53133 = ~n53141;
  assign n53080 = ~n53074;
  assign n49247 = n53142 ^ n53143;
  assign n53137 = n53156 & n53157;
  assign n53159 = n53164 & n53165;
  assign n52927 = ~n52920;
  assign n53113 = ~n53130;
  assign n53122 = n49247 & n51846;
  assign n53123 = n49247 & n53131;
  assign n53124 = n49247 & n50510;
  assign n53111 = n53133 & n53134;
  assign n53116 = n53137 ^ n53138;
  assign n49236 = ~n49247;
  assign n53140 = ~n53137;
  assign n53144 = ~n53159;
  assign n53088 = n343 ^ n53111;
  assign n53069 = n53116 ^ n53117;
  assign n53112 = ~n53111;
  assign n53120 = n49236 & n51894;
  assign n53114 = ~n53122;
  assign n51897 = ~n53123;
  assign n51862 = ~n53124;
  assign n53132 = n53139 & n53140;
  assign n53125 = n53144 & n53145;
  assign n53066 = n53088 ^ n53089;
  assign n53097 = n53069 & n342;
  assign n53104 = n53112 & n53113;
  assign n53096 = ~n53069;
  assign n53017 = n53114 & n53115;
  assign n51917 = ~n53120;
  assign n53105 = n53125 ^ n53126;
  assign n53118 = ~n53132;
  assign n53127 = ~n53125;
  assign n51666 = n53065 ^ n53066;
  assign n53067 = ~n53066;
  assign n53092 = n53096 & n12940;
  assign n53050 = ~n53097;
  assign n53094 = n53017 & n53098;
  assign n53090 = ~n53104;
  assign n53093 = ~n53017;
  assign n49193 = n50490 ^ n53105;
  assign n53106 = n53105 & n50441;
  assign n53099 = n53118 & n53119;
  assign n53121 = n53127 & n53128;
  assign n52885 = ~n51666;
  assign n53026 = n53067 & n53065;
  assign n53068 = n53090 & n53091;
  assign n53071 = ~n53092;
  assign n53081 = n53093 & n53038;
  assign n53083 = n49193 & n51795;
  assign n53084 = n49193 & n51855;
  assign n53040 = ~n53094;
  assign n53075 = n53099 ^ n53100;
  assign n49223 = ~n49193;
  assign n53103 = n53099 & n53100;
  assign n51814 = ~n53106;
  assign n53101 = ~n53099;
  assign n53107 = ~n53121;
  assign n53048 = n53068 ^ n53069;
  assign n53011 = n53074 ^ n53075;
  assign n53070 = ~n53068;
  assign n53021 = ~n53081;
  assign n53077 = n49223 & n53082;
  assign n53072 = ~n53083;
  assign n51858 = ~n53084;
  assign n53095 = n53101 & n53102;
  assign n53079 = ~n53103;
  assign n53085 = n53107 & n53108;
  assign n53027 = n342 ^ n53048;
  assign n53055 = n53011 & n12900;
  assign n53058 = n53070 & n53071;
  assign n53056 = ~n53011;
  assign n52976 = n53072 & n53073;
  assign n51878 = ~n53077;
  assign n53076 = n53079 & n53080;
  assign n53061 = n53085 ^ n50451;
  assign n53060 = ~n53095;
  assign n53086 = ~n53085;
  assign n51625 = n53026 ^ n53027;
  assign n53028 = ~n53027;
  assign n53030 = ~n53055;
  assign n53051 = n53056 & n341;
  assign n53053 = n52976 & n53057;
  assign n53049 = ~n53058;
  assign n53052 = ~n52976;
  assign n49178 = n53061 ^ n53062;
  assign n53059 = ~n53076;
  assign n53078 = n53086 & n53087;
  assign n52848 = ~n51625;
  assign n52986 = n53028 & n53026;
  assign n53029 = n53049 & n53050;
  assign n53013 = ~n53051;
  assign n53041 = n53052 & n52999;
  assign n53042 = n49178 & n51767;
  assign n53001 = ~n53053;
  assign n53043 = n49178 & n53054;
  assign n53044 = n49178 & n50451;
  assign n49134 = ~n49178;
  assign n53037 = n53059 & n53060;
  assign n53063 = ~n53078;
  assign n52985 = ~n52986;
  assign n53010 = n341 ^ n53029;
  assign n53031 = ~n53029;
  assign n53018 = n53037 ^ n53038;
  assign n52979 = ~n53041;
  assign n53035 = n49134 & n51816;
  assign n53032 = ~n53042;
  assign n51819 = ~n53043;
  assign n51785 = ~n53044;
  assign n53039 = ~n53037;
  assign n53045 = n53063 & n53064;
  assign n52987 = n53010 ^ n53011;
  assign n52989 = n53017 ^ n53018;
  assign n53019 = n53030 & n53031;
  assign n52937 = n53032 & n53033;
  assign n51840 = ~n53035;
  assign n53034 = n53039 & n53040;
  assign n53023 = n53045 ^ n50288;
  assign n53046 = ~n53045;
  assign n51536 = n52986 ^ n52987;
  assign n52984 = ~n52987;
  assign n52997 = n52989 & n340;
  assign n52996 = ~n52989;
  assign n53016 = n52937 & n52957;
  assign n53012 = ~n53019;
  assign n53014 = ~n52937;
  assign n49114 = n53022 ^ n53023;
  assign n53020 = ~n53034;
  assign n53036 = n53046 & n53047;
  assign n52798 = ~n51536;
  assign n52942 = n52984 & n52985;
  assign n52992 = n52996 & n12857;
  assign n52953 = ~n52997;
  assign n52988 = n53012 & n53013;
  assign n53002 = n53014 & n53015;
  assign n52959 = ~n53016;
  assign n53004 = n49114 & n51651;
  assign n53005 = n49114 & n51775;
  assign n53006 = n49114 & n50288;
  assign n49137 = ~n49114;
  assign n52998 = n53020 & n53021;
  assign n53024 = ~n53036;
  assign n52945 = ~n52942;
  assign n52969 = n52988 ^ n52989;
  assign n52974 = ~n52992;
  assign n52975 = ~n52988;
  assign n52977 = n52998 ^ n52999;
  assign n52932 = ~n53002;
  assign n52994 = n49137 & n53003;
  assign n52990 = ~n53004;
  assign n51777 = ~n53005;
  assign n51742 = ~n53006;
  assign n53000 = ~n52998;
  assign n53007 = n53024 & n53025;
  assign n52943 = n340 ^ n52969;
  assign n52973 = n52974 & n52975;
  assign n52934 = n52976 ^ n52977;
  assign n52894 = n52990 & n52991;
  assign n51802 = ~n52994;
  assign n52993 = n53000 & n53001;
  assign n52981 = n53007 ^ n50213;
  assign n53008 = ~n53007;
  assign n51476 = n52942 ^ n52943;
  assign n52944 = ~n52943;
  assign n52955 = n52934 & n339;
  assign n52952 = ~n52973;
  assign n52954 = ~n52934;
  assign n52972 = n52894 & n52914;
  assign n52970 = ~n52894;
  assign n49069 = n52980 ^ n52981;
  assign n52978 = ~n52993;
  assign n52995 = n53008 & n53009;
  assign n52760 = ~n51476;
  assign n52888 = n52944 & n52945;
  assign n52933 = n52952 & n52953;
  assign n52948 = n52954 & n12818;
  assign n52910 = ~n52955;
  assign n52960 = n52970 & n52971;
  assign n52961 = n49069 & n51732;
  assign n52962 = n49069 & n51674;
  assign n52916 = ~n52972;
  assign n52964 = n49069 & n50213;
  assign n49076 = ~n49069;
  assign n52956 = n52978 & n52979;
  assign n52982 = ~n52995;
  assign n52908 = n52933 ^ n52934;
  assign n52935 = ~n52933;
  assign n52936 = ~n52948;
  assign n52938 = n52956 ^ n52957;
  assign n52897 = ~n52960;
  assign n51734 = ~n52961;
  assign n52946 = ~n52962;
  assign n52950 = n49076 & n52963;
  assign n51697 = ~n52964;
  assign n52958 = ~n52956;
  assign n52965 = n52982 & n52983;
  assign n52891 = n339 ^ n52908;
  assign n52929 = n52935 & n52936;
  assign n52893 = n52937 ^ n52938;
  assign n52857 = n52946 & n52947;
  assign n51761 = ~n52950;
  assign n52949 = n52958 & n52959;
  assign n52939 = n52965 ^ n52966;
  assign n52967 = ~n52965;
  assign n51404 = n52888 ^ n52891;
  assign n52887 = ~n52891;
  assign n52911 = n52893 & n12767;
  assign n52909 = ~n52929;
  assign n52912 = ~n52893;
  assign n52928 = n52857 & n52930;
  assign n52926 = ~n52857;
  assign n49027 = n52939 ^ n50126;
  assign n52931 = ~n52949;
  assign n52951 = n52967 & n52968;
  assign n52711 = ~n51404;
  assign n52851 = n52887 & n52888;
  assign n52892 = n52909 & n52910;
  assign n52890 = ~n52911;
  assign n52904 = n52912 & n338;
  assign n52917 = n52926 & n52879;
  assign n52918 = n49027 & n52927;
  assign n52872 = ~n52928;
  assign n52919 = n49027 & n51547;
  assign n52921 = n49027 & n50140;
  assign n49022 = ~n49027;
  assign n52913 = n52931 & n52932;
  assign n52940 = ~n52951;
  assign n52873 = n52892 ^ n52893;
  assign n52889 = ~n52892;
  assign n52875 = ~n52904;
  assign n52895 = n52913 ^ n52914;
  assign n52860 = ~n52917;
  assign n51718 = ~n52918;
  assign n52902 = ~n52919;
  assign n52906 = n49022 & n52920;
  assign n51677 = ~n52921;
  assign n52915 = ~n52913;
  assign n52922 = n52940 & n52941;
  assign n52852 = n338 ^ n52873;
  assign n52886 = n52889 & n52890;
  assign n52854 = n52894 ^ n52895;
  assign n52787 = n52902 & n52903;
  assign n51691 = ~n52906;
  assign n52905 = n52915 & n52916;
  assign n52898 = n52922 ^ n52923;
  assign n52924 = ~n52922;
  assign n51324 = n52851 ^ n52852;
  assign n52813 = n52852 & n52851;
  assign n52876 = n52854 & n12734;
  assign n52874 = ~n52886;
  assign n52877 = ~n52854;
  assign n51715 = n51691 & n51718;
  assign n49004 = n52898 ^ n49964;
  assign n52899 = n52898 & n50141;
  assign n52896 = ~n52905;
  assign n52907 = n52924 & n52925;
  assign n52672 = ~n51324;
  assign n52812 = ~n52813;
  assign n52853 = n52874 & n52875;
  assign n52856 = ~n52876;
  assign n52867 = n52877 & n337;
  assign n52880 = n49004 & n51418;
  assign n52881 = n49004 & n52885;
  assign n48949 = ~n49004;
  assign n52878 = n52896 & n52897;
  assign n51604 = ~n52899;
  assign n52900 = ~n52907;
  assign n52829 = n52853 ^ n52854;
  assign n52855 = ~n52853;
  assign n52831 = ~n52867;
  assign n52858 = n52878 ^ n52879;
  assign n52865 = ~n52880;
  assign n52869 = n48949 & n51666;
  assign n51646 = ~n52881;
  assign n52871 = ~n52878;
  assign n52882 = n52900 & n52901;
  assign n52814 = n337 ^ n52829;
  assign n52849 = n52855 & n52856;
  assign n52816 = n52857 ^ n52858;
  assign n52784 = n52865 & n52866;
  assign n51668 = ~n52869;
  assign n52868 = n52871 & n52872;
  assign n52862 = n52882 ^ n49917;
  assign n52883 = ~n52882;
  assign n52636 = n52813 ^ n52814;
  assign n52811 = ~n52814;
  assign n52833 = n52816 & n336;
  assign n52830 = ~n52849;
  assign n52832 = ~n52816;
  assign n52845 = n52784 & n52850;
  assign n52844 = ~n52784;
  assign n48910 = n52861 ^ n52862;
  assign n52859 = ~n52868;
  assign n52870 = n52883 & n52884;
  assign n52771 = n52811 & n52812;
  assign n52815 = n52830 & n52831;
  assign n52825 = n52832 & n12647;
  assign n52795 = ~n52833;
  assign n52836 = n52844 & n52765;
  assign n52837 = n48910 & n51518;
  assign n52786 = ~n52845;
  assign n52839 = n48910 & n50041;
  assign n52840 = n48910 & n52848;
  assign n48968 = ~n48910;
  assign n52846 = n52859 & n52860;
  assign n52863 = ~n52870;
  assign n52774 = ~n52771;
  assign n52793 = n52815 ^ n52816;
  assign n52809 = ~n52815;
  assign n52810 = ~n52825;
  assign n52767 = ~n52836;
  assign n52823 = ~n52837;
  assign n51545 = ~n52839;
  assign n52827 = n48968 & n51625;
  assign n51598 = ~n52840;
  assign n52838 = n52846 & n52847;
  assign n52834 = ~n52846;
  assign n52841 = n52863 & n52864;
  assign n52772 = n336 ^ n52793;
  assign n52806 = n52809 & n52810;
  assign n52716 = n52823 & n52824;
  assign n51627 = ~n52827;
  assign n52826 = n52834 & n52835;
  assign n52818 = ~n52838;
  assign n52820 = n52841 ^ n49836;
  assign n52842 = ~n52841;
  assign n52750 = n52771 ^ n52772;
  assign n52773 = ~n52772;
  assign n52794 = ~n52806;
  assign n52805 = n52716 & n52807;
  assign n52804 = ~n52716;
  assign n48895 = n52819 ^ n52820;
  assign n52817 = n52818 & n52787;
  assign n52803 = ~n52826;
  assign n52828 = n52842 & n52843;
  assign n48749 = n52750 ^ n50634;
  assign n52751 = n52750 & n50634;
  assign n52657 = n52750 & n50636;
  assign n52726 = n52773 & n52774;
  assign n52775 = n52794 & n52795;
  assign n52796 = n52804 & n52739;
  assign n52743 = ~n52805;
  assign n52797 = n48895 & n51536;
  assign n48928 = ~n48895;
  assign n52802 = ~n52817;
  assign n52808 = n52803 & n52818;
  assign n52821 = ~n52828;
  assign n48751 = ~n48749;
  assign n51637 = ~n52751;
  assign n52752 = n351 ^ n52775;
  assign n52749 = ~n52775;
  assign n52719 = ~n52796;
  assign n52789 = n48928 & n51442;
  assign n52790 = n48928 & n49967;
  assign n51574 = ~n52797;
  assign n52791 = n48928 & n52798;
  assign n52783 = n52802 & n52803;
  assign n52788 = ~n52808;
  assign n52799 = n52821 & n52822;
  assign n52724 = n48751 & n51614;
  assign n52764 = n52783 ^ n52784;
  assign n52753 = n52787 ^ n52788;
  assign n52776 = ~n52789;
  assign n51475 = ~n52790;
  assign n51539 = ~n52791;
  assign n52785 = ~n52783;
  assign n52780 = n52799 ^ n49753;
  assign n52800 = ~n52799;
  assign n52705 = ~n52724;
  assign n52727 = n52752 ^ n52753;
  assign n52701 = n52764 ^ n52765;
  assign n52769 = n52753 & n12617;
  assign n52667 = n52776 & n52777;
  assign n48882 = n52779 ^ n52780;
  assign n52778 = n52785 & n52786;
  assign n52770 = ~n52753;
  assign n52792 = n52800 & n52801;
  assign n52677 = n52705 & n52706;
  assign n52715 = n52726 ^ n52727;
  assign n52645 = n52727 & n52726;
  assign n52737 = n52701 & n350;
  assign n52736 = ~n52701;
  assign n52756 = n48882 & n51230;
  assign n52757 = n52667 & n52693;
  assign n52758 = n48882 & n51476;
  assign n52759 = n48882 & n49753;
  assign n52748 = ~n52769;
  assign n52768 = n52770 & n351;
  assign n52754 = ~n52667;
  assign n48855 = ~n48882;
  assign n52766 = ~n52778;
  assign n52781 = ~n52792;
  assign n52655 = n52677 ^ n52678;
  assign n52679 = ~n52677;
  assign n52708 = n52715 & n50516;
  assign n52707 = ~n52715;
  assign n52648 = ~n52645;
  assign n52728 = n52736 & n12503;
  assign n52683 = ~n52737;
  assign n52744 = n52748 & n52749;
  assign n52745 = n52754 & n52755;
  assign n52740 = ~n52756;
  assign n52695 = ~n52757;
  assign n51479 = ~n52758;
  assign n51403 = ~n52759;
  assign n52746 = n48855 & n52760;
  assign n52738 = n52766 & n52767;
  assign n52730 = ~n52768;
  assign n52761 = n52781 & n52782;
  assign n50816 = n487 ^ n52655;
  assign n52472 = n52655 & n487;
  assign n52542 = n52679 & n52680;
  assign n52698 = n52707 & n50522;
  assign n52659 = ~n52708;
  assign n52709 = ~n52728;
  assign n52717 = n52738 ^ n52739;
  assign n52618 = n52740 & n52741;
  assign n52729 = ~n52744;
  assign n52670 = ~n52745;
  assign n51512 = ~n52746;
  assign n52742 = ~n52738;
  assign n52733 = n52761 ^ n49781;
  assign n52762 = ~n52761;
  assign n50836 = ~n50816;
  assign n52681 = ~n52698;
  assign n52661 = n52716 ^ n52717;
  assign n52722 = n52618 & n52640;
  assign n52725 = n52729 & n52730;
  assign n52720 = ~n52618;
  assign n48815 = n52732 ^ n52733;
  assign n52731 = n52742 & n52743;
  assign n52747 = n52762 & n52763;
  assign n52675 = n52681 & n52657;
  assign n52656 = n52681 & n52659;
  assign n52691 = n52661 & n349;
  assign n52690 = ~n52661;
  assign n52710 = n52720 & n52721;
  assign n52642 = ~n52722;
  assign n52712 = n48815 & n51404;
  assign n52700 = ~n52725;
  assign n48846 = ~n48815;
  assign n52718 = ~n52731;
  assign n52734 = ~n52747;
  assign n48688 = n52656 ^ n52657;
  assign n52658 = ~n52675;
  assign n52684 = n52690 & n12444;
  assign n52631 = ~n52691;
  assign n52676 = n52700 ^ n52701;
  assign n52699 = n52709 & n52700;
  assign n52621 = ~n52710;
  assign n52702 = n48846 & n51167;
  assign n52703 = n48846 & n49675;
  assign n52704 = n48846 & n52711;
  assign n51447 = ~n52712;
  assign n52692 = n52718 & n52719;
  assign n52713 = n52734 & n52735;
  assign n52626 = n48688 & n51514;
  assign n52627 = n48688 & n50522;
  assign n48695 = ~n48688;
  assign n52628 = n52658 & n52659;
  assign n52646 = n350 ^ n52676;
  assign n52662 = ~n52684;
  assign n52668 = n52692 ^ n52693;
  assign n52682 = ~n52699;
  assign n52686 = ~n52702;
  assign n51323 = ~n52703;
  assign n51407 = ~n52704;
  assign n52694 = ~n52692;
  assign n52689 = n52713 ^ n49605;
  assign n52714 = n52713 & n52723;
  assign n52615 = ~n52626;
  assign n51541 = ~n52627;
  assign n52602 = n52628 ^ n50463;
  assign n52601 = ~n52628;
  assign n52603 = n52645 ^ n52646;
  assign n52647 = ~n52646;
  assign n52609 = n52667 ^ n52668;
  assign n52660 = n52682 & n52683;
  assign n52566 = n52686 & n52687;
  assign n48787 = n52688 ^ n52689;
  assign n52685 = n52694 & n52695;
  assign n52696 = ~n52714;
  assign n48654 = n52602 ^ n52603;
  assign n52593 = n52615 & n52616;
  assign n52623 = n52603 & n50463;
  assign n52622 = ~n52603;
  assign n52604 = n52647 & n52648;
  assign n52637 = n52609 & n12352;
  assign n52629 = n52660 ^ n52661;
  assign n52638 = ~n52609;
  assign n52665 = n52566 & n52671;
  assign n52666 = n48787 & n52672;
  assign n52663 = ~n52660;
  assign n52664 = ~n52566;
  assign n48807 = ~n48787;
  assign n52669 = ~n52685;
  assign n52673 = n52696 & n52697;
  assign n52586 = n52593 & n52594;
  assign n48676 = ~n48654;
  assign n52584 = ~n52593;
  assign n52617 = n52622 & n50419;
  assign n52600 = ~n52623;
  assign n52605 = n349 ^ n52629;
  assign n52607 = ~n52604;
  assign n52611 = ~n52637;
  assign n52632 = n52638 & n348;
  assign n52649 = n52662 & n52663;
  assign n52650 = n52664 & n52590;
  assign n52651 = n48807 & n51106;
  assign n52592 = ~n52665;
  assign n52653 = n48807 & n49702;
  assign n51340 = ~n52666;
  assign n52654 = n48807 & n51324;
  assign n52639 = n52669 & n52670;
  assign n48802 = n52673 ^ n52674;
  assign n52570 = n48676 & n51449;
  assign n52571 = n48676 & n50463;
  assign n52574 = n52584 & n52585;
  assign n52565 = ~n52586;
  assign n52595 = n52600 & n52601;
  assign n52529 = n52604 ^ n52605;
  assign n52578 = ~n52617;
  assign n52606 = ~n52605;
  assign n52581 = ~n52632;
  assign n52619 = n52639 ^ n52640;
  assign n52630 = ~n52649;
  assign n52569 = ~n52650;
  assign n52633 = ~n52651;
  assign n52643 = n48802 & n52652;
  assign n51257 = ~n52653;
  assign n52644 = n48802 & n49647;
  assign n51381 = ~n52654;
  assign n52641 = ~n52639;
  assign n49724 = ~n48802;
  assign n52564 = n52565 & n52542;
  assign n52555 = ~n52570;
  assign n51481 = ~n52571;
  assign n52551 = ~n52574;
  assign n52576 = n52529 & n50382;
  assign n52575 = ~n52529;
  assign n52577 = ~n52595;
  assign n52558 = n52606 & n52607;
  assign n52561 = n52618 ^ n52619;
  assign n52608 = n52630 & n52631;
  assign n52523 = n52633 & n52634;
  assign n51301 = n52636 ^ n49724;
  assign n52635 = n52641 & n52642;
  assign n52624 = ~n52643;
  assign n51235 = ~n52644;
  assign n52494 = n52555 & n52556;
  assign n52550 = ~n52564;
  assign n52541 = n52551 & n52565;
  assign n52572 = n52575 & n50339;
  assign n52532 = ~n52576;
  assign n52573 = n52577 & n52578;
  assign n52587 = n52561 & n12313;
  assign n52579 = n52608 ^ n52609;
  assign n52588 = ~n52561;
  assign n52614 = n52523 & n52547;
  assign n52610 = ~n52608;
  assign n52612 = ~n52523;
  assign n52597 = n52624 & n52625;
  assign n52620 = ~n52635;
  assign n52535 = n52494 & n52522;
  assign n52527 = n52541 ^ n52542;
  assign n52533 = ~n52494;
  assign n52543 = n52550 & n52551;
  assign n52557 = ~n52572;
  assign n52553 = ~n52573;
  assign n52559 = n348 ^ n52579;
  assign n52563 = ~n52587;
  assign n52582 = n52588 & n347;
  assign n52480 = n52597 ^ n52598;
  assign n52596 = n52610 & n52611;
  assign n52599 = n52612 & n52613;
  assign n52549 = ~n52614;
  assign n52589 = n52620 & n52621;
  assign n52521 = n52527 & n486;
  assign n52528 = n52533 & n52534;
  assign n52518 = ~n52535;
  assign n52520 = ~n52527;
  assign n52519 = ~n52543;
  assign n52530 = n52553 ^ n50382;
  assign n52552 = n52553 & n52557;
  assign n52483 = n52558 ^ n52559;
  assign n52512 = n52559 & n52558;
  assign n52538 = ~n52582;
  assign n52567 = n52589 ^ n52590;
  assign n52580 = ~n52596;
  assign n52526 = ~n52599;
  assign n52591 = ~n52589;
  assign n52507 = n52518 & n52519;
  assign n52508 = n52520 & n9791;
  assign n52475 = ~n52521;
  assign n52495 = n52519 ^ n52522;
  assign n52497 = ~n52528;
  assign n48644 = n52529 ^ n52530;
  assign n52531 = ~n52552;
  assign n52515 = n52566 ^ n52567;
  assign n52560 = n52580 & n52581;
  assign n52583 = n52591 & n52592;
  assign n52448 = n52494 ^ n52495;
  assign n52496 = ~n52507;
  assign n52498 = ~n52508;
  assign n52503 = n48644 & n51342;
  assign n52504 = n48644 & n50339;
  assign n48624 = ~n48644;
  assign n52509 = n52531 & n52532;
  assign n52545 = n52515 & n346;
  assign n52536 = n52560 ^ n52561;
  assign n52544 = ~n52515;
  assign n52562 = ~n52560;
  assign n52568 = ~n52583;
  assign n52470 = n52448 & n485;
  assign n52469 = ~n52448;
  assign n52473 = n52496 & n52497;
  assign n52482 = n52498 & n52472;
  assign n52471 = n52498 & n52475;
  assign n52485 = ~n52503;
  assign n51409 = ~n52504;
  assign n52484 = n52509 ^ n50251;
  assign n52511 = n52509 & n50295;
  assign n52510 = ~n52509;
  assign n52513 = n347 ^ n52536;
  assign n52539 = n52544 & n12199;
  assign n52492 = ~n52545;
  assign n52554 = n52562 & n52563;
  assign n52546 = n52568 & n52569;
  assign n52458 = n52469 & n9753;
  assign n52427 = ~n52470;
  assign n52442 = n52471 ^ n52472;
  assign n52444 = n52473 ^ n52460;
  assign n52450 = ~n52473;
  assign n52474 = ~n52482;
  assign n48588 = n52483 ^ n52484;
  assign n52443 = n52485 & n52486;
  assign n52505 = n52510 & n50251;
  assign n52499 = ~n52511;
  assign n52428 = n52512 ^ n52513;
  assign n52462 = n52513 & n52512;
  assign n52517 = ~n52539;
  assign n52524 = n52546 ^ n52547;
  assign n52537 = ~n52554;
  assign n52548 = ~n52546;
  assign n50789 = n52442 ^ n50816;
  assign n52407 = n52443 ^ n52444;
  assign n52403 = n52442 & n50816;
  assign n52445 = ~n52458;
  assign n52447 = n52474 & n52475;
  assign n52461 = n52443 & n52476;
  assign n48609 = ~n48588;
  assign n52459 = ~n52443;
  assign n52487 = n52499 & n52483;
  assign n52489 = n52428 & n50195;
  assign n52478 = ~n52505;
  assign n52488 = ~n52428;
  assign n52466 = n52523 ^ n52524;
  assign n52514 = n52537 & n52538;
  assign n52540 = n52548 & n52549;
  assign n52424 = n52407 & n484;
  assign n52035 = ~n50789;
  assign n52423 = ~n52407;
  assign n52425 = n52447 ^ n52448;
  assign n52446 = ~n52447;
  assign n52454 = n48609 & n51292;
  assign n52455 = n48609 & n50295;
  assign n52456 = n52459 & n52460;
  assign n52449 = ~n52461;
  assign n52477 = ~n52487;
  assign n52481 = n52488 & n50173;
  assign n52433 = ~n52489;
  assign n52500 = n52466 & n12147;
  assign n52490 = n52514 ^ n52515;
  assign n52501 = ~n52466;
  assign n52516 = ~n52514;
  assign n52525 = ~n52540;
  assign n52418 = n52423 & n9721;
  assign n52380 = ~n52424;
  assign n52404 = n485 ^ n52425;
  assign n52434 = n52445 & n52446;
  assign n52437 = n52449 & n52450;
  assign n52435 = ~n52454;
  assign n51332 = ~n52455;
  assign n52431 = ~n52456;
  assign n52451 = n52477 & n52478;
  assign n52453 = ~n52481;
  assign n52463 = n346 ^ n52490;
  assign n52468 = ~n52500;
  assign n52493 = n52501 & n345;
  assign n52506 = n52516 & n52517;
  assign n52502 = n52525 & n52526;
  assign n50774 = n52403 ^ n52404;
  assign n52401 = ~n52418;
  assign n52405 = ~n52404;
  assign n52426 = ~n52434;
  assign n52381 = n52435 & n52436;
  assign n52430 = ~n52437;
  assign n52429 = n52451 ^ n50173;
  assign n52452 = ~n52451;
  assign n52384 = n52462 ^ n52463;
  assign n52464 = ~n52463;
  assign n52441 = ~n52493;
  assign n52479 = n344 ^ n52502;
  assign n52491 = ~n52506;
  assign n52016 = ~n50774;
  assign n52366 = n52405 & n52403;
  assign n52406 = n52426 & n52427;
  assign n48553 = n52428 ^ n52429;
  assign n52410 = n52430 & n52431;
  assign n52390 = ~n52381;
  assign n52438 = n52452 & n52453;
  assign n52392 = ~n52384;
  assign n52419 = n52464 & n52462;
  assign n52422 = n52479 ^ n52480;
  assign n52465 = n52491 & n52492;
  assign n52378 = n52406 ^ n52407;
  assign n52382 = n52410 ^ n52411;
  assign n52408 = n48553 & n51192;
  assign n52409 = n48553 & n50173;
  assign n52413 = n52410 & n52417;
  assign n52402 = ~n52406;
  assign n48577 = ~n48553;
  assign n52412 = ~n52410;
  assign n52432 = ~n52438;
  assign n52439 = n52465 ^ n52466;
  assign n52467 = ~n52465;
  assign n52367 = n484 ^ n52378;
  assign n52353 = n52381 ^ n52382;
  assign n52394 = n52401 & n52402;
  assign n52387 = ~n52408;
  assign n51248 = ~n52409;
  assign n52395 = n52412 & n52411;
  assign n52389 = ~n52413;
  assign n52414 = n52432 & n52433;
  assign n52420 = n345 ^ n52439;
  assign n52457 = n52467 & n52468;
  assign n50733 = n52366 ^ n52367;
  assign n52368 = ~n52367;
  assign n52337 = n52387 & n52388;
  assign n52385 = n52389 & n52390;
  assign n52379 = ~n52394;
  assign n52372 = ~n52395;
  assign n52383 = n52414 ^ n50138;
  assign n52416 = n52414 & n50138;
  assign n52415 = ~n52414;
  assign n52340 = n52419 ^ n52420;
  assign n52399 = n52420 & n52419;
  assign n52440 = ~n52457;
  assign n51963 = ~n50733;
  assign n52332 = n52368 & n52366;
  assign n52369 = n52379 & n52380;
  assign n52345 = ~n52337;
  assign n48514 = n52383 ^ n52384;
  assign n52371 = ~n52385;
  assign n52396 = n52415 & n50084;
  assign n52398 = n52340 & n49999;
  assign n52391 = ~n52416;
  assign n52397 = ~n52340;
  assign n52421 = n52440 & n52441;
  assign n52346 = n52369 ^ n52353;
  assign n52370 = n52369 & n9697;
  assign n52354 = n52371 & n52372;
  assign n52365 = ~n52369;
  assign n48516 = ~n48514;
  assign n52386 = n52391 & n52392;
  assign n52374 = ~n52396;
  assign n52393 = n52397 & n50052;
  assign n52343 = ~n52398;
  assign n52400 = n52421 ^ n52422;
  assign n52333 = n483 ^ n52346;
  assign n52338 = n52354 ^ n52355;
  assign n52357 = n52354 & n52362;
  assign n52361 = n52365 & n483;
  assign n52352 = ~n52370;
  assign n52363 = n48516 & n51151;
  assign n52364 = n48516 & n50138;
  assign n52356 = ~n52354;
  assign n52373 = ~n52386;
  assign n52360 = ~n52393;
  assign n52307 = n52399 ^ n52400;
  assign n50677 = n52332 ^ n52333;
  assign n52312 = n52337 ^ n52338;
  assign n52334 = ~n52333;
  assign n52347 = n52352 & n52353;
  assign n52350 = n52356 & n52355;
  assign n52344 = ~n52357;
  assign n52336 = ~n52361;
  assign n52348 = ~n52363;
  assign n51179 = ~n52364;
  assign n52358 = n52373 & n52374;
  assign n52377 = n52307 & n49962;
  assign n52376 = ~n52307;
  assign n51923 = ~n50677;
  assign n52291 = n52334 & n52332;
  assign n52341 = n52344 & n52345;
  assign n52335 = ~n52347;
  assign n52298 = n52348 & n52349;
  assign n52331 = ~n52350;
  assign n52339 = n52358 ^ n50052;
  assign n52359 = ~n52358;
  assign n52375 = n52376 & n49910;
  assign n52329 = ~n52377;
  assign n52323 = n52335 & n52336;
  assign n48463 = n52339 ^ n52340;
  assign n52330 = ~n52341;
  assign n52303 = ~n52298;
  assign n52351 = n52359 & n52360;
  assign n52310 = ~n52375;
  assign n52304 = n52323 ^ n52312;
  assign n52324 = n52323 & n9663;
  assign n52325 = n48463 & n51073;
  assign n52326 = n48463 & n50052;
  assign n52315 = n52330 & n52331;
  assign n52322 = ~n52323;
  assign n48496 = ~n48463;
  assign n52342 = ~n52351;
  assign n52292 = n482 ^ n52304;
  assign n52299 = n52315 ^ n52316;
  assign n52318 = n52315 & n52320;
  assign n52319 = n52322 & n482;
  assign n52311 = ~n52324;
  assign n52313 = ~n52325;
  assign n51110 = ~n52326;
  assign n52317 = ~n52315;
  assign n52327 = n52342 & n52343;
  assign n50655 = n52291 ^ n52292;
  assign n52270 = n52298 ^ n52299;
  assign n52293 = ~n52292;
  assign n52305 = n52311 & n52312;
  assign n52253 = n52313 & n52314;
  assign n52308 = n52317 & n52316;
  assign n52302 = ~n52318;
  assign n52297 = ~n52319;
  assign n52306 = n52327 ^ n49962;
  assign n52328 = ~n52327;
  assign n51885 = ~n50655;
  assign n52245 = n52293 & n52291;
  assign n52300 = n52302 & n52303;
  assign n52296 = ~n52305;
  assign n52260 = ~n52253;
  assign n48419 = n52306 ^ n52307;
  assign n52287 = ~n52308;
  assign n52321 = n52328 & n52329;
  assign n52282 = n52296 & n52297;
  assign n52286 = ~n52300;
  assign n48455 = ~n48419;
  assign n52309 = ~n52321;
  assign n52263 = n52282 ^ n52270;
  assign n52271 = n52286 & n52287;
  assign n52284 = n52282 & n9619;
  assign n52283 = ~n52282;
  assign n52288 = n48455 & n51000;
  assign n52289 = n48455 & n49962;
  assign n52301 = n52309 & n52310;
  assign n52246 = n481 ^ n52263;
  assign n52254 = n52271 ^ n52272;
  assign n52275 = n52271 & n52272;
  assign n52277 = n52283 & n481;
  assign n52269 = ~n52284;
  assign n52273 = ~n52271;
  assign n52278 = ~n52288;
  assign n51046 = ~n52289;
  assign n52295 = n52301 & n49878;
  assign n52294 = ~n52301;
  assign n50578 = n52245 ^ n52246;
  assign n52237 = n52253 ^ n52254;
  assign n52247 = ~n52246;
  assign n52264 = n52269 & n52270;
  assign n52266 = n52273 & n52274;
  assign n52259 = ~n52275;
  assign n52252 = ~n52277;
  assign n52210 = n52278 & n52279;
  assign n52290 = n52294 & n49826;
  assign n52281 = ~n52295;
  assign n51837 = ~n50578;
  assign n52202 = n52247 & n52245;
  assign n52224 = ~n52237;
  assign n52255 = n52259 & n52260;
  assign n52251 = ~n52264;
  assign n52262 = n52210 & n52265;
  assign n52243 = ~n52266;
  assign n52261 = ~n52210;
  assign n52280 = n52281 & n52285;
  assign n52268 = ~n52290;
  assign n52205 = ~n52202;
  assign n52236 = n52251 & n52252;
  assign n52242 = ~n52255;
  assign n52256 = n52261 & n52226;
  assign n52228 = ~n52262;
  assign n52267 = ~n52280;
  assign n52276 = n52268 & n52281;
  assign n52220 = n52236 ^ n52237;
  assign n52239 = n52236 & n9577;
  assign n52225 = n52242 & n52243;
  assign n52238 = ~n52236;
  assign n52213 = ~n52256;
  assign n52248 = n52267 & n52268;
  assign n52257 = ~n52276;
  assign n52203 = n480 ^ n52220;
  assign n52211 = n52225 ^ n52226;
  assign n52231 = n52238 & n480;
  assign n52223 = ~n52239;
  assign n52227 = ~n52225;
  assign n52232 = n52248 ^ n49761;
  assign n48381 = n52257 ^ n52258;
  assign n52249 = ~n52248;
  assign n50525 = n52202 ^ n52203;
  assign n52175 = n52210 ^ n52211;
  assign n52204 = ~n52203;
  assign n52221 = n52223 & n52224;
  assign n52222 = n52227 & n52228;
  assign n52209 = ~n52231;
  assign n48341 = n52232 ^ n52233;
  assign n52240 = n48381 & n50940;
  assign n52241 = n48381 & n49878;
  assign n52244 = n52249 & n52250;
  assign n48413 = ~n48381;
  assign n51807 = ~n50525;
  assign n52156 = n52204 & n52205;
  assign n52208 = ~n52221;
  assign n52215 = n48341 & n50904;
  assign n52216 = n48341 & n49747;
  assign n52212 = ~n52222;
  assign n48372 = ~n48341;
  assign n52229 = ~n52240;
  assign n50995 = ~n52241;
  assign n52234 = ~n52244;
  assign n52155 = ~n52156;
  assign n52189 = n52208 & n52209;
  assign n52193 = n52212 & n52213;
  assign n52206 = ~n52215;
  assign n50949 = ~n52216;
  assign n52170 = n52229 & n52230;
  assign n52217 = n52234 & n52235;
  assign n52168 = n52189 ^ n52175;
  assign n52171 = n52193 ^ n52194;
  assign n52191 = n52189 & n9544;
  assign n52196 = n52193 & n52197;
  assign n52190 = ~n52189;
  assign n52124 = n52206 & n52207;
  assign n52195 = ~n52193;
  assign n52198 = n52217 ^ n49711;
  assign n52177 = ~n52170;
  assign n52218 = ~n52217;
  assign n52157 = n495 ^ n52168;
  assign n52133 = n52170 ^ n52171;
  assign n52185 = n52190 & n495;
  assign n52174 = ~n52191;
  assign n52187 = n52124 & n52192;
  assign n52188 = n52195 & n52194;
  assign n52176 = ~n52196;
  assign n52186 = ~n52124;
  assign n48300 = n52198 ^ n52199;
  assign n52214 = n52218 & n52219;
  assign n50460 = n52156 ^ n52157;
  assign n52154 = ~n52157;
  assign n52169 = n52174 & n52175;
  assign n52172 = n52176 & n52177;
  assign n52159 = ~n52185;
  assign n52178 = n52186 & n52142;
  assign n52179 = n48300 & n50861;
  assign n52144 = ~n52187;
  assign n52180 = n48300 & n49711;
  assign n52161 = ~n52188;
  assign n48331 = ~n48300;
  assign n52200 = ~n52214;
  assign n51757 = ~n50460;
  assign n52101 = n52154 & n52155;
  assign n52158 = ~n52169;
  assign n52160 = ~n52172;
  assign n52127 = ~n52178;
  assign n52166 = ~n52179;
  assign n50901 = ~n52180;
  assign n52181 = n52200 & n52201;
  assign n52104 = ~n52101;
  assign n52150 = n52158 & n52159;
  assign n52141 = n52160 & n52161;
  assign n52088 = n52166 & n52167;
  assign n52162 = n52181 ^ n52182;
  assign n52183 = ~n52181;
  assign n52125 = n52141 ^ n52142;
  assign n52140 = n52150 & n9510;
  assign n52136 = ~n52150;
  assign n52153 = n52088 & n52110;
  assign n52143 = ~n52141;
  assign n52151 = ~n52088;
  assign n48259 = n49577 ^ n52162;
  assign n52163 = n52162 & n49608;
  assign n52173 = n52183 & n52184;
  assign n52086 = n52124 ^ n52125;
  assign n52122 = n52136 ^ n52133;
  assign n52139 = n52136 & n494;
  assign n52132 = ~n52140;
  assign n52137 = n52143 & n52144;
  assign n52145 = n52151 & n52152;
  assign n52146 = n48259 & n50819;
  assign n52112 = ~n52153;
  assign n48291 = ~n48259;
  assign n50872 = ~n52163;
  assign n52164 = ~n52173;
  assign n52102 = n494 ^ n52122;
  assign n52123 = n52132 & n52133;
  assign n52126 = ~n52137;
  assign n52118 = ~n52139;
  assign n52093 = ~n52145;
  assign n52134 = ~n52146;
  assign n52147 = n52164 & n52165;
  assign n51711 = n52101 ^ n52102;
  assign n52103 = ~n52102;
  assign n52117 = ~n52123;
  assign n52109 = n52126 & n52127;
  assign n52051 = n52134 & n52135;
  assign n52128 = n52147 ^ n49546;
  assign n52148 = ~n52147;
  assign n50390 = ~n51711;
  assign n52059 = n52103 & n52104;
  assign n52089 = n52109 ^ n52110;
  assign n52098 = n52117 & n52118;
  assign n52121 = n52051 & n52072;
  assign n52111 = ~n52109;
  assign n52119 = ~n52051;
  assign n48218 = n52128 ^ n52129;
  assign n52138 = n52148 & n52149;
  assign n52047 = n52088 ^ n52089;
  assign n52083 = n52098 ^ n52086;
  assign n52100 = n52098 & n9459;
  assign n52099 = ~n52098;
  assign n52105 = n52111 & n52112;
  assign n52113 = n52119 & n52120;
  assign n52074 = ~n52121;
  assign n48242 = ~n48218;
  assign n52130 = ~n52138;
  assign n52060 = n493 ^ n52083;
  assign n52069 = n52047 & n9421;
  assign n52070 = ~n52047;
  assign n52087 = n52099 & n493;
  assign n52085 = ~n52100;
  assign n52092 = ~n52105;
  assign n52054 = ~n52113;
  assign n52106 = n48242 & n50785;
  assign n52107 = n48242 & n49546;
  assign n52114 = n52130 & n52131;
  assign n51700 = n52059 ^ n52060;
  assign n52002 = n52060 & n52059;
  assign n52049 = ~n52069;
  assign n52065 = n52070 & n492;
  assign n52084 = n52085 & n52086;
  assign n52064 = ~n52087;
  assign n52071 = n52092 & n52093;
  assign n52090 = ~n52106;
  assign n50828 = ~n52107;
  assign n52095 = n52114 ^ n49458;
  assign n52115 = ~n52114;
  assign n51687 = ~n51700;
  assign n52009 = ~n52002;
  assign n52022 = ~n52065;
  assign n52052 = n52071 ^ n52072;
  assign n52063 = ~n52084;
  assign n52073 = ~n52071;
  assign n52010 = n52090 & n52091;
  assign n48174 = n52094 ^ n52095;
  assign n52108 = n52115 & n52116;
  assign n52005 = n52051 ^ n52052;
  assign n52046 = n52063 & n52064;
  assign n52066 = n52073 & n52074;
  assign n52077 = n48174 & n50752;
  assign n52078 = n52010 & n52031;
  assign n52079 = n48174 & n49458;
  assign n52075 = ~n52010;
  assign n48210 = ~n48174;
  assign n52096 = ~n52108;
  assign n52028 = n52005 & n9407;
  assign n52023 = n52046 ^ n52047;
  assign n52029 = ~n52005;
  assign n52048 = ~n52046;
  assign n52053 = ~n52066;
  assign n52067 = n52075 & n52076;
  assign n52061 = ~n52077;
  assign n52033 = ~n52078;
  assign n50781 = ~n52079;
  assign n52080 = n52096 & n52097;
  assign n52003 = n492 ^ n52023;
  assign n52001 = ~n52028;
  assign n52024 = n52029 & n491;
  assign n52043 = n52048 & n52049;
  assign n52030 = n52053 & n52054;
  assign n51970 = n52061 & n52062;
  assign n52013 = ~n52067;
  assign n52055 = n52080 ^ n49435;
  assign n52081 = ~n52080;
  assign n50271 = n52002 ^ n52003;
  assign n51964 = n52003 & n52009;
  assign n51980 = ~n52024;
  assign n52011 = n52030 ^ n52031;
  assign n52021 = ~n52043;
  assign n52045 = n51970 & n52050;
  assign n52032 = ~n52030;
  assign n52044 = ~n51970;
  assign n48132 = n52055 ^ n52056;
  assign n52068 = n52081 & n52082;
  assign n51632 = ~n50271;
  assign n51967 = n52010 ^ n52011;
  assign n52004 = n52021 & n52022;
  assign n52025 = n52032 & n52033;
  assign n52034 = n52044 & n51987;
  assign n51989 = ~n52045;
  assign n52036 = n48132 & n50741;
  assign n52037 = n48132 & n50789;
  assign n52038 = n48132 & n49435;
  assign n48166 = ~n48132;
  assign n52057 = ~n52068;
  assign n51985 = n51967 & n9340;
  assign n51978 = n52004 ^ n52005;
  assign n51984 = ~n51967;
  assign n52000 = ~n52004;
  assign n52012 = ~n52025;
  assign n51973 = ~n52034;
  assign n52026 = n48166 & n52035;
  assign n52019 = ~n52036;
  assign n50791 = ~n52037;
  assign n50763 = ~n52038;
  assign n52040 = n52057 & n52058;
  assign n51965 = n491 ^ n51978;
  assign n51981 = n51984 & n490;
  assign n51969 = ~n51985;
  assign n51995 = n52000 & n52001;
  assign n51986 = n52012 & n52013;
  assign n51933 = n52019 & n52020;
  assign n50805 = ~n52026;
  assign n48070 = n52039 ^ n52040;
  assign n52041 = ~n52040;
  assign n50191 = n51964 ^ n51965;
  assign n51924 = n51965 & n51964;
  assign n51945 = ~n51981;
  assign n51971 = n51986 ^ n51987;
  assign n51979 = ~n51995;
  assign n51997 = n51933 & n52006;
  assign n51988 = ~n51986;
  assign n51996 = ~n51933;
  assign n52014 = n48070 & n50774;
  assign n52015 = n48070 & n50641;
  assign n48122 = ~n48070;
  assign n52027 = n52041 & n52042;
  assign n51571 = ~n50191;
  assign n51927 = ~n51924;
  assign n51929 = n51970 ^ n51971;
  assign n51966 = n51979 & n51980;
  assign n51982 = n51988 & n51989;
  assign n51990 = n51996 & n51953;
  assign n51955 = ~n51997;
  assign n50776 = ~n52014;
  assign n51998 = ~n52015;
  assign n52007 = n48122 & n52016;
  assign n52008 = n48122 & n49389;
  assign n52017 = ~n52027;
  assign n51951 = n51929 & n489;
  assign n51943 = n51966 ^ n51967;
  assign n51950 = ~n51929;
  assign n51968 = ~n51966;
  assign n51972 = ~n51982;
  assign n51936 = ~n51990;
  assign n51871 = n51998 & n51999;
  assign n50758 = ~n52007;
  assign n50715 = ~n52008;
  assign n51991 = n52017 & n52018;
  assign n51925 = n490 ^ n51943;
  assign n51946 = n51950 & n9304;
  assign n51901 = ~n51951;
  assign n51962 = n51968 & n51969;
  assign n51952 = n51972 & n51973;
  assign n51974 = n51991 ^ n51992;
  assign n51993 = ~n51991;
  assign n51521 = n51924 ^ n51925;
  assign n51926 = ~n51925;
  assign n51931 = ~n51946;
  assign n51934 = n51952 ^ n51953;
  assign n51944 = ~n51962;
  assign n51954 = ~n51952;
  assign n48032 = n51974 ^ n49319;
  assign n51975 = n51974 & n49348;
  assign n51983 = n51993 & n51994;
  assign n50062 = ~n51521;
  assign n51886 = n51926 & n51927;
  assign n51889 = n51933 ^ n51934;
  assign n51928 = n51944 & n51945;
  assign n51947 = n51954 & n51955;
  assign n51956 = n48032 & n50620;
  assign n51957 = n48032 & n51963;
  assign n48084 = ~n48032;
  assign n50675 = ~n51975;
  assign n51976 = ~n51983;
  assign n51908 = n51889 & n488;
  assign n51902 = n51928 ^ n51929;
  assign n51907 = ~n51889;
  assign n51930 = ~n51928;
  assign n51935 = ~n51947;
  assign n51941 = ~n51956;
  assign n51948 = n48084 & n50733;
  assign n50719 = ~n51957;
  assign n51958 = n51976 & n51977;
  assign n51887 = n489 ^ n51902;
  assign n51903 = n51907 & n9262;
  assign n51867 = ~n51908;
  assign n51918 = n51930 & n51931;
  assign n51920 = n51935 & n51936;
  assign n51860 = n51941 & n51942;
  assign n50735 = ~n51948;
  assign n51937 = n51958 ^ n51959;
  assign n51960 = ~n51958;
  assign n51457 = n51886 ^ n51887;
  assign n51848 = n51887 & n51886;
  assign n51891 = ~n51903;
  assign n51900 = ~n51918;
  assign n51913 = n51920 & n51921;
  assign n51922 = n51860 & n51932;
  assign n51910 = ~n51920;
  assign n51919 = ~n51860;
  assign n48012 = n51937 ^ n49291;
  assign n51938 = n51937 & n49280;
  assign n51949 = n51960 & n51961;
  assign n49974 = ~n51457;
  assign n51888 = n51900 & n51901;
  assign n51904 = n51910 & n51911;
  assign n51893 = ~n51913;
  assign n51909 = n51919 & n51842;
  assign n51912 = n48012 & n50534;
  assign n51864 = ~n51922;
  assign n51914 = n48012 & n51923;
  assign n48021 = ~n48012;
  assign n50626 = ~n51938;
  assign n51939 = ~n51949;
  assign n51865 = n51888 ^ n51889;
  assign n51890 = ~n51888;
  assign n51892 = n51893 & n51871;
  assign n51881 = ~n51904;
  assign n51844 = ~n51909;
  assign n51898 = ~n51912;
  assign n50679 = ~n51914;
  assign n51905 = n48021 & n50677;
  assign n51915 = n51939 & n51940;
  assign n51849 = n488 ^ n51865;
  assign n51879 = n51890 & n51891;
  assign n51880 = ~n51892;
  assign n51870 = n51881 & n51893;
  assign n51803 = n51898 & n51899;
  assign n50699 = ~n51905;
  assign n51895 = n51915 ^ n49247;
  assign n51916 = ~n51915;
  assign n51380 = n51848 ^ n51849;
  assign n51808 = n51849 & n51848;
  assign n51827 = n51870 ^ n51871;
  assign n51866 = ~n51879;
  assign n51859 = n51880 & n51881;
  assign n51884 = n51803 & n51823;
  assign n51882 = ~n51803;
  assign n47958 = n51894 ^ n51895;
  assign n51906 = n51916 & n51917;
  assign n49887 = ~n51380;
  assign n51853 = n51827 & n503;
  assign n51841 = n51859 ^ n51860;
  assign n51850 = n51866 & n51867;
  assign n51852 = ~n51827;
  assign n51863 = ~n51859;
  assign n51872 = n51882 & n51883;
  assign n51825 = ~n51884;
  assign n51873 = n47958 & n50571;
  assign n51874 = n47958 & n51885;
  assign n51875 = n47958 & n49236;
  assign n48003 = ~n47958;
  assign n51896 = ~n51906;
  assign n51791 = n51841 ^ n51842;
  assign n51826 = n503 ^ n51850;
  assign n51851 = n51852 & n9219;
  assign n51811 = ~n51853;
  assign n51834 = ~n51850;
  assign n51854 = n51863 & n51864;
  assign n51806 = ~n51872;
  assign n51868 = n48003 & n50655;
  assign n51861 = ~n51873;
  assign n50630 = ~n51874;
  assign n50593 = ~n51875;
  assign n51876 = n51896 & n51897;
  assign n51809 = n51826 ^ n51827;
  assign n51821 = n51791 & n502;
  assign n51820 = ~n51791;
  assign n51833 = ~n51851;
  assign n51843 = ~n51854;
  assign n51762 = n51861 & n51862;
  assign n50657 = ~n51868;
  assign n51856 = n51876 ^ n49193;
  assign n51877 = ~n51876;
  assign n49805 = n51808 ^ n51809;
  assign n51746 = n51809 & n51808;
  assign n51812 = n51820 & n9190;
  assign n51770 = ~n51821;
  assign n51828 = n51833 & n51834;
  assign n51822 = n51843 & n51844;
  assign n51847 = n51762 & n51781;
  assign n51845 = ~n51762;
  assign n47918 = n51855 ^ n51856;
  assign n51869 = n51877 & n51878;
  assign n51289 = ~n49805;
  assign n51749 = ~n51746;
  assign n51792 = ~n51812;
  assign n51804 = n51822 ^ n51823;
  assign n51810 = ~n51828;
  assign n51824 = ~n51822;
  assign n51835 = n51845 & n51846;
  assign n51783 = ~n51847;
  assign n51836 = n47918 & n50578;
  assign n47949 = ~n47918;
  assign n51857 = ~n51869;
  assign n51751 = n51803 ^ n51804;
  assign n51790 = n51810 & n51811;
  assign n51815 = n51824 & n51825;
  assign n51765 = ~n51835;
  assign n51829 = n47949 & n50490;
  assign n50607 = ~n51836;
  assign n51830 = n47949 & n51837;
  assign n51831 = n47949 & n49223;
  assign n51838 = n51857 & n51858;
  assign n51778 = n51751 & n9138;
  assign n51771 = n51790 ^ n51791;
  assign n51779 = ~n51751;
  assign n51793 = ~n51790;
  assign n51805 = ~n51815;
  assign n51813 = ~n51829;
  assign n50581 = ~n51830;
  assign n50524 = ~n51831;
  assign n51817 = n51838 ^ n49178;
  assign n51839 = ~n51838;
  assign n51747 = n502 ^ n51771;
  assign n51753 = ~n51778;
  assign n51772 = n51779 & n501;
  assign n51786 = n51792 & n51793;
  assign n51780 = n51805 & n51806;
  assign n51719 = n51813 & n51814;
  assign n47878 = n51816 ^ n51817;
  assign n51832 = n51839 & n51840;
  assign n51258 = n51746 ^ n51747;
  assign n51748 = ~n51747;
  assign n51727 = ~n51772;
  assign n51763 = n51780 ^ n51781;
  assign n51769 = ~n51786;
  assign n51782 = ~n51780;
  assign n51796 = n47878 & n50369;
  assign n51797 = n51719 & n51738;
  assign n51798 = n47878 & n51807;
  assign n51799 = n47878 & n49134;
  assign n51794 = ~n51719;
  assign n47923 = ~n47878;
  assign n51818 = ~n51832;
  assign n51704 = n51748 & n51749;
  assign n51707 = n51762 ^ n51763;
  assign n51750 = n51769 & n51770;
  assign n51773 = n51782 & n51783;
  assign n51787 = n51794 & n51795;
  assign n51784 = ~n51796;
  assign n51740 = ~n51797;
  assign n50528 = ~n51798;
  assign n51788 = n47923 & n50525;
  assign n50473 = ~n51799;
  assign n51800 = n51818 & n51819;
  assign n51735 = n51707 & n9098;
  assign n51728 = n51750 ^ n51751;
  assign n51736 = ~n51707;
  assign n51752 = ~n51750;
  assign n51764 = ~n51773;
  assign n51669 = n51784 & n51785;
  assign n51722 = ~n51787;
  assign n50554 = ~n51788;
  assign n51774 = n51800 ^ n49137;
  assign n51801 = ~n51800;
  assign n51705 = n501 ^ n51728;
  assign n51709 = ~n51735;
  assign n51729 = n51736 & n500;
  assign n51743 = n51752 & n51753;
  assign n51737 = n51764 & n51765;
  assign n51768 = n51669 & n51695;
  assign n51766 = ~n51669;
  assign n47836 = n51774 ^ n51775;
  assign n51789 = n51801 & n51802;
  assign n51681 = n51704 ^ n51705;
  assign n51658 = n51705 & n51704;
  assign n51680 = ~n51729;
  assign n51720 = n51737 ^ n51738;
  assign n51726 = ~n51743;
  assign n51739 = ~n51737;
  assign n51754 = n51766 & n51767;
  assign n51755 = n47836 & n50373;
  assign n51699 = ~n51768;
  assign n51756 = n47836 & n50460;
  assign n51758 = n47836 & n49137;
  assign n47884 = ~n47836;
  assign n51776 = ~n51789;
  assign n47588 = n51681 ^ n48749;
  assign n51586 = n51681 & n48751;
  assign n51682 = n51681 & n48749;
  assign n51661 = n51719 ^ n51720;
  assign n51706 = n51726 & n51727;
  assign n51730 = n51739 & n51740;
  assign n51672 = ~n51754;
  assign n51741 = ~n51755;
  assign n50462 = ~n51756;
  assign n51744 = n47884 & n51757;
  assign n50404 = ~n51758;
  assign n51759 = n51776 & n51777;
  assign n47590 = ~n47588;
  assign n50663 = ~n51682;
  assign n51692 = n51661 & n9053;
  assign n51683 = n51706 ^ n51707;
  assign n51693 = ~n51661;
  assign n51708 = ~n51706;
  assign n51721 = ~n51730;
  assign n51628 = n51741 & n51742;
  assign n50498 = ~n51744;
  assign n51731 = n51759 ^ n49076;
  assign n51760 = ~n51759;
  assign n51654 = n47590 & n50636;
  assign n51659 = n500 ^ n51683;
  assign n51663 = ~n51692;
  assign n51684 = n51693 & n499;
  assign n51701 = n51708 & n51709;
  assign n51694 = n51721 & n51722;
  assign n51724 = n51628 & n51725;
  assign n51723 = ~n51628;
  assign n47792 = n51731 ^ n51732;
  assign n51745 = n51760 & n51761;
  assign n51636 = ~n51654;
  assign n51647 = n51658 ^ n51659;
  assign n51611 = n51659 & n51658;
  assign n51635 = ~n51684;
  assign n51670 = n51694 ^ n51695;
  assign n51679 = ~n51701;
  assign n51698 = ~n51694;
  assign n51713 = n47792 & n50390;
  assign n51714 = n47792 & n49076;
  assign n51710 = n51723 & n51651;
  assign n51712 = n47792 & n50292;
  assign n51653 = ~n51724;
  assign n47842 = ~n47792;
  assign n51733 = ~n51745;
  assign n51615 = n51636 & n51637;
  assign n51639 = n51647 & n48688;
  assign n51638 = ~n51647;
  assign n51619 = n51669 ^ n51670;
  assign n51660 = n51679 & n51680;
  assign n51685 = n51698 & n51699;
  assign n51631 = ~n51710;
  assign n51702 = n47842 & n51711;
  assign n51696 = ~n51712;
  assign n50392 = ~n51713;
  assign n50326 = ~n51714;
  assign n51716 = n51733 & n51734;
  assign n51584 = n51615 ^ n51616;
  assign n51613 = ~n51615;
  assign n51633 = n51638 & n48695;
  assign n51588 = ~n51639;
  assign n51648 = n51619 & n9015;
  assign n51640 = n51660 ^ n51661;
  assign n51649 = ~n51619;
  assign n51662 = ~n51660;
  assign n51671 = ~n51685;
  assign n51575 = n51696 & n51697;
  assign n50431 = ~n51702;
  assign n47736 = n51715 ^ n51716;
  assign n51717 = ~n51716;
  assign n49269 = n135 ^ n51584;
  assign n51329 = n51584 & n135;
  assign n51452 = n51613 & n51614;
  assign n51617 = ~n51633;
  assign n51612 = n499 ^ n51640;
  assign n51621 = ~n51648;
  assign n51641 = n51649 & n498;
  assign n51655 = n51662 & n51663;
  assign n51650 = n51671 & n51672;
  assign n51675 = n51575 & n51602;
  assign n51673 = ~n51575;
  assign n51686 = n47736 & n50126;
  assign n51688 = n47736 & n51700;
  assign n51689 = n47736 & n49027;
  assign n47796 = ~n47736;
  assign n51703 = n51717 & n51718;
  assign n50572 = ~n49269;
  assign n51525 = n51611 ^ n51612;
  assign n51607 = n51617 & n51586;
  assign n51585 = n51617 & n51588;
  assign n51560 = n51612 & n51611;
  assign n51592 = ~n51641;
  assign n51629 = n51650 ^ n51651;
  assign n51634 = ~n51655;
  assign n51652 = ~n51650;
  assign n51664 = n51673 & n51674;
  assign n51606 = ~n51675;
  assign n51676 = ~n51686;
  assign n51678 = n47796 & n51687;
  assign n50356 = ~n51688;
  assign n50269 = ~n51689;
  assign n51690 = ~n51703;
  assign n47494 = n51585 ^ n51586;
  assign n51589 = n51525 & n48676;
  assign n51587 = ~n51607;
  assign n51583 = ~n51525;
  assign n51563 = ~n51560;
  assign n51565 = n51628 ^ n51629;
  assign n51618 = n51634 & n51635;
  assign n51642 = n51652 & n51653;
  assign n51578 = ~n51664;
  assign n51485 = n51676 & n51677;
  assign n50312 = ~n51678;
  assign n51665 = n51690 & n51691;
  assign n51555 = n47494 & n50516;
  assign n51556 = n47494 & n48695;
  assign n47509 = ~n47494;
  assign n51581 = n51583 & n48654;
  assign n51557 = n51587 & n51588;
  assign n51528 = ~n51589;
  assign n51600 = n51565 & n497;
  assign n51590 = n51618 ^ n51619;
  assign n51599 = ~n51565;
  assign n51620 = ~n51618;
  assign n51630 = ~n51642;
  assign n51656 = n50356 & n50312;
  assign n51643 = n51665 ^ n51666;
  assign n51667 = ~n51665;
  assign n51540 = ~n51555;
  assign n50540 = ~n51556;
  assign n51526 = n51557 ^ n48654;
  assign n51559 = ~n51557;
  assign n51558 = ~n51581;
  assign n51561 = n498 ^ n51590;
  assign n51593 = n51599 & n8981;
  assign n51533 = ~n51600;
  assign n51608 = n51620 & n51621;
  assign n51601 = n51630 & n51631;
  assign n47689 = n49004 ^ n51643;
  assign n51644 = n51643 & n48949;
  assign n50354 = ~n51656;
  assign n51657 = n51667 & n51668;
  assign n47435 = n51525 ^ n51526;
  assign n51522 = n51540 & n51541;
  assign n51549 = n51558 & n51559;
  assign n51465 = n51560 ^ n51561;
  assign n51562 = ~n51561;
  assign n51567 = ~n51593;
  assign n51576 = n51601 ^ n51602;
  assign n51591 = ~n51608;
  assign n51605 = ~n51601;
  assign n51622 = n47689 & n49964;
  assign n51623 = n47689 & n51632;
  assign n47719 = ~n47689;
  assign n50167 = ~n51644;
  assign n51645 = ~n51657;
  assign n51497 = n47435 & n50419;
  assign n51498 = n47435 & n48654;
  assign n51515 = n51522 & n51523;
  assign n47465 = ~n47435;
  assign n51513 = ~n51522;
  assign n51529 = n51465 & n48624;
  assign n51527 = ~n51549;
  assign n51530 = ~n51465;
  assign n51500 = n51562 & n51563;
  assign n51505 = n51575 ^ n51576;
  assign n51564 = n51591 & n51592;
  assign n51594 = n51605 & n51606;
  assign n51609 = n47719 & n50271;
  assign n51603 = ~n51622;
  assign n50230 = ~n51623;
  assign n51624 = n51645 & n51646;
  assign n51480 = ~n51497;
  assign n50484 = ~n51498;
  assign n51496 = n51513 & n51514;
  assign n51483 = ~n51515;
  assign n51499 = n51527 & n51528;
  assign n51494 = ~n51529;
  assign n51524 = n51530 & n48644;
  assign n51503 = ~n51500;
  assign n51542 = n51505 & n8944;
  assign n51531 = n51564 ^ n51565;
  assign n51543 = ~n51505;
  assign n51566 = ~n51564;
  assign n51577 = ~n51594;
  assign n51462 = n51603 & n51604;
  assign n50273 = ~n51609;
  assign n51595 = n51624 ^ n51625;
  assign n51626 = ~n51624;
  assign n51371 = n51480 & n51481;
  assign n51482 = n51483 & n51452;
  assign n51459 = ~n51496;
  assign n51466 = n51499 ^ n48644;
  assign n51495 = ~n51499;
  assign n51468 = ~n51524;
  assign n51501 = n497 ^ n51531;
  assign n51507 = ~n51542;
  assign n51534 = n51543 & n496;
  assign n51550 = n51566 & n51567;
  assign n51551 = n51577 & n51578;
  assign n51580 = n51462 & n51582;
  assign n51579 = ~n51462;
  assign n47649 = n48910 ^ n51595;
  assign n51596 = n51595 & n48968;
  assign n51610 = n51626 & n51627;
  assign n51450 = n51371 & n51414;
  assign n51448 = ~n51371;
  assign n47383 = n51465 ^ n51466;
  assign n51458 = ~n51482;
  assign n51451 = n51459 & n51483;
  assign n51486 = n51494 & n51495;
  assign n51393 = n51500 ^ n51501;
  assign n51502 = ~n51501;
  assign n51473 = ~n51534;
  assign n51532 = ~n51550;
  assign n51548 = n51551 & n51552;
  assign n51546 = ~n51551;
  assign n51568 = n51579 & n51418;
  assign n51569 = n47649 & n49917;
  assign n51464 = ~n51580;
  assign n51570 = n47649 & n50191;
  assign n47716 = ~n47649;
  assign n50061 = ~n51596;
  assign n51597 = ~n51610;
  assign n51429 = n51448 & n51449;
  assign n51430 = n47383 & n50382;
  assign n51419 = ~n51450;
  assign n51431 = n47383 & n48624;
  assign n51420 = n51451 ^ n51452;
  assign n51453 = n51458 & n51459;
  assign n47411 = ~n47383;
  assign n51469 = n51393 & n48609;
  assign n51467 = ~n51486;
  assign n51470 = ~n51393;
  assign n51435 = n51502 & n51503;
  assign n51504 = n51532 & n51533;
  assign n51535 = n51546 & n51547;
  assign n51519 = ~n51548;
  assign n51423 = ~n51568;
  assign n51544 = ~n51569;
  assign n50151 = ~n51570;
  assign n51553 = n47716 & n51571;
  assign n51572 = n51597 & n51598;
  assign n51412 = n51420 & n134;
  assign n51383 = ~n51429;
  assign n51408 = ~n51430;
  assign n50414 = ~n51431;
  assign n51411 = ~n51420;
  assign n51413 = ~n51453;
  assign n51432 = n51467 & n51468;
  assign n51396 = ~n51469;
  assign n51460 = n51470 & n48588;
  assign n51438 = ~n51435;
  assign n51471 = n51504 ^ n51505;
  assign n51506 = ~n51504;
  assign n51516 = n51519 & n51485;
  assign n51489 = ~n51535;
  assign n51346 = n51544 & n51545;
  assign n50193 = ~n51553;
  assign n51537 = n51572 ^ n48895;
  assign n51573 = ~n51572;
  assign n51302 = n51408 & n51409;
  assign n51392 = n51411 & n6633;
  assign n51334 = ~n51412;
  assign n51372 = n51413 ^ n51414;
  assign n51410 = n51419 & n51413;
  assign n51394 = n51432 ^ n48588;
  assign n51433 = ~n51432;
  assign n51434 = ~n51460;
  assign n51436 = n496 ^ n51471;
  assign n51487 = n51506 & n51507;
  assign n51488 = ~n51516;
  assign n51484 = n51489 & n51519;
  assign n51520 = n51346 & n51389;
  assign n51517 = ~n51346;
  assign n47602 = n51536 ^ n51537;
  assign n51554 = n51573 & n51574;
  assign n51277 = n51371 ^ n51372;
  assign n51374 = n51302 & n51384;
  assign n51373 = ~n51302;
  assign n51370 = ~n51392;
  assign n47306 = n51393 ^ n51394;
  assign n51382 = ~n51410;
  assign n51421 = n51433 & n51434;
  assign n51313 = n51435 ^ n51436;
  assign n51437 = ~n51436;
  assign n51400 = n51484 ^ n51485;
  assign n51472 = ~n51487;
  assign n51461 = n51488 & n51489;
  assign n51508 = n51517 & n51518;
  assign n51391 = ~n51520;
  assign n51509 = n47602 & n51521;
  assign n47673 = ~n47602;
  assign n51538 = ~n51554;
  assign n51327 = n51277 & n133;
  assign n51326 = ~n51277;
  assign n51356 = n51370 & n51329;
  assign n51357 = n51373 & n51342;
  assign n51328 = n51370 & n51334;
  assign n51358 = n47306 & n50251;
  assign n51343 = ~n51374;
  assign n51359 = n47306 & n48588;
  assign n51341 = n51382 & n51383;
  assign n47336 = ~n47306;
  assign n51398 = n51313 & n48577;
  assign n51395 = ~n51421;
  assign n51397 = ~n51313;
  assign n51354 = n51437 & n51438;
  assign n51455 = n51400 & n511;
  assign n51417 = n51461 ^ n51462;
  assign n51439 = n51472 & n51473;
  assign n51454 = ~n51400;
  assign n51463 = ~n51461;
  assign n51349 = ~n51508;
  assign n51490 = n47673 & n49836;
  assign n50106 = ~n51509;
  assign n51491 = n47673 & n50062;
  assign n51492 = n47673 & n48895;
  assign n51510 = n51538 & n51539;
  assign n51315 = n51326 & n6535;
  assign n51244 = ~n51327;
  assign n49227 = n51328 ^ n51329;
  assign n51303 = n51341 ^ n51342;
  assign n51333 = ~n51356;
  assign n51305 = ~n51357;
  assign n51331 = ~n51358;
  assign n50314 = ~n51359;
  assign n51344 = ~n51341;
  assign n51360 = n51395 & n51396;
  assign n51385 = n51397 & n48553;
  assign n51361 = ~n51398;
  assign n51336 = n51417 ^ n51418;
  assign n51364 = ~n51354;
  assign n51399 = n511 ^ n51439;
  assign n51440 = n51454 & n8895;
  assign n51376 = ~n51455;
  assign n51416 = ~n51439;
  assign n51456 = n51463 & n51464;
  assign n51474 = ~n51490;
  assign n50065 = ~n51491;
  assign n49991 = ~n51492;
  assign n51477 = n51510 ^ n48882;
  assign n51511 = ~n51510;
  assign n51204 = n51302 ^ n51303;
  assign n51290 = ~n51315;
  assign n50491 = ~n49227;
  assign n51224 = n51331 & n51332;
  assign n51316 = n51333 & n51334;
  assign n51330 = n51343 & n51344;
  assign n51314 = n51360 ^ n48553;
  assign n51362 = ~n51360;
  assign n51318 = ~n51385;
  assign n51355 = n51399 ^ n51400;
  assign n51387 = n51336 & n510;
  assign n51386 = ~n51336;
  assign n51415 = ~n51440;
  assign n51422 = ~n51456;
  assign n51268 = n51474 & n51475;
  assign n47552 = n51476 ^ n51477;
  assign n51493 = n51511 & n51512;
  assign n51262 = n51204 & n132;
  assign n51261 = ~n51204;
  assign n51293 = n51224 & n51264;
  assign n47248 = n51313 ^ n51314;
  assign n51291 = ~n51224;
  assign n51276 = ~n51316;
  assign n51304 = ~n51330;
  assign n51238 = n51354 ^ n51355;
  assign n51345 = n51361 & n51362;
  assign n51363 = ~n51355;
  assign n51377 = n51386 & n8851;
  assign n51296 = ~n51387;
  assign n51401 = n51415 & n51416;
  assign n51388 = n51422 & n51423;
  assign n51443 = n51268 & n51310;
  assign n51444 = n47552 & n51457;
  assign n51441 = ~n51268;
  assign n47623 = ~n47552;
  assign n51478 = ~n51493;
  assign n51245 = n51261 & n6467;
  assign n51176 = ~n51262;
  assign n51236 = n51276 ^ n51277;
  assign n51275 = n51290 & n51276;
  assign n51278 = n51291 & n51292;
  assign n51265 = ~n51293;
  assign n51279 = n47248 & n50195;
  assign n51280 = n47248 & n48577;
  assign n51263 = n51304 & n51305;
  assign n47292 = ~n47248;
  assign n51319 = n51238 & n48516;
  assign n51317 = ~n51345;
  assign n51320 = ~n51238;
  assign n51249 = n51363 & n51364;
  assign n51337 = ~n51377;
  assign n51347 = n51388 ^ n51389;
  assign n51375 = ~n51401;
  assign n51390 = ~n51388;
  assign n51424 = n51441 & n51442;
  assign n51312 = ~n51443;
  assign n51425 = n47623 & n49865;
  assign n51426 = n47623 & n49974;
  assign n51427 = n47623 & n48855;
  assign n50027 = ~n51444;
  assign n51445 = n51478 & n51479;
  assign n49183 = n133 ^ n51236;
  assign n51212 = ~n51245;
  assign n51225 = n51263 ^ n51264;
  assign n51243 = ~n51275;
  assign n51223 = ~n51278;
  assign n51247 = ~n51279;
  assign n50238 = ~n51280;
  assign n51266 = ~n51263;
  assign n51281 = n51317 & n51318;
  assign n51241 = ~n51319;
  assign n51306 = n51320 & n48514;
  assign n51253 = n51346 ^ n51347;
  assign n51335 = n51375 & n51376;
  assign n51378 = n51390 & n51391;
  assign n51271 = ~n51424;
  assign n51402 = ~n51425;
  assign n49977 = ~n51426;
  assign n49902 = ~n51427;
  assign n51405 = n51445 ^ n48815;
  assign n51446 = ~n51445;
  assign n51147 = n51224 ^ n51225;
  assign n50428 = ~n49183;
  assign n51237 = n51243 & n51244;
  assign n51160 = n51247 & n51248;
  assign n51246 = n51265 & n51266;
  assign n51239 = n51281 ^ n48514;
  assign n51282 = ~n51281;
  assign n51283 = ~n51306;
  assign n51307 = n51253 & n8797;
  assign n51294 = n51335 ^ n51336;
  assign n51308 = ~n51253;
  assign n51338 = ~n51335;
  assign n51348 = ~n51378;
  assign n51196 = n51402 & n51403;
  assign n47505 = n51404 ^ n51405;
  assign n51428 = n51446 & n51447;
  assign n51189 = n51147 & n6372;
  assign n51190 = ~n51147;
  assign n51214 = n51160 & n51226;
  assign n51203 = ~n51237;
  assign n51213 = ~n51160;
  assign n47232 = n51238 ^ n51239;
  assign n51222 = ~n51246;
  assign n51267 = n51282 & n51283;
  assign n51250 = n510 ^ n51294;
  assign n51254 = ~n51307;
  assign n51297 = n51308 & n509;
  assign n51321 = n51337 & n51338;
  assign n51309 = n51348 & n51349;
  assign n51366 = n51196 & n51379;
  assign n51367 = n47505 & n51380;
  assign n51365 = ~n51196;
  assign n47559 = ~n47505;
  assign n51406 = ~n51428;
  assign n51148 = ~n51189;
  assign n51177 = n51190 & n131;
  assign n51170 = n51203 ^ n51204;
  assign n51202 = n51212 & n51203;
  assign n51205 = n51213 & n51192;
  assign n51206 = n47232 & n50084;
  assign n51194 = ~n51214;
  assign n51207 = n47232 & n48514;
  assign n51191 = n51222 & n51223;
  assign n47251 = ~n47232;
  assign n51172 = n51249 ^ n51250;
  assign n51240 = ~n51267;
  assign n51251 = ~n51250;
  assign n51217 = ~n51297;
  assign n51269 = n51309 ^ n51310;
  assign n51295 = ~n51321;
  assign n51311 = ~n51309;
  assign n51350 = n51365 & n51230;
  assign n51351 = n47559 & n49781;
  assign n51232 = ~n51366;
  assign n51352 = n47559 & n48815;
  assign n51353 = n47559 & n49887;
  assign n49938 = ~n51367;
  assign n51368 = n51406 & n51407;
  assign n49122 = n132 ^ n51170;
  assign n51115 = ~n51177;
  assign n51161 = n51191 ^ n51192;
  assign n51175 = ~n51202;
  assign n51163 = ~n51205;
  assign n51178 = ~n51206;
  assign n50155 = ~n51207;
  assign n51193 = ~n51191;
  assign n51208 = n51240 & n51241;
  assign n51182 = ~n51172;
  assign n51183 = n51251 & n51249;
  assign n51186 = n51268 ^ n51269;
  assign n51252 = n51295 & n51296;
  assign n51298 = n51311 & n51312;
  assign n51199 = ~n51350;
  assign n51322 = ~n51351;
  assign n49818 = ~n51352;
  assign n49890 = ~n51353;
  assign n51325 = n51368 ^ n48787;
  assign n51369 = n51368 & n51381;
  assign n49156 = ~n49122;
  assign n51085 = n51160 ^ n51161;
  assign n51146 = n51175 & n51176;
  assign n51098 = n51178 & n51179;
  assign n51180 = n51193 & n51194;
  assign n51171 = n51208 ^ n48496;
  assign n51210 = n51208 & n48496;
  assign n51209 = ~n51208;
  assign n51227 = n51186 & n8745;
  assign n51215 = n51252 ^ n51253;
  assign n51228 = ~n51186;
  assign n51255 = ~n51252;
  assign n51270 = ~n51298;
  assign n51137 = n51322 & n51323;
  assign n47454 = n51324 ^ n51325;
  assign n51339 = ~n51369;
  assign n51130 = n51085 & n130;
  assign n51113 = n51146 ^ n51147;
  assign n51129 = ~n51085;
  assign n51152 = n51098 & n51132;
  assign n51149 = ~n51146;
  assign n51150 = ~n51098;
  assign n47195 = n51171 ^ n51172;
  assign n51162 = ~n51180;
  assign n51195 = n51209 & n48463;
  assign n51181 = ~n51210;
  assign n51184 = n509 ^ n51215;
  assign n51188 = ~n51227;
  assign n51218 = n51228 & n508;
  assign n51242 = n51254 & n51255;
  assign n51229 = n51270 & n51271;
  assign n51288 = n47454 & n51289;
  assign n51285 = n47454 & n49605;
  assign n51286 = n51137 & n51299;
  assign n51287 = n47454 & n48787;
  assign n51284 = ~n51137;
  assign n47462 = ~n47454;
  assign n51300 = n51339 & n51340;
  assign n51083 = n131 ^ n51113;
  assign n51116 = n51129 & n6286;
  assign n51055 = ~n51130;
  assign n51141 = n51148 & n51149;
  assign n51142 = n51150 & n51151;
  assign n51134 = ~n51152;
  assign n51131 = n51162 & n51163;
  assign n47202 = ~n47195;
  assign n51173 = n51181 & n51182;
  assign n51088 = n51183 ^ n51184;
  assign n51145 = ~n51195;
  assign n51121 = n51184 & n51183;
  assign n51157 = ~n51218;
  assign n51197 = n51229 ^ n51230;
  assign n51216 = ~n51242;
  assign n51231 = ~n51229;
  assign n51272 = n51284 & n51167;
  assign n51256 = ~n51285;
  assign n51169 = ~n51286;
  assign n49722 = ~n51287;
  assign n49807 = ~n51288;
  assign n51274 = n47462 & n49805;
  assign n49725 = n51300 ^ n51301;
  assign n50327 = n51083 ^ n49122;
  assign n51027 = n51083 & n49122;
  assign n51086 = ~n51116;
  assign n51099 = n51131 ^ n51132;
  assign n51114 = ~n51141;
  assign n51101 = ~n51142;
  assign n51135 = n47202 & n49999;
  assign n51136 = n47202 & n48496;
  assign n51133 = ~n51131;
  assign n51154 = n51088 & n48455;
  assign n51144 = ~n51173;
  assign n51153 = ~n51088;
  assign n51124 = ~n51121;
  assign n51126 = n51196 ^ n51197;
  assign n51185 = n51216 & n51217;
  assign n51219 = n51231 & n51232;
  assign n51076 = n51256 & n51257;
  assign n49769 = n51258 ^ n49725;
  assign n51140 = ~n51272;
  assign n51259 = n49725 & n51273;
  assign n51260 = n49725 & n48802;
  assign n49854 = ~n51274;
  assign n47468 = ~n49725;
  assign n50310 = ~n50327;
  assign n51031 = n51098 ^ n51099;
  assign n51084 = n51114 & n51115;
  assign n51117 = n51133 & n51134;
  assign n51109 = ~n51135;
  assign n50069 = ~n51136;
  assign n51118 = n51144 & n51145;
  assign n51143 = n51153 & n48419;
  assign n51091 = ~n51154;
  assign n51165 = n51126 & n507;
  assign n51155 = n51185 ^ n51186;
  assign n51164 = ~n51126;
  assign n51187 = ~n51185;
  assign n51198 = ~n51219;
  assign n51221 = n51076 & n51233;
  assign n51220 = ~n51076;
  assign n51234 = ~n51259;
  assign n49686 = ~n51260;
  assign n51071 = n51031 & n6214;
  assign n51056 = n51084 ^ n51085;
  assign n51070 = ~n51031;
  assign n51087 = ~n51084;
  assign n51042 = n51109 & n51110;
  assign n51100 = ~n51117;
  assign n51089 = n51118 ^ n48419;
  assign n51119 = ~n51118;
  assign n51120 = ~n51143;
  assign n51122 = n508 ^ n51155;
  assign n51158 = n51164 & n8665;
  assign n51095 = ~n51165;
  assign n51174 = n51187 & n51188;
  assign n51166 = n51198 & n51199;
  assign n51211 = n51220 & n51106;
  assign n51108 = ~n51221;
  assign n51200 = n51234 & n51235;
  assign n51028 = n130 ^ n51056;
  assign n51057 = n51070 & n129;
  assign n51032 = ~n51071;
  assign n51080 = n51086 & n51087;
  assign n47150 = n51088 ^ n51089;
  assign n51072 = n51100 & n51101;
  assign n51051 = ~n51042;
  assign n51111 = n51119 & n51120;
  assign n51102 = n51121 ^ n51122;
  assign n51123 = ~n51122;
  assign n51128 = ~n51158;
  assign n51138 = n51166 ^ n51167;
  assign n51156 = ~n51174;
  assign n51168 = ~n51166;
  assign n51023 = n51200 ^ n51201;
  assign n51079 = ~n51211;
  assign n49073 = n51027 ^ n51028;
  assign n51029 = ~n51028;
  assign n51007 = ~n51057;
  assign n51043 = n51072 ^ n51073;
  assign n51059 = n47150 & n49910;
  assign n51060 = n47150 & n48419;
  assign n51054 = ~n51080;
  assign n51075 = n51072 & n51081;
  assign n47166 = ~n47150;
  assign n51074 = ~n51072;
  assign n51092 = n51102 & n48413;
  assign n51090 = ~n51111;
  assign n51035 = ~n51102;
  assign n51064 = n51123 & n51124;
  assign n51067 = n51137 ^ n51138;
  assign n51125 = n51156 & n51157;
  assign n51159 = n51168 & n51169;
  assign n50216 = ~n49073;
  assign n50977 = n51029 & n51027;
  assign n50965 = n51042 ^ n51043;
  assign n51030 = n51054 & n51055;
  assign n51045 = ~n51059;
  assign n49980 = ~n51060;
  assign n51058 = n51074 & n51073;
  assign n51050 = ~n51075;
  assign n51061 = n51090 & n51091;
  assign n51082 = n51035 & n48381;
  assign n51063 = ~n51092;
  assign n51104 = n51067 & n506;
  assign n51093 = n51125 ^ n51126;
  assign n51103 = ~n51067;
  assign n51127 = ~n51125;
  assign n51139 = ~n51159;
  assign n50980 = ~n50977;
  assign n51005 = n51030 ^ n51031;
  assign n50972 = n51045 & n51046;
  assign n51033 = ~n51030;
  assign n51044 = n51050 & n51051;
  assign n51026 = ~n51058;
  assign n51034 = n51061 ^ n48413;
  assign n51062 = ~n51061;
  assign n51037 = ~n51082;
  assign n51065 = n507 ^ n51093;
  assign n51096 = n51103 & n8632;
  assign n51040 = ~n51104;
  assign n51112 = n51127 & n51128;
  assign n51105 = n51139 & n51140;
  assign n50978 = n129 ^ n51005;
  assign n51024 = n51032 & n51033;
  assign n50985 = ~n50972;
  assign n47110 = n51034 ^ n51035;
  assign n51025 = ~n51044;
  assign n51052 = n51062 & n51063;
  assign n50986 = n51064 ^ n51065;
  assign n51014 = n51065 & n51064;
  assign n51069 = ~n51096;
  assign n51077 = n51105 ^ n51106;
  assign n51094 = ~n51112;
  assign n51107 = ~n51105;
  assign n49015 = n50977 ^ n50978;
  assign n50979 = ~n50978;
  assign n51009 = n47110 & n49826;
  assign n51010 = n47110 & n48413;
  assign n51006 = ~n51024;
  assign n50999 = n51025 & n51026;
  assign n47140 = ~n47110;
  assign n51036 = ~n51052;
  assign n50998 = ~n50986;
  assign n51017 = ~n51014;
  assign n51019 = n51076 ^ n51077;
  assign n51066 = n51094 & n51095;
  assign n51097 = n51107 & n51108;
  assign n50102 = ~n49015;
  assign n50937 = n50979 & n50980;
  assign n50973 = n50999 ^ n51000;
  assign n50981 = n51006 & n51007;
  assign n51002 = n50999 & n51008;
  assign n50994 = ~n51009;
  assign n49893 = ~n51010;
  assign n51001 = ~n50999;
  assign n51011 = n51036 & n51037;
  assign n51048 = n51019 & n505;
  assign n51038 = n51066 ^ n51067;
  assign n51047 = ~n51019;
  assign n51068 = ~n51066;
  assign n51078 = ~n51097;
  assign n50920 = n50972 ^ n50973;
  assign n50955 = n50981 ^ n50965;
  assign n50983 = n50981 & n6136;
  assign n50923 = n50994 & n50995;
  assign n50982 = ~n50981;
  assign n50996 = n51001 & n51000;
  assign n50984 = ~n51002;
  assign n50987 = n51011 ^ n48341;
  assign n51013 = n51011 & n48372;
  assign n51012 = ~n51011;
  assign n51015 = n506 ^ n51038;
  assign n51041 = n51047 & n8583;
  assign n50993 = ~n51048;
  assign n51053 = n51068 & n51069;
  assign n51049 = n51078 & n51079;
  assign n50938 = n128 ^ n50955;
  assign n50967 = n50923 & n50975;
  assign n50974 = n50982 & n128;
  assign n50964 = ~n50983;
  assign n50971 = n50984 & n50985;
  assign n50966 = ~n50923;
  assign n47075 = n50986 ^ n50987;
  assign n50958 = ~n50996;
  assign n51003 = n51012 & n48341;
  assign n50997 = ~n51013;
  assign n50930 = n51014 ^ n51015;
  assign n51016 = ~n51015;
  assign n51021 = ~n51041;
  assign n51022 = n504 ^ n51049;
  assign n51039 = ~n51053;
  assign n50024 = n50937 ^ n50938;
  assign n50890 = n50938 & n50937;
  assign n50956 = n50964 & n50965;
  assign n50959 = n50966 & n50940;
  assign n50942 = ~n50967;
  assign n50960 = n47075 & n49761;
  assign n50961 = n47075 & n48372;
  assign n50957 = ~n50971;
  assign n50947 = ~n50974;
  assign n47081 = ~n47075;
  assign n50988 = n50997 & n50998;
  assign n50989 = n50930 & n48300;
  assign n50969 = ~n51003;
  assign n50990 = ~n50930;
  assign n50962 = n51016 & n51017;
  assign n50934 = n51022 ^ n51023;
  assign n51018 = n51039 & n51040;
  assign n48982 = ~n50024;
  assign n50946 = ~n50956;
  assign n50939 = n50957 & n50958;
  assign n50922 = ~n50959;
  assign n50948 = ~n50960;
  assign n49801 = ~n50961;
  assign n50968 = ~n50988;
  assign n50932 = ~n50989;
  assign n50976 = n50990 & n48331;
  assign n50970 = ~n50962;
  assign n50991 = n51018 ^ n51019;
  assign n51020 = ~n51018;
  assign n50924 = n50939 ^ n50940;
  assign n50926 = n50946 & n50947;
  assign n50887 = n50948 & n50949;
  assign n50941 = ~n50939;
  assign n50950 = n50968 & n50969;
  assign n50952 = ~n50976;
  assign n50963 = n505 ^ n50991;
  assign n51004 = n51020 & n51021;
  assign n50875 = n50923 ^ n50924;
  assign n50909 = n50926 ^ n50920;
  assign n50928 = n50926 & n6045;
  assign n50927 = ~n50926;
  assign n50935 = n50941 & n50942;
  assign n50893 = ~n50887;
  assign n50929 = n50950 ^ n48331;
  assign n50951 = ~n50950;
  assign n50895 = n50962 ^ n50963;
  assign n50954 = n50963 & n50970;
  assign n50992 = ~n51004;
  assign n50891 = n143 ^ n50909;
  assign n50925 = n50927 & n143;
  assign n50919 = ~n50928;
  assign n47025 = n50929 ^ n50930;
  assign n50921 = ~n50935;
  assign n50943 = n50951 & n50952;
  assign n50945 = n50895 & n48259;
  assign n50944 = ~n50895;
  assign n50953 = n50992 & n50993;
  assign n49935 = n50890 ^ n50891;
  assign n50849 = n50891 & n50890;
  assign n50910 = n50919 & n50920;
  assign n50912 = n47025 & n49652;
  assign n50913 = n47025 & n48331;
  assign n50903 = n50921 & n50922;
  assign n50899 = ~n50925;
  assign n47049 = ~n47025;
  assign n50931 = ~n50943;
  assign n50936 = n50944 & n48291;
  assign n50897 = ~n50945;
  assign n50933 = n50953 ^ n50954;
  assign n48939 = ~n49935;
  assign n50888 = n50903 ^ n50904;
  assign n50898 = ~n50910;
  assign n50906 = n50903 & n50911;
  assign n50900 = ~n50912;
  assign n49728 = ~n50913;
  assign n50905 = ~n50903;
  assign n50914 = n50931 & n50932;
  assign n50864 = n50933 ^ n50934;
  assign n50916 = ~n50936;
  assign n50830 = n50887 ^ n50888;
  assign n50884 = n50898 & n50899;
  assign n50843 = n50900 & n50901;
  assign n50902 = n50905 & n50904;
  assign n50892 = ~n50906;
  assign n50894 = n50914 ^ n48291;
  assign n50917 = n50864 & n48218;
  assign n50915 = ~n50914;
  assign n50918 = ~n50864;
  assign n50868 = n50884 ^ n50875;
  assign n50886 = n50884 & n5959;
  assign n50885 = ~n50884;
  assign n50889 = n50892 & n50893;
  assign n50852 = ~n50843;
  assign n46987 = n50894 ^ n50895;
  assign n50878 = ~n50902;
  assign n50907 = n50915 & n50916;
  assign n50883 = ~n50917;
  assign n50908 = n50918 & n48242;
  assign n50850 = n142 ^ n50868;
  assign n50876 = n50885 & n142;
  assign n50874 = ~n50886;
  assign n50879 = n46987 & n49577;
  assign n50880 = n46987 & n48291;
  assign n50877 = ~n50889;
  assign n47015 = ~n46987;
  assign n50896 = ~n50907;
  assign n50867 = ~n50908;
  assign n48903 = n50849 ^ n50850;
  assign n50808 = n50850 & n50849;
  assign n50869 = n50874 & n50875;
  assign n50857 = ~n50876;
  assign n50860 = n50877 & n50878;
  assign n50871 = ~n50879;
  assign n49637 = ~n50880;
  assign n50881 = n50896 & n50897;
  assign n49867 = ~n48903;
  assign n50807 = ~n50808;
  assign n50844 = n50860 ^ n50861;
  assign n50856 = ~n50869;
  assign n50863 = n50860 & n50870;
  assign n50799 = n50871 & n50872;
  assign n50862 = ~n50860;
  assign n50865 = n50881 ^ n48218;
  assign n50882 = ~n50881;
  assign n50783 = n50843 ^ n50844;
  assign n50837 = n50856 & n50857;
  assign n50854 = n50799 & n50859;
  assign n50858 = n50862 & n50861;
  assign n50851 = ~n50863;
  assign n50853 = ~n50799;
  assign n46949 = n50864 ^ n50865;
  assign n50873 = n50882 & n50883;
  assign n50825 = n50837 ^ n50830;
  assign n50839 = n50837 & n5852;
  assign n50838 = ~n50837;
  assign n50845 = n50851 & n50852;
  assign n50846 = n50853 & n50819;
  assign n50821 = ~n50854;
  assign n50835 = ~n50858;
  assign n46969 = ~n46949;
  assign n50866 = ~n50873;
  assign n50809 = n141 ^ n50825;
  assign n50833 = n50838 & n141;
  assign n50829 = ~n50839;
  assign n50834 = ~n50845;
  assign n50802 = ~n50846;
  assign n50840 = n46969 & n49514;
  assign n50841 = n46969 & n48218;
  assign n50855 = n50866 & n50867;
  assign n48859 = n50808 ^ n50809;
  assign n50806 = ~n50809;
  assign n50826 = n50829 & n50830;
  assign n50812 = ~n50833;
  assign n50818 = n50834 & n50835;
  assign n50827 = ~n50840;
  assign n49568 = ~n50841;
  assign n50848 = n50855 & n48210;
  assign n50847 = ~n50855;
  assign n49783 = ~n48859;
  assign n49723 = n50806 & n50807;
  assign n50800 = n50818 ^ n50819;
  assign n50811 = ~n50826;
  assign n50767 = n50827 & n50828;
  assign n50820 = ~n50818;
  assign n50842 = n50847 & n48174;
  assign n50832 = ~n50848;
  assign n50760 = ~n49723;
  assign n50737 = n50799 ^ n50800;
  assign n50798 = n50811 & n50812;
  assign n50813 = n50820 & n50821;
  assign n50815 = n50767 & n50822;
  assign n50814 = ~n50767;
  assign n50831 = n50832 & n50836;
  assign n50824 = ~n50842;
  assign n50796 = n50798 & n5747;
  assign n50792 = ~n50798;
  assign n50801 = ~n50813;
  assign n50810 = n50814 & n50785;
  assign n50787 = ~n50815;
  assign n50823 = ~n50831;
  assign n50817 = n50824 & n50832;
  assign n50777 = n50792 ^ n50783;
  assign n50793 = n50792 & n140;
  assign n50782 = ~n50796;
  assign n50784 = n50801 & n50802;
  assign n50770 = ~n50810;
  assign n46909 = n50816 ^ n50817;
  assign n50803 = n50823 & n50824;
  assign n49682 = n140 ^ n50777;
  assign n50778 = n50782 & n50783;
  assign n50768 = n50784 ^ n50785;
  assign n50766 = ~n50793;
  assign n50786 = ~n50784;
  assign n50788 = n50803 ^ n48166;
  assign n46938 = ~n46909;
  assign n50804 = ~n50803;
  assign n50759 = ~n49682;
  assign n50703 = n50767 ^ n50768;
  assign n50765 = ~n50778;
  assign n50779 = n50786 & n50787;
  assign n46866 = n50788 ^ n50789;
  assign n50794 = n46938 & n49468;
  assign n50795 = n46938 & n48210;
  assign n50797 = n50804 & n50805;
  assign n50711 = n50759 & n50760;
  assign n50750 = n50703 & n138;
  assign n50748 = ~n50703;
  assign n50746 = n50765 & n50766;
  assign n50771 = n46866 & n49400;
  assign n50772 = n46866 & n48166;
  assign n50769 = ~n50779;
  assign n46901 = ~n46866;
  assign n50780 = ~n50794;
  assign n49491 = ~n50795;
  assign n50790 = ~n50797;
  assign n50726 = n50746 ^ n50737;
  assign n50744 = n50748 & n5626;
  assign n50682 = ~n50750;
  assign n50749 = n50746 & n5694;
  assign n50747 = ~n50746;
  assign n50751 = n50769 & n50770;
  assign n50762 = ~n50771;
  assign n49450 = ~n50772;
  assign n50728 = n50780 & n50781;
  assign n50773 = n50790 & n50791;
  assign n50712 = n139 ^ n50726;
  assign n50701 = ~n50744;
  assign n50743 = n50747 & n139;
  assign n50736 = ~n50749;
  assign n50729 = n50751 ^ n50752;
  assign n50754 = n50751 & n50761;
  assign n50683 = n50762 & n50763;
  assign n50753 = ~n50751;
  assign n50755 = n50773 ^ n50774;
  assign n50739 = ~n50728;
  assign n50775 = ~n50773;
  assign n50691 = n50711 ^ n50712;
  assign n50664 = n50712 & n50711;
  assign n50667 = n50728 ^ n50729;
  assign n50727 = n50736 & n50737;
  assign n50721 = ~n50743;
  assign n50742 = n50683 & n50705;
  assign n50745 = n50753 & n50752;
  assign n50738 = ~n50754;
  assign n50740 = ~n50683;
  assign n46802 = n48070 ^ n50755;
  assign n50756 = n50755 & n48070;
  assign n50764 = n50775 & n50776;
  assign n46551 = n50691 ^ n47588;
  assign n50692 = ~n50691;
  assign n50713 = n50667 & n137;
  assign n50710 = ~n50667;
  assign n50720 = ~n50727;
  assign n50730 = n50738 & n50739;
  assign n50731 = n50740 & n50741;
  assign n50707 = ~n50742;
  assign n50723 = ~n50745;
  assign n46849 = ~n46802;
  assign n49402 = ~n50756;
  assign n50757 = ~n50764;
  assign n50673 = n46551 & n48751;
  assign n46549 = ~n46551;
  assign n50583 = n50692 & n47590;
  assign n50687 = n50692 & n47588;
  assign n50709 = n50710 & n5602;
  assign n50632 = ~n50713;
  assign n50702 = n50720 & n50721;
  assign n50722 = ~n50730;
  assign n50686 = ~n50731;
  assign n50724 = n46849 & n49337;
  assign n50732 = n50757 & n50758;
  assign n50662 = ~n50673;
  assign n48763 = ~n50687;
  assign n50680 = n50702 ^ n50703;
  assign n50661 = ~n50709;
  assign n50700 = ~n50702;
  assign n50704 = n50722 & n50723;
  assign n50714 = ~n50724;
  assign n50716 = n50732 ^ n50733;
  assign n50734 = ~n50732;
  assign n50633 = n50662 & n50663;
  assign n50665 = n138 ^ n50680;
  assign n50693 = n50700 & n50701;
  assign n50684 = n50704 ^ n50705;
  assign n50706 = ~n50704;
  assign n50671 = n50714 & n50715;
  assign n46784 = n50716 ^ n48084;
  assign n50717 = n50716 & n48084;
  assign n50725 = n50734 & n50735;
  assign n50610 = n50633 ^ n50634;
  assign n50635 = ~n50633;
  assign n50644 = n50664 ^ n50665;
  assign n50613 = n50665 & n50664;
  assign n50616 = n50683 ^ n50684;
  assign n50681 = ~n50693;
  assign n50694 = n50706 & n50707;
  assign n50696 = n50671 & n50708;
  assign n50695 = ~n50671;
  assign n46813 = ~n46784;
  assign n49360 = ~n50717;
  assign n50718 = ~n50725;
  assign n48629 = n295 ^ n50610;
  assign n50331 = n50610 & n295;
  assign n50450 = n50635 & n50636;
  assign n50637 = n50644 & n47509;
  assign n50638 = ~n50644;
  assign n50668 = n50616 & n5544;
  assign n50669 = ~n50616;
  assign n50666 = n50681 & n50682;
  assign n50685 = ~n50694;
  assign n50688 = n50695 & n50641;
  assign n50659 = ~n50696;
  assign n50689 = n46813 & n49319;
  assign n50697 = n50718 & n50719;
  assign n50259 = ~n48629;
  assign n50612 = ~n50637;
  assign n50624 = n50638 & n47494;
  assign n50639 = n50666 ^ n50667;
  assign n50609 = ~n50668;
  assign n50650 = n50669 & n136;
  assign n50660 = ~n50666;
  assign n50670 = n50685 & n50686;
  assign n50643 = ~n50688;
  assign n50674 = ~n50689;
  assign n50676 = n50697 ^ n48021;
  assign n50698 = ~n50697;
  assign n50611 = n50612 & n50583;
  assign n50596 = ~n50624;
  assign n50614 = n137 ^ n50639;
  assign n50587 = ~n50650;
  assign n50649 = n50660 & n50661;
  assign n50640 = n50670 ^ n50671;
  assign n50658 = ~n50670;
  assign n50588 = n50674 & n50675;
  assign n46720 = n50676 ^ n50677;
  assign n50690 = n50698 & n50699;
  assign n50595 = ~n50611;
  assign n50582 = n50612 & n50596;
  assign n50594 = n50613 ^ n50614;
  assign n50560 = n50614 & n50613;
  assign n50530 = n50640 ^ n50641;
  assign n50631 = ~n50649;
  assign n50651 = n50658 & n50659;
  assign n50653 = n50588 & n50672;
  assign n50652 = ~n50588;
  assign n46772 = ~n46720;
  assign n50678 = ~n50690;
  assign n46432 = n50582 ^ n50583;
  assign n50584 = n50594 & n47465;
  assign n50574 = n50595 & n50596;
  assign n50538 = ~n50594;
  assign n50618 = n50530 & n151;
  assign n50617 = ~n50530;
  assign n50615 = n50631 & n50632;
  assign n50646 = n46772 & n49291;
  assign n50642 = ~n50651;
  assign n50645 = n50652 & n50620;
  assign n50622 = ~n50653;
  assign n50647 = n46772 & n48021;
  assign n50654 = n50678 & n50679;
  assign n50557 = n46432 & n48688;
  assign n50558 = n46432 & n47509;
  assign n50537 = n50574 ^ n47465;
  assign n46439 = ~n46432;
  assign n50576 = ~n50574;
  assign n50575 = ~n50584;
  assign n50577 = n50538 & n47435;
  assign n50585 = n50615 ^ n50616;
  assign n50600 = n50617 & n5509;
  assign n50532 = ~n50618;
  assign n50608 = ~n50615;
  assign n50619 = n50642 & n50643;
  assign n50591 = ~n50645;
  assign n50625 = ~n50646;
  assign n49308 = ~n50647;
  assign n50627 = n50654 ^ n50655;
  assign n50656 = ~n50654;
  assign n46371 = n50537 ^ n50538;
  assign n50539 = ~n50557;
  assign n48702 = ~n50558;
  assign n50559 = n50575 & n50576;
  assign n50546 = ~n50577;
  assign n50561 = n136 ^ n50585;
  assign n50565 = ~n50600;
  assign n50599 = n50608 & n50609;
  assign n50589 = n50619 ^ n50620;
  assign n50621 = ~n50619;
  assign n50569 = n50625 & n50626;
  assign n46699 = n47958 ^ n50627;
  assign n50628 = n50627 & n48003;
  assign n50648 = n50656 & n50657;
  assign n50513 = n46371 & n48676;
  assign n50514 = n46371 & n47465;
  assign n46335 = ~n46371;
  assign n50521 = n50539 & n50540;
  assign n50545 = ~n50559;
  assign n50475 = n50560 ^ n50561;
  assign n50562 = ~n50561;
  assign n50504 = n50588 ^ n50589;
  assign n50586 = ~n50599;
  assign n50601 = n50621 & n50622;
  assign n50603 = n50569 & n50623;
  assign n50604 = n46699 & n49247;
  assign n50602 = ~n50569;
  assign n46734 = ~n46699;
  assign n49267 = ~n50628;
  assign n50629 = ~n50648;
  assign n50483 = ~n50513;
  assign n48685 = ~n50514;
  assign n50517 = n50521 & n50522;
  assign n50515 = ~n50521;
  assign n50518 = n50545 & n50546;
  assign n50501 = n50562 & n50560;
  assign n50567 = n50504 & n150;
  assign n50566 = ~n50504;
  assign n50563 = n50586 & n50587;
  assign n50590 = ~n50601;
  assign n50597 = n50602 & n50534;
  assign n50556 = ~n50603;
  assign n50592 = ~n50604;
  assign n50605 = n50629 & n50630;
  assign n50377 = n50483 & n50484;
  assign n50499 = n50515 & n50516;
  assign n50477 = ~n50517;
  assign n50474 = n50518 ^ n47411;
  assign n50520 = n50518 & n47411;
  assign n50519 = ~n50518;
  assign n50529 = n151 ^ n50563;
  assign n50548 = n50566 & n5464;
  assign n50467 = ~n50567;
  assign n50564 = ~n50563;
  assign n50568 = n50590 & n50591;
  assign n50468 = n50592 & n50593;
  assign n50536 = ~n50597;
  assign n50579 = n50605 ^ n47918;
  assign n50606 = ~n50605;
  assign n50455 = n50377 & n50463;
  assign n50454 = ~n50377;
  assign n46262 = n50474 ^ n50475;
  assign n50476 = n50477 & n50450;
  assign n50457 = ~n50499;
  assign n50500 = n50519 & n47383;
  assign n50485 = ~n50520;
  assign n50502 = n50529 ^ n50530;
  assign n50506 = ~n50548;
  assign n50547 = n50564 & n50565;
  assign n50533 = n50568 ^ n50569;
  assign n50573 = n50468 & n50510;
  assign n50555 = ~n50568;
  assign n50570 = ~n50468;
  assign n46660 = n50578 ^ n50579;
  assign n50598 = n50606 & n50607;
  assign n50446 = n50454 & n50419;
  assign n50415 = ~n50455;
  assign n50447 = n46262 & n48644;
  assign n50448 = n46262 & n47411;
  assign n46303 = ~n46262;
  assign n50456 = ~n50476;
  assign n50449 = n50457 & n50477;
  assign n50478 = n50485 & n50475;
  assign n50453 = ~n50500;
  assign n50479 = n50501 ^ n50502;
  assign n50432 = n50502 & n50501;
  assign n50435 = n50533 ^ n50534;
  assign n50531 = ~n50547;
  assign n50549 = n50555 & n50556;
  assign n50550 = n50570 & n50571;
  assign n50551 = n46660 & n50572;
  assign n50512 = ~n50573;
  assign n46688 = ~n46660;
  assign n50580 = ~n50598;
  assign n50380 = ~n50446;
  assign n50413 = ~n50447;
  assign n48656 = ~n50448;
  assign n50417 = n50449 ^ n50450;
  assign n50418 = n50456 & n50457;
  assign n50452 = ~n50478;
  assign n50464 = n50479 & n47336;
  assign n50385 = ~n50479;
  assign n50508 = n50435 & n149;
  assign n50507 = ~n50435;
  assign n50503 = n50531 & n50532;
  assign n50535 = ~n50549;
  assign n50471 = ~n50550;
  assign n49295 = ~n50551;
  assign n50541 = n46688 & n49193;
  assign n50542 = n46688 & n49269;
  assign n50543 = n46688 & n47918;
  assign n50552 = n50580 & n50581;
  assign n50302 = n50413 & n50414;
  assign n50407 = n50417 & n294;
  assign n50378 = n50418 ^ n50419;
  assign n50406 = ~n50417;
  assign n50416 = ~n50418;
  assign n50420 = n50452 & n50453;
  assign n50458 = n50385 & n47306;
  assign n50412 = ~n50464;
  assign n50465 = n50503 ^ n50504;
  assign n50487 = n50507 & n5423;
  assign n50398 = ~n50508;
  assign n50505 = ~n50503;
  assign n50509 = n50535 & n50536;
  assign n50523 = ~n50541;
  assign n49272 = ~n50542;
  assign n49240 = ~n50543;
  assign n50526 = n50552 ^ n47878;
  assign n50553 = ~n50552;
  assign n50280 = n50377 ^ n50378;
  assign n50383 = n50302 & n50339;
  assign n50381 = ~n50302;
  assign n50393 = n50406 & n2545;
  assign n50333 = ~n50407;
  assign n50405 = n50415 & n50416;
  assign n50384 = n50420 ^ n47336;
  assign n50411 = ~n50420;
  assign n50387 = ~n50458;
  assign n50433 = n150 ^ n50465;
  assign n50437 = ~n50487;
  assign n50486 = n50505 & n50506;
  assign n50469 = n50509 ^ n50510;
  assign n50511 = ~n50509;
  assign n50399 = n50523 & n50524;
  assign n46616 = n50525 ^ n50526;
  assign n50544 = n50553 & n50554;
  assign n50337 = n50280 & n293;
  assign n50336 = ~n50280;
  assign n50376 = n50381 & n50382;
  assign n50340 = ~n50383;
  assign n46182 = n50384 ^ n50385;
  assign n50375 = ~n50393;
  assign n50379 = ~n50405;
  assign n50408 = n50411 & n50412;
  assign n50304 = n50432 ^ n50433;
  assign n50358 = n50433 & n50432;
  assign n50363 = n50468 ^ n50469;
  assign n50466 = ~n50486;
  assign n50488 = n50511 & n50512;
  assign n50492 = n46616 & n49227;
  assign n50493 = n46616 & n49178;
  assign n50494 = n50399 & n50441;
  assign n50495 = n46616 & n47923;
  assign n50489 = ~n50399;
  assign n46650 = ~n46616;
  assign n50527 = ~n50544;
  assign n50329 = n50336 & n2430;
  assign n50250 = ~n50337;
  assign n50342 = n46182 & n48609;
  assign n50343 = n46182 & n47336;
  assign n50330 = n50375 & n50333;
  assign n50301 = ~n50376;
  assign n50357 = n50375 & n50331;
  assign n46224 = ~n46182;
  assign n50338 = n50379 & n50380;
  assign n50386 = ~n50408;
  assign n50394 = n50304 & n47292;
  assign n50395 = ~n50304;
  assign n50361 = ~n50358;
  assign n50438 = n50363 & n5391;
  assign n50439 = ~n50363;
  assign n50434 = n50466 & n50467;
  assign n50470 = ~n50488;
  assign n50480 = n50489 & n50490;
  assign n50481 = n46650 & n50491;
  assign n49229 = ~n50492;
  assign n50472 = ~n50493;
  assign n50443 = ~n50494;
  assign n49195 = ~n50495;
  assign n50496 = n50527 & n50528;
  assign n50294 = ~n50329;
  assign n48568 = n50330 ^ n50331;
  assign n50303 = n50338 ^ n50339;
  assign n50313 = ~n50342;
  assign n48626 = ~n50343;
  assign n50332 = ~n50357;
  assign n50341 = ~n50338;
  assign n50344 = n50386 & n50387;
  assign n50346 = ~n50394;
  assign n50388 = n50395 & n47248;
  assign n50396 = n50434 ^ n50435;
  assign n50365 = ~n50438;
  assign n50422 = n50439 & n148;
  assign n50436 = ~n50434;
  assign n50440 = n50470 & n50471;
  assign n50321 = n50472 & n50473;
  assign n50402 = ~n50480;
  assign n49253 = ~n50481;
  assign n50459 = n50496 ^ n47884;
  assign n50497 = ~n50496;
  assign n50202 = n50302 ^ n50303;
  assign n50218 = n50313 & n50314;
  assign n48598 = ~n48568;
  assign n50315 = n50332 & n50333;
  assign n50328 = n50340 & n50341;
  assign n50305 = n50344 ^ n47248;
  assign n50345 = ~n50344;
  assign n50307 = ~n50388;
  assign n50359 = n149 ^ n50396;
  assign n50320 = ~n50422;
  assign n50421 = n50436 & n50437;
  assign n50400 = n50440 ^ n50441;
  assign n50445 = n50321 & n50451;
  assign n50442 = ~n50440;
  assign n50444 = ~n50321;
  assign n46565 = n50459 ^ n50460;
  assign n50482 = n50497 & n50498;
  assign n50255 = n50202 & n2338;
  assign n50254 = ~n50202;
  assign n50278 = n50218 & n50295;
  assign n50277 = ~n50218;
  assign n46091 = n50304 ^ n50305;
  assign n50279 = ~n50315;
  assign n50300 = ~n50328;
  assign n50334 = n50345 & n50346;
  assign n50223 = n50358 ^ n50359;
  assign n50360 = ~n50359;
  assign n50284 = n50399 ^ n50400;
  assign n50397 = ~n50421;
  assign n50423 = n50442 & n50443;
  assign n50424 = n50444 & n50369;
  assign n50425 = n46565 & n49183;
  assign n50371 = ~n50445;
  assign n50426 = n46565 & n49114;
  assign n50427 = n46565 & n47884;
  assign n46606 = ~n46565;
  assign n50461 = ~n50482;
  assign n50246 = n50254 & n292;
  assign n50217 = ~n50255;
  assign n50256 = n50277 & n50251;
  assign n50257 = n46091 & n48553;
  assign n50247 = ~n50278;
  assign n50258 = n46091 & n47292;
  assign n50260 = n46091 & n48629;
  assign n50235 = n50279 ^ n50280;
  assign n50276 = n50294 & n50279;
  assign n46111 = ~n46091;
  assign n50296 = n50300 & n50301;
  assign n50306 = ~n50334;
  assign n50316 = n50223 & n47232;
  assign n50317 = ~n50223;
  assign n50281 = n50360 & n50361;
  assign n50366 = n50284 & n5352;
  assign n50367 = ~n50284;
  assign n50362 = n50397 & n50398;
  assign n50401 = ~n50423;
  assign n50324 = ~n50424;
  assign n49186 = ~n50425;
  assign n50403 = ~n50426;
  assign n49143 = ~n50427;
  assign n50409 = n46606 & n50428;
  assign n50429 = n50461 & n50462;
  assign n50198 = n293 ^ n50235;
  assign n50169 = ~n50246;
  assign n50221 = ~n50256;
  assign n50237 = ~n50257;
  assign n48590 = ~n50258;
  assign n50252 = n46111 & n50259;
  assign n48632 = ~n50260;
  assign n50249 = ~n50276;
  assign n50248 = ~n50296;
  assign n50261 = n50306 & n50307;
  assign n50225 = ~n50316;
  assign n50308 = n50317 & n47251;
  assign n50318 = n50362 ^ n50363;
  assign n50275 = ~n50366;
  assign n50348 = n50367 & n147;
  assign n50364 = ~n50362;
  assign n50368 = n50401 & n50402;
  assign n50231 = n50403 & n50404;
  assign n49207 = ~n50409;
  assign n50389 = n50429 ^ n47842;
  assign n50430 = ~n50429;
  assign n48541 = n50198 ^ n48568;
  assign n50200 = ~n50198;
  assign n50130 = n50237 & n50238;
  assign n50236 = n50247 & n50248;
  assign n50239 = n50249 & n50250;
  assign n50219 = n50248 ^ n50251;
  assign n48648 = ~n50252;
  assign n50222 = n50261 ^ n47251;
  assign n50262 = ~n50261;
  assign n50263 = ~n50308;
  assign n50282 = n148 ^ n50318;
  assign n50244 = ~n50348;
  assign n50347 = n50364 & n50365;
  assign n50322 = n50368 ^ n50369;
  assign n50374 = n50231 & n50288;
  assign n50370 = ~n50368;
  assign n50372 = ~n50231;
  assign n46512 = n50389 ^ n50390;
  assign n50410 = n50430 & n50431;
  assign n50112 = ~n48541;
  assign n50107 = n50200 & n48598;
  assign n50133 = n50218 ^ n50219;
  assign n50203 = n50130 & n50173;
  assign n50194 = ~n50130;
  assign n45997 = n50222 ^ n50223;
  assign n50220 = ~n50236;
  assign n50201 = ~n50239;
  assign n50245 = n50262 & n50263;
  assign n50143 = n50281 ^ n50282;
  assign n50196 = n50282 & n50281;
  assign n50207 = n50321 ^ n50322;
  assign n50319 = ~n50347;
  assign n50349 = n50370 & n50371;
  assign n50350 = n50372 & n50373;
  assign n50351 = n46512 & n49069;
  assign n50290 = ~n50374;
  assign n50352 = n46512 & n47842;
  assign n46553 = ~n46512;
  assign n50391 = ~n50410;
  assign n50110 = ~n50107;
  assign n50170 = n50133 & n2210;
  assign n50179 = n50194 & n50195;
  assign n50171 = ~n50133;
  assign n50152 = n50201 ^ n50202;
  assign n50180 = n45997 & n48516;
  assign n50174 = ~n50203;
  assign n50181 = n45997 & n47251;
  assign n50199 = n50217 & n50201;
  assign n50172 = n50220 & n50221;
  assign n46037 = ~n45997;
  assign n50224 = ~n50245;
  assign n50240 = n50143 & n47202;
  assign n50241 = ~n50143;
  assign n50205 = ~n50196;
  assign n50286 = n50207 & n146;
  assign n50285 = ~n50207;
  assign n50283 = n50319 & n50320;
  assign n50323 = ~n50349;
  assign n50234 = ~n50350;
  assign n50325 = ~n50351;
  assign n49082 = ~n50352;
  assign n50353 = n50391 & n50392;
  assign n50108 = n292 ^ n50152;
  assign n50134 = ~n50170;
  assign n50153 = n50171 & n291;
  assign n50131 = n50172 ^ n50173;
  assign n50137 = ~n50179;
  assign n50154 = ~n50180;
  assign n48538 = ~n50181;
  assign n50168 = ~n50199;
  assign n50175 = ~n50172;
  assign n50182 = n50224 & n50225;
  assign n50146 = ~n50240;
  assign n50226 = n50241 & n47195;
  assign n50242 = n50283 ^ n50284;
  assign n50265 = n50285 & n5311;
  assign n50161 = ~n50286;
  assign n50274 = ~n50283;
  assign n50287 = n50323 & n50324;
  assign n50162 = n50325 & n50326;
  assign n46422 = n50353 ^ n50354;
  assign n50355 = ~n50353;
  assign n48499 = n50107 ^ n50108;
  assign n50049 = n50130 ^ n50131;
  assign n50109 = ~n50108;
  assign n50082 = ~n50153;
  assign n50046 = n50154 & n50155;
  assign n50132 = n50168 & n50169;
  assign n50156 = n50174 & n50175;
  assign n50144 = n50182 ^ n47195;
  assign n50183 = ~n50182;
  assign n50184 = ~n50226;
  assign n50197 = n147 ^ n50242;
  assign n50209 = ~n50265;
  assign n50264 = n50274 & n50275;
  assign n50232 = n50287 ^ n50288;
  assign n50293 = n50162 & n50213;
  assign n50289 = ~n50287;
  assign n50291 = ~n50162;
  assign n50309 = n46422 & n50327;
  assign n46498 = ~n46422;
  assign n50335 = n50355 & n50356;
  assign n50079 = n50049 & n2109;
  assign n50010 = ~n48499;
  assign n50042 = n50109 & n50110;
  assign n50080 = ~n50049;
  assign n50078 = n50132 ^ n50133;
  assign n50114 = n50046 & n50138;
  assign n45936 = n50143 ^ n50144;
  assign n50113 = ~n50046;
  assign n50135 = ~n50132;
  assign n50136 = ~n50156;
  assign n50176 = n50183 & n50184;
  assign n50055 = n50196 ^ n50197;
  assign n50204 = ~n50197;
  assign n50120 = n50231 ^ n50232;
  assign n50243 = ~n50264;
  assign n50266 = n50289 & n50290;
  assign n50267 = n50291 & n50292;
  assign n50215 = ~n50293;
  assign n49099 = ~n50309;
  assign n50297 = n46498 & n49022;
  assign n50298 = n46498 & n47736;
  assign n50299 = n46498 & n50310;
  assign n50311 = ~n50335;
  assign n50043 = n291 ^ n50078;
  assign n50044 = ~n50079;
  assign n50067 = n50080 & n290;
  assign n50091 = n45936 & n50112;
  assign n50092 = n50113 & n50084;
  assign n50085 = ~n50114;
  assign n50093 = n45936 & n48463;
  assign n50094 = n45936 & n47195;
  assign n50111 = n50134 & n50135;
  assign n50083 = n50136 & n50137;
  assign n45963 = ~n45936;
  assign n50145 = ~n50176;
  assign n50157 = n50055 & n47166;
  assign n50158 = ~n50055;
  assign n50115 = n50204 & n50205;
  assign n50210 = n50120 & n5261;
  assign n50211 = ~n50120;
  assign n50206 = n50243 & n50244;
  assign n50233 = ~n50266;
  assign n50165 = ~n50267;
  assign n50268 = ~n50297;
  assign n49078 = ~n50298;
  assign n49120 = ~n50299;
  assign n50270 = n50311 & n50312;
  assign n48461 = n50042 ^ n50043;
  assign n49950 = n50043 & n50042;
  assign n49994 = ~n50067;
  assign n50047 = n50083 ^ n50084;
  assign n50087 = n45963 & n48541;
  assign n48543 = ~n50091;
  assign n50051 = ~n50092;
  assign n50068 = ~n50093;
  assign n48509 = ~n50094;
  assign n50081 = ~n50111;
  assign n50086 = ~n50083;
  assign n50095 = n50145 & n50146;
  assign n50097 = ~n50157;
  assign n50147 = n50158 & n47150;
  assign n50118 = ~n50115;
  assign n50159 = n50206 ^ n50207;
  assign n50122 = ~n50210;
  assign n50186 = n50211 & n145;
  assign n50208 = ~n50206;
  assign n50212 = n50233 & n50234;
  assign n50040 = n50268 & n50269;
  assign n49117 = n49120 & n49099;
  assign n50227 = n50270 ^ n50271;
  assign n50272 = ~n50270;
  assign n49923 = ~n48461;
  assign n49953 = ~n49950;
  assign n49955 = n50046 ^ n50047;
  assign n49958 = n50068 & n50069;
  assign n50048 = n50081 & n50082;
  assign n50066 = n50085 & n50086;
  assign n48564 = ~n50087;
  assign n50056 = n50095 ^ n47150;
  assign n50096 = ~n50095;
  assign n50058 = ~n50147;
  assign n50116 = n146 ^ n50159;
  assign n50074 = ~n50186;
  assign n50185 = n50208 & n50209;
  assign n50163 = n50212 ^ n50213;
  assign n50214 = ~n50212;
  assign n46435 = n50227 ^ n47689;
  assign n50228 = n50227 & n47719;
  assign n50253 = n50272 & n50273;
  assign n49996 = n49955 & n289;
  assign n49995 = ~n49955;
  assign n49992 = n50048 ^ n50049;
  assign n50032 = n49958 & n50052;
  assign n50031 = ~n49958;
  assign n45883 = n50055 ^ n50056;
  assign n50050 = ~n50066;
  assign n50045 = ~n50048;
  assign n50077 = n50096 & n50097;
  assign n49969 = n50115 ^ n50116;
  assign n50117 = ~n50116;
  assign n50038 = n50162 ^ n50163;
  assign n50160 = ~n50185;
  assign n50187 = n50214 & n50215;
  assign n50188 = n46435 & n49004;
  assign n50189 = n46435 & n50216;
  assign n46357 = ~n46435;
  assign n49020 = ~n50228;
  assign n50229 = ~n50253;
  assign n49951 = n290 ^ n49992;
  assign n49978 = n49995 & n2069;
  assign n49905 = ~n49996;
  assign n50013 = n45883 & n48455;
  assign n50011 = n45883 & n48499;
  assign n50012 = n50031 & n49999;
  assign n50000 = ~n50032;
  assign n50014 = n45883 & n47166;
  assign n50030 = n50044 & n50045;
  assign n49998 = n50050 & n50051;
  assign n45909 = ~n45883;
  assign n50057 = ~n50077;
  assign n50070 = n49969 & n47110;
  assign n50071 = ~n49969;
  assign n50033 = n50117 & n50118;
  assign n50123 = n50038 & n5208;
  assign n50124 = ~n50038;
  assign n50119 = n50160 & n50161;
  assign n50164 = ~n50187;
  assign n50166 = ~n50188;
  assign n50177 = n46357 & n49073;
  assign n49057 = ~n50189;
  assign n50190 = n50229 & n50230;
  assign n48422 = n49950 ^ n49951;
  assign n49952 = ~n49951;
  assign n49956 = ~n49978;
  assign n49959 = n49998 ^ n49999;
  assign n49997 = n45909 & n50010;
  assign n48503 = ~n50011;
  assign n49961 = ~n50012;
  assign n49979 = ~n50013;
  assign n48471 = ~n50014;
  assign n49993 = ~n50030;
  assign n50001 = ~n49998;
  assign n50015 = n50057 & n50058;
  assign n49971 = ~n50070;
  assign n50059 = n50071 & n47140;
  assign n50036 = ~n50033;
  assign n50072 = n50119 ^ n50120;
  assign n50029 = ~n50123;
  assign n50099 = n50124 & n144;
  assign n50121 = ~n50119;
  assign n50139 = n50164 & n50165;
  assign n50004 = n50166 & n50167;
  assign n49075 = ~n50177;
  assign n50148 = n50190 ^ n50191;
  assign n50192 = ~n50190;
  assign n49841 = ~n48422;
  assign n49868 = n49952 & n49953;
  assign n49871 = n49958 ^ n49959;
  assign n49874 = n49979 & n49980;
  assign n49954 = n49993 & n49994;
  assign n48528 = ~n49997;
  assign n49981 = n50000 & n50001;
  assign n49968 = n50015 ^ n47140;
  assign n50016 = ~n50015;
  assign n50017 = ~n50059;
  assign n50034 = n145 ^ n50072;
  assign n49986 = ~n50099;
  assign n50098 = n50121 & n50122;
  assign n50127 = n50139 & n50140;
  assign n50129 = n50004 & n50141;
  assign n50125 = ~n50139;
  assign n50128 = ~n50004;
  assign n46321 = n47649 ^ n50148;
  assign n50149 = ~n50148;
  assign n50178 = n50192 & n50193;
  assign n49907 = n49871 & n288;
  assign n49906 = ~n49871;
  assign n49903 = n49954 ^ n49955;
  assign n49941 = n49874 & n49962;
  assign n49940 = ~n49874;
  assign n45842 = n49968 ^ n49969;
  assign n49957 = ~n49954;
  assign n49960 = ~n49981;
  assign n50002 = n50016 & n50017;
  assign n49884 = n50033 ^ n50034;
  assign n50035 = ~n50034;
  assign n50073 = ~n50098;
  assign n50100 = n50125 & n50126;
  assign n50076 = ~n50127;
  assign n50101 = n50128 & n49964;
  assign n50006 = ~n50129;
  assign n50103 = n46321 & n49015;
  assign n46361 = ~n46321;
  assign n50142 = n50149 & n47716;
  assign n50150 = ~n50178;
  assign n49869 = n289 ^ n49903;
  assign n49891 = n49906 & n2009;
  assign n49821 = ~n49907;
  assign n49922 = n45842 & n48461;
  assign n49924 = n49940 & n49910;
  assign n49925 = n45842 & n48381;
  assign n49911 = ~n49941;
  assign n49926 = n45842 & n47140;
  assign n49939 = n49956 & n49957;
  assign n49909 = n49960 & n49961;
  assign n45853 = ~n45842;
  assign n49970 = ~n50002;
  assign n49983 = n49884 & n47081;
  assign n49982 = ~n49884;
  assign n49942 = n50035 & n50036;
  assign n50037 = n50073 & n50074;
  assign n50075 = n50076 & n50040;
  assign n50054 = ~n50100;
  assign n49966 = ~n50101;
  assign n50088 = n46361 & n48910;
  assign n50089 = n46361 & n50102;
  assign n49038 = ~n50103;
  assign n48980 = ~n50142;
  assign n50104 = n50150 & n50151;
  assign n48387 = n49868 ^ n49869;
  assign n49784 = n49869 & n49868;
  assign n49873 = ~n49891;
  assign n49875 = n49909 ^ n49910;
  assign n48465 = ~n49922;
  assign n49908 = n45853 & n49923;
  assign n49877 = ~n49924;
  assign n49892 = ~n49925;
  assign n48430 = ~n49926;
  assign n49904 = ~n49939;
  assign n49912 = ~n49909;
  assign n49927 = n49970 & n49971;
  assign n49972 = n49982 & n47075;
  assign n49929 = ~n49983;
  assign n49984 = n50037 ^ n50038;
  assign n50028 = ~n50037;
  assign n50053 = ~n50075;
  assign n50039 = n50054 & n50076;
  assign n50060 = ~n50088;
  assign n49018 = ~n50089;
  assign n50063 = n50104 ^ n47602;
  assign n50105 = ~n50104;
  assign n49770 = ~n48387;
  assign n49787 = n49874 ^ n49875;
  assign n49790 = n49892 & n49893;
  assign n49870 = n49904 & n49905;
  assign n48483 = ~n49908;
  assign n49894 = n49911 & n49912;
  assign n49883 = n49927 ^ n47081;
  assign n49928 = ~n49927;
  assign n49886 = ~n49972;
  assign n49943 = n144 ^ n49984;
  assign n50018 = n50028 & n50029;
  assign n49896 = n50039 ^ n50040;
  assign n50003 = n50053 & n50054;
  assign n49879 = n50060 & n50061;
  assign n46240 = n50062 ^ n50063;
  assign n50090 = n50105 & n50106;
  assign n49823 = n49787 & n303;
  assign n49822 = ~n49787;
  assign n49819 = n49870 ^ n49871;
  assign n49857 = n49790 & n49878;
  assign n49856 = ~n49790;
  assign n45788 = n49883 ^ n49884;
  assign n49872 = ~n49870;
  assign n49876 = ~n49894;
  assign n49913 = n49928 & n49929;
  assign n49799 = n49942 ^ n49943;
  assign n49944 = ~n49943;
  assign n49988 = n49896 & n159;
  assign n49963 = n50003 ^ n50004;
  assign n49985 = ~n50018;
  assign n49987 = ~n49896;
  assign n50005 = ~n50003;
  assign n50020 = n49879 & n50041;
  assign n50021 = n46240 & n48928;
  assign n50022 = n46240 & n47602;
  assign n50023 = n46240 & n48982;
  assign n50019 = ~n49879;
  assign n46306 = ~n46240;
  assign n50064 = ~n50090;
  assign n49785 = n288 ^ n49819;
  assign n49808 = n49822 & n1922;
  assign n49743 = ~n49823;
  assign n49842 = n45788 & n48422;
  assign n49843 = n49856 & n49826;
  assign n49828 = ~n49857;
  assign n49855 = n49872 & n49873;
  assign n49825 = n49876 & n49877;
  assign n45809 = ~n45788;
  assign n49885 = ~n49913;
  assign n49858 = n49944 & n49942;
  assign n49861 = n49963 ^ n49964;
  assign n49945 = n49985 & n49986;
  assign n49973 = n49987 & n5179;
  assign n49898 = ~n49988;
  assign n49989 = n50005 & n50006;
  assign n50007 = n50019 & n49917;
  assign n49919 = ~n50020;
  assign n49990 = ~n50021;
  assign n48946 = ~n50022;
  assign n48984 = ~n50023;
  assign n50008 = n46306 & n50024;
  assign n50025 = n50064 & n50065;
  assign n49649 = n49784 ^ n49785;
  assign n49705 = n49785 & n49784;
  assign n49788 = ~n49808;
  assign n49791 = n49825 ^ n49826;
  assign n49824 = n45809 & n49841;
  assign n48445 = ~n49842;
  assign n49793 = ~n49843;
  assign n49829 = n45809 & n48341;
  assign n49830 = n45809 & n47081;
  assign n49820 = ~n49855;
  assign n49827 = ~n49825;
  assign n49844 = n49885 & n49886;
  assign n49915 = n49861 & n158;
  assign n49895 = n159 ^ n49945;
  assign n49914 = ~n49861;
  assign n49946 = ~n49945;
  assign n49947 = ~n49973;
  assign n49965 = ~n49989;
  assign n49794 = n49990 & n49991;
  assign n49882 = ~n50007;
  assign n49001 = ~n50008;
  assign n49975 = n50025 ^ n47552;
  assign n50026 = ~n50025;
  assign n48346 = ~n49649;
  assign n49708 = n49790 ^ n49791;
  assign n49786 = n49820 & n49821;
  assign n48425 = ~n49824;
  assign n49809 = n49827 & n49828;
  assign n49800 = ~n49829;
  assign n48385 = ~n49830;
  assign n49798 = n49844 ^ n47049;
  assign n49846 = n49844 & n47049;
  assign n49845 = ~n49844;
  assign n49859 = n49895 ^ n49896;
  assign n49899 = n49914 & n5130;
  assign n49814 = ~n49915;
  assign n49930 = n49946 & n49947;
  assign n49916 = n49965 & n49966;
  assign n49949 = n49794 & n49967;
  assign n49948 = ~n49794;
  assign n46161 = n49974 ^ n49975;
  assign n50009 = n50026 & n50027;
  assign n49745 = n49708 & n302;
  assign n49744 = ~n49708;
  assign n49740 = n49786 ^ n49787;
  assign n45748 = n49798 ^ n49799;
  assign n49703 = n49800 & n49801;
  assign n49789 = ~n49786;
  assign n49792 = ~n49809;
  assign n49831 = n49845 & n47025;
  assign n49810 = ~n49846;
  assign n49832 = n49858 ^ n49859;
  assign n49774 = n49859 & n49858;
  assign n49863 = ~n49899;
  assign n49880 = n49916 ^ n49917;
  assign n49897 = ~n49930;
  assign n49918 = ~n49916;
  assign n49931 = n49948 & n49836;
  assign n49932 = n46161 & n48882;
  assign n49838 = ~n49949;
  assign n49933 = n46161 & n47552;
  assign n49934 = n46161 & n48939;
  assign n46227 = ~n46161;
  assign n49976 = ~n50009;
  assign n49706 = n303 ^ n49740;
  assign n49726 = n49744 & n1874;
  assign n49669 = ~n49745;
  assign n49759 = n45748 & n49770;
  assign n49762 = n45748 & n48300;
  assign n49763 = n49703 & n49747;
  assign n49764 = n45748 & n47049;
  assign n49771 = n49788 & n49789;
  assign n49746 = n49792 & n49793;
  assign n49760 = ~n49703;
  assign n45763 = ~n45748;
  assign n49802 = n49810 & n49799;
  assign n49773 = ~n49831;
  assign n49811 = n49832 & n47015;
  assign n49693 = ~n49832;
  assign n49777 = n49879 ^ n49880;
  assign n49860 = n49897 & n49898;
  assign n49900 = n49918 & n49919;
  assign n49797 = ~n49931;
  assign n49901 = ~n49932;
  assign n48902 = ~n49933;
  assign n48942 = ~n49934;
  assign n49920 = n46227 & n49935;
  assign n49936 = n49976 & n49977;
  assign n48306 = n49705 ^ n49706;
  assign n49630 = n49706 & n49705;
  assign n49710 = ~n49726;
  assign n49704 = n49746 ^ n49747;
  assign n48389 = ~n49759;
  assign n49741 = n45763 & n48387;
  assign n49748 = n49760 & n49761;
  assign n49727 = ~n49762;
  assign n49730 = ~n49763;
  assign n48345 = ~n49764;
  assign n49742 = ~n49771;
  assign n49729 = ~n49746;
  assign n49772 = ~n49802;
  assign n49803 = n49693 & n46987;
  assign n49733 = ~n49811;
  assign n49834 = n49777 & n157;
  assign n49812 = n49860 ^ n49861;
  assign n49833 = ~n49777;
  assign n49862 = ~n49860;
  assign n49881 = ~n49900;
  assign n49712 = n49901 & n49902;
  assign n48965 = ~n49920;
  assign n49888 = n49936 ^ n47505;
  assign n49937 = ~n49936;
  assign n49597 = ~n48306;
  assign n49633 = n49703 ^ n49704;
  assign n49629 = ~n49630;
  assign n49614 = n49727 & n49728;
  assign n49718 = n49729 & n49730;
  assign n48404 = ~n49741;
  assign n49707 = n49742 & n49743;
  assign n49689 = ~n49748;
  assign n49731 = n49772 & n49773;
  assign n49695 = ~n49803;
  assign n49775 = n158 ^ n49812;
  assign n49815 = n49833 & n5088;
  assign n49737 = ~n49834;
  assign n49847 = n49862 & n49863;
  assign n49835 = n49881 & n49882;
  assign n49866 = n49712 & n49753;
  assign n49864 = ~n49712;
  assign n46082 = n49887 ^ n49888;
  assign n49921 = n49937 & n49938;
  assign n49670 = n49633 & n1851;
  assign n49671 = ~n49633;
  assign n49667 = n49707 ^ n49708;
  assign n49691 = n49614 & n49711;
  assign n49690 = ~n49614;
  assign n49688 = ~n49718;
  assign n49709 = ~n49707;
  assign n49692 = n49731 ^ n47015;
  assign n49732 = ~n49731;
  assign n49749 = n49774 ^ n49775;
  assign n49696 = n49775 & n49774;
  assign n49779 = ~n49815;
  assign n49795 = n49835 ^ n49836;
  assign n49813 = ~n49847;
  assign n49837 = ~n49835;
  assign n49848 = n49864 & n49865;
  assign n49849 = n46082 & n48846;
  assign n49755 = ~n49866;
  assign n49850 = n46082 & n47505;
  assign n49851 = n46082 & n49867;
  assign n46149 = ~n46082;
  assign n49889 = ~n49921;
  assign n49631 = n302 ^ n49667;
  assign n49634 = ~n49670;
  assign n49650 = n49671 & n301;
  assign n49651 = n49688 & n49689;
  assign n49679 = n49690 & n49652;
  assign n49654 = ~n49691;
  assign n45723 = n49692 ^ n49693;
  assign n49687 = n49709 & n49710;
  assign n49719 = n49732 & n49733;
  assign n49734 = n49749 & n46949;
  assign n49618 = ~n49749;
  assign n49699 = n49794 ^ n49795;
  assign n49776 = n49813 & n49814;
  assign n49816 = n49837 & n49838;
  assign n49715 = ~n49848;
  assign n49817 = ~n49849;
  assign n48863 = ~n49850;
  assign n49839 = n46149 & n48903;
  assign n48906 = ~n49851;
  assign n49852 = n49889 & n49890;
  assign n48264 = n49630 ^ n49631;
  assign n49628 = ~n49631;
  assign n49599 = ~n49650;
  assign n49615 = n49651 ^ n49652;
  assign n49648 = n45723 & n48346;
  assign n49655 = n45723 & n48259;
  assign n49656 = n45723 & n47015;
  assign n49653 = ~n49651;
  assign n49617 = ~n49679;
  assign n45710 = ~n45723;
  assign n49668 = ~n49687;
  assign n49694 = ~n49719;
  assign n49720 = n49618 & n46969;
  assign n49659 = ~n49734;
  assign n49751 = n49699 & n156;
  assign n49735 = n49776 ^ n49777;
  assign n49750 = ~n49699;
  assign n49778 = ~n49776;
  assign n49796 = ~n49816;
  assign n49638 = n49817 & n49818;
  assign n48923 = ~n49839;
  assign n49804 = n49852 ^ n47462;
  assign n49853 = ~n49852;
  assign n49535 = ~n48264;
  assign n49565 = n49614 ^ n49615;
  assign n49560 = n49628 & n49629;
  assign n48349 = ~n49648;
  assign n49642 = n45710 & n49649;
  assign n49643 = n49653 & n49654;
  assign n49636 = ~n49655;
  assign n48302 = ~n49656;
  assign n49632 = n49668 & n49669;
  assign n49657 = n49694 & n49695;
  assign n49621 = ~n49720;
  assign n49697 = n157 ^ n49735;
  assign n49738 = n49750 & n5043;
  assign n49664 = ~n49751;
  assign n49765 = n49778 & n49779;
  assign n49752 = n49796 & n49797;
  assign n49782 = n49638 & n49675;
  assign n49780 = ~n49638;
  assign n46011 = n49804 ^ n49805;
  assign n49840 = n49853 & n49854;
  assign n49582 = n49565 & n300;
  assign n49581 = ~n49565;
  assign n49563 = ~n49560;
  assign n49596 = n49632 ^ n49633;
  assign n49542 = n49636 & n49637;
  assign n48369 = ~n49642;
  assign n49616 = ~n49643;
  assign n49635 = ~n49632;
  assign n49619 = n49657 ^ n46949;
  assign n49658 = ~n49657;
  assign n49550 = n49696 ^ n49697;
  assign n49611 = n49697 & n49696;
  assign n49701 = ~n49738;
  assign n49713 = n49752 ^ n49753;
  assign n49736 = ~n49765;
  assign n49754 = ~n49752;
  assign n49766 = n49780 & n49781;
  assign n49677 = ~n49782;
  assign n49767 = n46011 & n49783;
  assign n46063 = ~n46011;
  assign n49806 = ~n49840;
  assign n49574 = n49581 & n1797;
  assign n49523 = ~n49582;
  assign n49561 = n301 ^ n49596;
  assign n49601 = n49542 & n49608;
  assign n49600 = ~n49542;
  assign n49609 = n49616 & n49617;
  assign n45672 = n49618 ^ n49619;
  assign n49613 = n49634 & n49635;
  assign n49644 = n49658 & n49659;
  assign n49661 = n49550 & n46909;
  assign n49660 = ~n49550;
  assign n49623 = ~n49611;
  assign n49625 = n49712 ^ n49713;
  assign n49698 = n49736 & n49737;
  assign n49739 = n49754 & n49755;
  assign n49641 = ~n49766;
  assign n49756 = n46063 & n48807;
  assign n49757 = n46063 & n47462;
  assign n49758 = n46063 & n48859;
  assign n48865 = ~n49767;
  assign n49768 = n49806 & n49807;
  assign n49464 = n49560 ^ n49561;
  assign n49549 = ~n49574;
  assign n49562 = ~n49561;
  assign n49580 = n45672 & n49597;
  assign n49583 = n49600 & n49577;
  assign n49584 = n45672 & n48242;
  assign n49575 = ~n49601;
  assign n49585 = n45672 & n46949;
  assign n49576 = ~n49609;
  assign n45690 = ~n45672;
  assign n49598 = ~n49613;
  assign n49620 = ~n49644;
  assign n49645 = n49660 & n46938;
  assign n49588 = ~n49661;
  assign n49672 = n49625 & n5010;
  assign n49662 = n49698 ^ n49699;
  assign n49673 = ~n49625;
  assign n49700 = ~n49698;
  assign n49714 = ~n49739;
  assign n49721 = ~n49756;
  assign n48822 = ~n49757;
  assign n48891 = ~n49758;
  assign n45973 = n49768 ^ n49769;
  assign n48222 = ~n49464;
  assign n49504 = n49562 & n49563;
  assign n49566 = n49575 & n49576;
  assign n49543 = n49576 ^ n49577;
  assign n49573 = n45690 & n48306;
  assign n48308 = ~n49580;
  assign n49545 = ~n49583;
  assign n49567 = ~n49584;
  assign n48261 = ~n49585;
  assign n49564 = n49598 & n49599;
  assign n49586 = n49620 & n49621;
  assign n49553 = ~n49645;
  assign n49612 = n156 ^ n49662;
  assign n49627 = ~n49672;
  assign n49665 = n49673 & n155;
  assign n49680 = n49700 & n49701;
  assign n49674 = n49714 & n49715;
  assign n49569 = n49721 & n49722;
  assign n49681 = n49723 ^ n45973;
  assign n48834 = ~n45973;
  assign n49489 = n49542 ^ n49543;
  assign n49534 = n49564 ^ n49565;
  assign n49544 = ~n49566;
  assign n49480 = n49567 & n49568;
  assign n48330 = ~n49573;
  assign n49548 = ~n49564;
  assign n49551 = n49586 ^ n46909;
  assign n49587 = ~n49586;
  assign n49493 = n49611 ^ n49612;
  assign n49622 = ~n49612;
  assign n49593 = ~n49665;
  assign n49639 = n49674 ^ n49675;
  assign n49663 = ~n49680;
  assign n48849 = n49681 ^ n49682;
  assign n49676 = ~n49674;
  assign n49684 = n49569 & n49702;
  assign n49683 = ~n49569;
  assign n49716 = n48834 & n49724;
  assign n49717 = n48834 & n49725;
  assign n49511 = n49489 & n1764;
  assign n49505 = n300 ^ n49534;
  assign n49512 = ~n49489;
  assign n49513 = n49544 & n49545;
  assign n49537 = n49480 & n49546;
  assign n49541 = n49548 & n49549;
  assign n49536 = ~n49480;
  assign n45633 = n49550 ^ n49551;
  assign n49578 = n49587 & n49588;
  assign n49590 = n49493 & n46866;
  assign n49589 = ~n49493;
  assign n49554 = n49622 & n49623;
  assign n49557 = n49638 ^ n49639;
  assign n49624 = n49663 & n49664;
  assign n49666 = n49676 & n49677;
  assign n49678 = n49683 & n49605;
  assign n49607 = ~n49684;
  assign n49685 = ~n49716;
  assign n48819 = ~n49717;
  assign n48204 = n49504 ^ n49505;
  assign n49436 = n49505 & n49504;
  assign n49487 = ~n49511;
  assign n49506 = n49512 & n299;
  assign n49481 = n49513 ^ n49514;
  assign n49521 = n45633 & n49535;
  assign n49516 = ~n49513;
  assign n49524 = n49536 & n49514;
  assign n49515 = ~n49537;
  assign n49522 = ~n49541;
  assign n45629 = ~n45633;
  assign n49552 = ~n49578;
  assign n49579 = n49589 & n46901;
  assign n49495 = ~n49590;
  assign n49602 = n49557 & n4987;
  assign n49591 = n49624 ^ n49625;
  assign n49603 = ~n49557;
  assign n49626 = ~n49624;
  assign n49640 = ~n49666;
  assign n49572 = ~n49678;
  assign n49646 = n49685 & n49686;
  assign n49434 = n49480 ^ n49481;
  assign n49424 = ~n48204;
  assign n49447 = ~n49436;
  assign n49466 = ~n49506;
  assign n49507 = n49515 & n49516;
  assign n49510 = n45629 & n48264;
  assign n48290 = ~n49521;
  assign n49488 = n49522 & n49523;
  assign n49484 = ~n49524;
  assign n49517 = n45629 & n48174;
  assign n49518 = n45629 & n46909;
  assign n49525 = n49552 & n49553;
  assign n49527 = ~n49579;
  assign n49555 = n155 ^ n49591;
  assign n49559 = ~n49602;
  assign n49594 = n49603 & n154;
  assign n49610 = n49626 & n49627;
  assign n49604 = n49640 & n49641;
  assign n49509 = n49646 ^ n49647;
  assign n49455 = n49434 & n298;
  assign n49454 = ~n49434;
  assign n49462 = n49488 ^ n49489;
  assign n49483 = ~n49507;
  assign n48267 = ~n49510;
  assign n49486 = ~n49488;
  assign n49490 = ~n49517;
  assign n48226 = ~n49518;
  assign n49492 = n49525 ^ n46901;
  assign n49526 = ~n49525;
  assign n49439 = n49554 ^ n49555;
  assign n49496 = n49555 & n49554;
  assign n49532 = ~n49594;
  assign n49570 = n49604 ^ n49605;
  assign n49592 = ~n49610;
  assign n49606 = ~n49604;
  assign n49448 = n49454 & n1703;
  assign n49407 = ~n49455;
  assign n49437 = n299 ^ n49462;
  assign n49457 = n49483 & n49484;
  assign n49482 = n49486 & n49487;
  assign n49432 = n49490 & n49491;
  assign n45563 = n49492 ^ n49493;
  assign n49519 = n49526 & n49527;
  assign n49529 = n49439 & n46849;
  assign n49528 = ~n49439;
  assign n49499 = ~n49496;
  assign n49501 = n49569 ^ n49570;
  assign n49556 = n49592 & n49593;
  assign n49595 = n49606 & n49607;
  assign n48160 = n49436 ^ n49437;
  assign n49383 = n49437 & n49447;
  assign n49430 = ~n49448;
  assign n49433 = n49457 ^ n49458;
  assign n49463 = n45563 & n48222;
  assign n49452 = ~n49457;
  assign n49469 = n45563 & n48132;
  assign n49470 = n49432 & n49458;
  assign n49471 = n45563 & n46901;
  assign n49465 = ~n49482;
  assign n49467 = ~n49432;
  assign n45601 = ~n45563;
  assign n49494 = ~n49519;
  assign n49520 = n49528 & n46802;
  assign n49442 = ~n49529;
  assign n49539 = n49501 & n153;
  assign n49530 = n49556 ^ n49557;
  assign n49538 = ~n49501;
  assign n49558 = ~n49556;
  assign n49571 = ~n49595;
  assign n49375 = ~n48160;
  assign n49386 = n49432 ^ n49433;
  assign n48224 = ~n49463;
  assign n49456 = n45601 & n49464;
  assign n49453 = n49465 & n49466;
  assign n49459 = n49467 & n49468;
  assign n49449 = ~n49469;
  assign n49451 = ~n49470;
  assign n48182 = ~n49471;
  assign n49472 = n49494 & n49495;
  assign n49474 = ~n49520;
  assign n49497 = n154 ^ n49530;
  assign n49533 = n49538 & n4946;
  assign n49478 = ~n49539;
  assign n49547 = n49558 & n49559;
  assign n49540 = n49571 & n49572;
  assign n49408 = n49386 & n1678;
  assign n49409 = ~n49386;
  assign n49377 = n49449 & n49450;
  assign n49438 = n49451 & n49452;
  assign n49431 = ~n49453;
  assign n48250 = ~n49456;
  assign n49427 = ~n49459;
  assign n49440 = n49472 ^ n46802;
  assign n49473 = ~n49472;
  assign n49479 = n49496 ^ n49497;
  assign n49498 = ~n49497;
  assign n49503 = ~n49533;
  assign n49508 = n152 ^ n49540;
  assign n49531 = ~n49547;
  assign n49388 = ~n49408;
  assign n49398 = n49409 & n297;
  assign n49425 = n49430 & n49431;
  assign n49405 = n49431 ^ n49434;
  assign n49429 = n49377 & n49435;
  assign n49428 = ~n49377;
  assign n49426 = ~n49438;
  assign n45547 = n49439 ^ n49440;
  assign n49460 = n49473 & n49474;
  assign n49475 = n49479 & n46784;
  assign n49392 = ~n49479;
  assign n49443 = n49498 & n49499;
  assign n49446 = n49508 ^ n49509;
  assign n49500 = n49531 & n49532;
  assign n49365 = ~n49398;
  assign n49384 = n298 ^ n49405;
  assign n49413 = n45547 & n49424;
  assign n49406 = ~n49425;
  assign n49399 = n49426 & n49427;
  assign n49414 = n49428 & n49400;
  assign n49415 = n45547 & n48122;
  assign n49404 = ~n49429;
  assign n49416 = n45547 & n46802;
  assign n45489 = ~n45547;
  assign n49441 = ~n49460;
  assign n49419 = ~n49475;
  assign n49461 = n49392 & n46813;
  assign n49476 = n49500 ^ n49501;
  assign n49502 = ~n49500;
  assign n48095 = n49383 ^ n49384;
  assign n49342 = n49384 & n49383;
  assign n49378 = n49399 ^ n49400;
  assign n49385 = n49406 & n49407;
  assign n48180 = ~n49413;
  assign n49410 = n45489 & n48204;
  assign n49380 = ~n49414;
  assign n49401 = ~n49415;
  assign n48140 = ~n49416;
  assign n49403 = ~n49399;
  assign n49417 = n49441 & n49442;
  assign n49395 = ~n49461;
  assign n49444 = n153 ^ n49476;
  assign n49485 = n49502 & n49503;
  assign n49333 = ~n48095;
  assign n49347 = n49377 ^ n49378;
  assign n49345 = ~n49342;
  assign n49363 = n49385 ^ n49386;
  assign n49387 = ~n49385;
  assign n49358 = n49401 & n49402;
  assign n49391 = n49403 & n49404;
  assign n48206 = ~n49410;
  assign n49393 = n49417 ^ n46784;
  assign n49418 = ~n49417;
  assign n49351 = n49443 ^ n49444;
  assign n49422 = n49444 & n49443;
  assign n49477 = ~n49485;
  assign n49343 = n297 ^ n49363;
  assign n49356 = n49347 & n296;
  assign n49355 = ~n49347;
  assign n49376 = n49387 & n49388;
  assign n49382 = n49358 & n49389;
  assign n49381 = ~n49358;
  assign n49379 = ~n49391;
  assign n45503 = n49392 ^ n49393;
  assign n49411 = n49418 & n49419;
  assign n49421 = n49351 & n46720;
  assign n49420 = ~n49351;
  assign n49445 = n49477 & n49478;
  assign n49296 = n49342 ^ n49343;
  assign n49344 = ~n49343;
  assign n49349 = n49355 & n1618;
  assign n49315 = ~n49356;
  assign n49368 = n45503 & n49375;
  assign n49364 = ~n49376;
  assign n49357 = n49379 & n49380;
  assign n49369 = n49381 & n49337;
  assign n49370 = n45503 & n48032;
  assign n49362 = ~n49382;
  assign n49371 = n45503 & n46784;
  assign n45465 = ~n45503;
  assign n49394 = ~n49411;
  assign n49412 = n49420 & n46772;
  assign n49374 = ~n49421;
  assign n49423 = n49445 ^ n49446;
  assign n48053 = ~n49296;
  assign n49304 = n49344 & n49345;
  assign n49335 = ~n49349;
  assign n49336 = n49357 ^ n49358;
  assign n49346 = n49364 & n49365;
  assign n48138 = ~n49368;
  assign n49366 = n45465 & n48160;
  assign n49361 = ~n49357;
  assign n49339 = ~n49369;
  assign n49359 = ~n49370;
  assign n48100 = ~n49371;
  assign n49372 = n49394 & n49395;
  assign n49354 = ~n49412;
  assign n49311 = n49422 ^ n49423;
  assign n49274 = n49336 ^ n49337;
  assign n49322 = n49346 ^ n49347;
  assign n49334 = ~n49346;
  assign n49300 = n49359 & n49360;
  assign n49350 = n49361 & n49362;
  assign n48162 = ~n49366;
  assign n49352 = n49372 ^ n46720;
  assign n49373 = ~n49372;
  assign n49397 = n49311 & n46734;
  assign n49396 = ~n49311;
  assign n49305 = n296 ^ n49322;
  assign n49317 = n49274 & n311;
  assign n49316 = ~n49274;
  assign n49328 = n49334 & n49335;
  assign n49341 = n49300 & n49348;
  assign n49340 = ~n49300;
  assign n49338 = ~n49350;
  assign n45411 = n49351 ^ n49352;
  assign n49367 = n49373 & n49374;
  assign n49390 = n49396 & n46699;
  assign n49332 = ~n49397;
  assign n48016 = n49304 ^ n49305;
  assign n49254 = n49305 & n49304;
  assign n49306 = n49316 & n1559;
  assign n49276 = ~n49317;
  assign n49314 = ~n49328;
  assign n49327 = n45411 & n49333;
  assign n49318 = n49338 & n49339;
  assign n49329 = n49340 & n49319;
  assign n49321 = ~n49341;
  assign n45443 = ~n45411;
  assign n49353 = ~n49367;
  assign n49313 = ~n49390;
  assign n49256 = ~n48016;
  assign n49299 = ~n49306;
  assign n49297 = n49314 & n49315;
  assign n49301 = n49318 ^ n49319;
  assign n49323 = n45443 & n48095;
  assign n48120 = ~n49327;
  assign n49320 = ~n49318;
  assign n49303 = ~n49329;
  assign n49324 = n45443 & n48012;
  assign n49325 = n45443 & n46720;
  assign n49330 = n49353 & n49354;
  assign n49273 = n311 ^ n49297;
  assign n49258 = n49300 ^ n49301;
  assign n49298 = ~n49297;
  assign n49309 = n49320 & n49321;
  assign n48098 = ~n49323;
  assign n49307 = ~n49324;
  assign n48058 = ~n49325;
  assign n49310 = n49330 ^ n46734;
  assign n49331 = ~n49330;
  assign n49255 = n49273 ^ n49274;
  assign n49278 = n49258 & n310;
  assign n49277 = ~n49258;
  assign n49289 = n49298 & n49299;
  assign n49261 = n49307 & n49308;
  assign n49302 = ~n49309;
  assign n45343 = n49310 ^ n49311;
  assign n49326 = n49331 & n49332;
  assign n47970 = n49254 ^ n49255;
  assign n49211 = n49255 & n49254;
  assign n49265 = n49277 & n1507;
  assign n49232 = ~n49278;
  assign n49275 = ~n49289;
  assign n49288 = n45343 & n49296;
  assign n49279 = n49302 & n49303;
  assign n49292 = n49261 & n49280;
  assign n49290 = ~n49261;
  assign n45391 = ~n45343;
  assign n49312 = ~n49326;
  assign n49208 = ~n47970;
  assign n49214 = ~n49211;
  assign n49260 = ~n49265;
  assign n49257 = n49275 & n49276;
  assign n49262 = n49279 ^ n49280;
  assign n48080 = ~n49288;
  assign n49283 = n45391 & n48053;
  assign n49281 = ~n49279;
  assign n49284 = n49290 & n49291;
  assign n49285 = n45391 & n47958;
  assign n49282 = ~n49292;
  assign n49286 = n45391 & n46734;
  assign n49293 = n49312 & n49313;
  assign n49230 = n49257 ^ n49258;
  assign n49216 = n49261 ^ n49262;
  assign n49259 = ~n49257;
  assign n49268 = n49281 & n49282;
  assign n48056 = ~n49283;
  assign n49264 = ~n49284;
  assign n49266 = ~n49285;
  assign n48020 = ~n49286;
  assign n49270 = n49293 ^ n46660;
  assign n49294 = ~n49293;
  assign n49212 = n310 ^ n49230;
  assign n49233 = n49216 & n1450;
  assign n49234 = ~n49216;
  assign n49244 = n49259 & n49260;
  assign n49217 = n49266 & n49267;
  assign n49263 = ~n49268;
  assign n45272 = n49269 ^ n49270;
  assign n49287 = n49294 & n49295;
  assign n47927 = n49211 ^ n49212;
  assign n49213 = ~n49212;
  assign n49210 = ~n49233;
  assign n49224 = n49234 & n309;
  assign n49231 = ~n49244;
  assign n49245 = n45272 & n49256;
  assign n49235 = n49263 & n49264;
  assign n49248 = n45272 & n47949;
  assign n49249 = n49217 & n49236;
  assign n49250 = n45272 & n46660;
  assign n49246 = ~n49217;
  assign n45328 = ~n45272;
  assign n49271 = ~n49287;
  assign n49168 = ~n47927;
  assign n49166 = n49213 & n49214;
  assign n49189 = ~n49224;
  assign n49215 = n49231 & n49232;
  assign n49218 = n49235 ^ n49236;
  assign n48018 = ~n49245;
  assign n49241 = n45328 & n48016;
  assign n49238 = ~n49235;
  assign n49242 = n49246 & n49247;
  assign n49239 = ~n49248;
  assign n49237 = ~n49249;
  assign n47969 = ~n49250;
  assign n49251 = n49271 & n49272;
  assign n49187 = n49215 ^ n49216;
  assign n49170 = n49217 ^ n49218;
  assign n49209 = ~n49215;
  assign n49225 = n49237 & n49238;
  assign n49173 = n49239 & n49240;
  assign n48040 = ~n49241;
  assign n49220 = ~n49242;
  assign n49226 = n49251 ^ n46650;
  assign n49252 = ~n49251;
  assign n49167 = n309 ^ n49187;
  assign n49190 = n49170 & n1423;
  assign n49191 = ~n49170;
  assign n49201 = n49209 & n49210;
  assign n49222 = n49173 & n49223;
  assign n49219 = ~n49225;
  assign n49221 = ~n49173;
  assign n45157 = n49226 ^ n49227;
  assign n49243 = n49252 & n49253;
  assign n47888 = n49166 ^ n49167;
  assign n49127 = n49167 & n49166;
  assign n49171 = ~n49190;
  assign n49181 = n49191 & n308;
  assign n49188 = ~n49201;
  assign n49200 = n45157 & n49208;
  assign n49192 = n49219 & n49220;
  assign n49202 = n49221 & n49193;
  assign n49203 = n45157 & n47878;
  assign n49197 = ~n49222;
  assign n49204 = n45157 & n46650;
  assign n45258 = ~n45157;
  assign n49228 = ~n49243;
  assign n49101 = ~n47888;
  assign n49149 = ~n49181;
  assign n49169 = n49188 & n49189;
  assign n49174 = n49192 ^ n49193;
  assign n47973 = ~n49200;
  assign n49198 = n45258 & n47970;
  assign n49196 = ~n49192;
  assign n49176 = ~n49202;
  assign n49194 = ~n49203;
  assign n47936 = ~n49204;
  assign n49205 = n49228 & n49229;
  assign n49147 = n49169 ^ n49170;
  assign n49130 = n49173 ^ n49174;
  assign n49172 = ~n49169;
  assign n49153 = n49194 & n49195;
  assign n49182 = n49196 & n49197;
  assign n47996 = ~n49198;
  assign n49184 = n49205 ^ n46565;
  assign n49206 = ~n49205;
  assign n49128 = n308 ^ n49147;
  assign n49151 = n49130 & n307;
  assign n49150 = ~n49130;
  assign n49161 = n49171 & n49172;
  assign n49179 = n49153 & n49134;
  assign n49177 = ~n49153;
  assign n49175 = ~n49182;
  assign n45113 = n49183 ^ n49184;
  assign n49199 = n49206 & n49207;
  assign n47844 = n49127 ^ n49128;
  assign n49084 = n49128 & n49127;
  assign n49141 = n49150 & n1356;
  assign n49110 = ~n49151;
  assign n49148 = ~n49161;
  assign n49162 = n45113 & n49168;
  assign n49152 = n49175 & n49176;
  assign n49163 = n49177 & n49178;
  assign n49155 = ~n49179;
  assign n45174 = ~n45113;
  assign n49185 = ~n49199;
  assign n49100 = ~n47844;
  assign n49132 = ~n49141;
  assign n49129 = n49148 & n49149;
  assign n49133 = n49152 ^ n49153;
  assign n47956 = ~n49162;
  assign n49157 = n45174 & n47927;
  assign n49154 = ~n49152;
  assign n49136 = ~n49163;
  assign n49158 = n45174 & n47836;
  assign n49159 = n45174 & n46606;
  assign n49180 = n49185 & n49186;
  assign n49108 = n49129 ^ n49130;
  assign n49089 = n49133 ^ n49134;
  assign n49131 = ~n49129;
  assign n49144 = n49154 & n49155;
  assign n47930 = ~n49157;
  assign n49142 = ~n49158;
  assign n47896 = ~n49159;
  assign n49165 = n49180 & n46553;
  assign n49164 = ~n49180;
  assign n49085 = n307 ^ n49108;
  assign n49111 = n49089 & n1286;
  assign n49112 = ~n49089;
  assign n49124 = n49131 & n49132;
  assign n49093 = n49142 & n49143;
  assign n49135 = ~n49144;
  assign n49160 = n49164 & n46512;
  assign n49146 = ~n49165;
  assign n47827 = n49084 ^ n49085;
  assign n49086 = ~n49085;
  assign n49091 = ~n49111;
  assign n49105 = n49112 & n306;
  assign n49109 = ~n49124;
  assign n49113 = n49135 & n49136;
  assign n49126 = n49093 & n49137;
  assign n49125 = ~n49093;
  assign n49145 = n49146 & n49156;
  assign n49139 = ~n49160;
  assign n49039 = ~n47827;
  assign n49043 = n49086 & n49084;
  assign n49065 = ~n49105;
  assign n49088 = n49109 & n49110;
  assign n49094 = n49113 ^ n49114;
  assign n49115 = ~n49113;
  assign n49121 = n49125 & n49114;
  assign n49116 = ~n49126;
  assign n49138 = ~n49145;
  assign n49140 = n49139 & n49146;
  assign n49046 = ~n49043;
  assign n49063 = n49088 ^ n49089;
  assign n49048 = n49093 ^ n49094;
  assign n49090 = ~n49088;
  assign n49106 = n49115 & n49116;
  assign n49096 = ~n49121;
  assign n49118 = n49138 & n49139;
  assign n49123 = ~n49140;
  assign n49044 = n306 ^ n49063;
  assign n49067 = n49048 & n305;
  assign n49066 = ~n49048;
  assign n49080 = n49090 & n49091;
  assign n49095 = ~n49106;
  assign n44891 = n49117 ^ n49118;
  assign n45040 = n49122 ^ n49123;
  assign n49119 = ~n49118;
  assign n47760 = n49043 ^ n49044;
  assign n49045 = ~n49044;
  assign n49060 = n49066 & n1201;
  assign n49031 = ~n49067;
  assign n49064 = ~n49080;
  assign n49068 = n49095 & n49096;
  assign n49087 = n44891 & n49100;
  assign n49097 = n44891 & n47796;
  assign n49102 = n45040 & n47888;
  assign n49103 = n45040 & n47792;
  assign n49104 = n45040 & n46553;
  assign n45000 = ~n44891;
  assign n49107 = n49119 & n49120;
  assign n45056 = ~n45040;
  assign n48994 = ~n47760;
  assign n49008 = n49045 & n49046;
  assign n49050 = ~n49060;
  assign n49047 = n49064 & n49065;
  assign n49052 = n49068 ^ n49069;
  assign n49071 = n49068 & n49076;
  assign n49070 = ~n49068;
  assign n49079 = n45000 & n47844;
  assign n47872 = ~n49087;
  assign n49077 = ~n49097;
  assign n49083 = n45000 & n46498;
  assign n49092 = n45056 & n49101;
  assign n47890 = ~n49102;
  assign n49081 = ~n49103;
  assign n47857 = ~n49104;
  assign n49098 = ~n49107;
  assign n49032 = n49047 ^ n49048;
  assign n49049 = ~n49047;
  assign n49061 = n49070 & n49069;
  assign n49058 = ~n49071;
  assign n48986 = n49077 & n49078;
  assign n47847 = ~n49079;
  assign n49051 = n49081 & n49082;
  assign n47817 = ~n49083;
  assign n47914 = ~n49092;
  assign n49072 = n49098 & n49099;
  assign n49009 = n305 ^ n49032;
  assign n49042 = n49049 & n49050;
  assign n49011 = n49051 ^ n49052;
  assign n49041 = ~n49061;
  assign n49054 = n49072 ^ n49073;
  assign n49059 = ~n49051;
  assign n49074 = ~n49072;
  assign n48956 = n49008 ^ n49009;
  assign n48974 = n49009 & n49008;
  assign n49034 = n49011 & n304;
  assign n49030 = ~n49042;
  assign n49029 = ~n49011;
  assign n44851 = n46435 ^ n49054;
  assign n49053 = n49058 & n49059;
  assign n49055 = n49054 & n46357;
  assign n49062 = n49074 & n49075;
  assign n47724 = ~n48956;
  assign n49025 = n49029 & n1168;
  assign n49010 = n49030 & n49031;
  assign n48997 = ~n49034;
  assign n49033 = n44851 & n49039;
  assign n49035 = n44851 & n47689;
  assign n44946 = ~n44851;
  assign n49040 = ~n49053;
  assign n47773 = ~n49055;
  assign n49056 = ~n49062;
  assign n48993 = n49010 ^ n49011;
  assign n49012 = ~n49010;
  assign n49013 = ~n49025;
  assign n49024 = n44946 & n47827;
  assign n47803 = ~n49033;
  assign n49019 = ~n49035;
  assign n49026 = n49040 & n49041;
  assign n49036 = n49056 & n49057;
  assign n48975 = n304 ^ n48993;
  assign n49007 = n49012 & n49013;
  assign n48971 = n49019 & n49020;
  assign n47829 = ~n49024;
  assign n49023 = n49026 & n49027;
  assign n49021 = ~n49026;
  assign n49016 = n49036 ^ n46321;
  assign n49037 = ~n49036;
  assign n48924 = n48974 ^ n48975;
  assign n48936 = n48975 & n48974;
  assign n48996 = ~n49007;
  assign n49006 = n48971 & n48949;
  assign n49003 = ~n48971;
  assign n44768 = n49015 ^ n49016;
  assign n49014 = n49021 & n49022;
  assign n49005 = ~n49023;
  assign n49028 = n49037 & n49038;
  assign n47678 = ~n48924;
  assign n48976 = n48996 & n48997;
  assign n48995 = n44768 & n47760;
  assign n48998 = n49003 & n49004;
  assign n48973 = ~n49006;
  assign n49002 = n49005 & n48986;
  assign n44855 = ~n44768;
  assign n48989 = ~n49014;
  assign n49017 = ~n49028;
  assign n48954 = n319 ^ n48976;
  assign n48978 = n48976 & n1118;
  assign n48977 = ~n48976;
  assign n48987 = n44855 & n48994;
  assign n47785 = ~n48995;
  assign n48951 = ~n48998;
  assign n48990 = n44855 & n47649;
  assign n48991 = n44855 & n46321;
  assign n48988 = ~n49002;
  assign n48985 = n48989 & n49005;
  assign n48999 = n49017 & n49018;
  assign n48969 = n48977 & n319;
  assign n48966 = ~n48978;
  assign n48955 = n48985 ^ n48986;
  assign n47763 = ~n48987;
  assign n48970 = n48988 & n48989;
  assign n48979 = ~n48990;
  assign n47722 = ~n48991;
  assign n48981 = n48999 ^ n46306;
  assign n49000 = ~n48999;
  assign n48937 = n48954 ^ n48955;
  assign n48958 = n48966 & n48955;
  assign n48944 = ~n48969;
  assign n48948 = n48970 ^ n48971;
  assign n48933 = n48979 & n48980;
  assign n44685 = n48981 ^ n48982;
  assign n48972 = ~n48970;
  assign n48992 = n49000 & n49001;
  assign n47634 = n48936 ^ n48937;
  assign n48874 = n48937 & n48936;
  assign n48919 = n48948 ^ n48949;
  assign n48943 = ~n48958;
  assign n48957 = n44685 & n47724;
  assign n48960 = n48933 & n48968;
  assign n48961 = n44685 & n47673;
  assign n48962 = n44685 & n46306;
  assign n48967 = n48972 & n48973;
  assign n48959 = ~n48933;
  assign n44786 = ~n44685;
  assign n48983 = ~n48992;
  assign n48888 = ~n47634;
  assign n48931 = n48919 & n1025;
  assign n48877 = ~n48874;
  assign n48938 = n48943 & n48944;
  assign n48930 = ~n48919;
  assign n48947 = n44786 & n48956;
  assign n47726 = ~n48957;
  assign n48952 = n48959 & n48910;
  assign n48935 = ~n48960;
  assign n48945 = ~n48961;
  assign n47691 = ~n48962;
  assign n48950 = ~n48967;
  assign n48963 = n48983 & n48984;
  assign n48925 = n48930 & n318;
  assign n48916 = ~n48931;
  assign n48917 = ~n48938;
  assign n48867 = n48945 & n48946;
  assign n47749 = ~n48947;
  assign n48932 = n48950 & n48951;
  assign n48912 = ~n48952;
  assign n48940 = n48963 ^ n46161;
  assign n48964 = ~n48963;
  assign n48907 = n48916 & n48917;
  assign n48898 = n48917 ^ n48919;
  assign n48900 = ~n48925;
  assign n48909 = n48932 ^ n48933;
  assign n48929 = n48867 & n48895;
  assign n48927 = ~n48867;
  assign n44689 = n48939 ^ n48940;
  assign n48934 = ~n48932;
  assign n48953 = n48964 & n48965;
  assign n48875 = n318 ^ n48898;
  assign n48899 = ~n48907;
  assign n48879 = n48909 ^ n48910;
  assign n48918 = n44689 & n48924;
  assign n48920 = n48927 & n48928;
  assign n48897 = ~n48929;
  assign n48926 = n48934 & n48935;
  assign n44668 = ~n44689;
  assign n48941 = ~n48953;
  assign n47584 = n48874 ^ n48875;
  assign n48876 = ~n48875;
  assign n48878 = n48899 & n48900;
  assign n48893 = n48879 & n317;
  assign n48892 = ~n48879;
  assign n48908 = n44668 & n47678;
  assign n47707 = ~n48918;
  assign n48872 = ~n48920;
  assign n48913 = n44668 & n47623;
  assign n48914 = n44668 & n46227;
  assign n48911 = ~n48926;
  assign n48921 = n48941 & n48942;
  assign n48839 = ~n47584;
  assign n48835 = n48876 & n48877;
  assign n48858 = n48878 ^ n48879;
  assign n48869 = ~n48878;
  assign n48889 = n48892 & n970;
  assign n48851 = ~n48893;
  assign n47681 = ~n48908;
  assign n48894 = n48911 & n48912;
  assign n48901 = ~n48913;
  assign n47647 = ~n48914;
  assign n48904 = n48921 ^ n46082;
  assign n48922 = ~n48921;
  assign n48836 = n317 ^ n48858;
  assign n48870 = ~n48889;
  assign n48868 = n48894 ^ n48895;
  assign n48830 = n48901 & n48902;
  assign n44513 = n48903 ^ n48904;
  assign n48896 = ~n48894;
  assign n48915 = n48922 & n48923;
  assign n47531 = n48835 ^ n48836;
  assign n48837 = ~n48836;
  assign n48827 = n48867 ^ n48868;
  assign n48861 = n48869 & n48870;
  assign n48880 = n44513 & n48888;
  assign n48883 = n48830 & n48855;
  assign n48884 = n44513 & n47559;
  assign n48885 = n44513 & n46149;
  assign n48890 = n48896 & n48897;
  assign n48881 = ~n48830;
  assign n44602 = ~n44513;
  assign n48905 = ~n48915;
  assign n48791 = n48837 & n48835;
  assign n48852 = n48827 & n901;
  assign n48850 = ~n48861;
  assign n48853 = ~n48827;
  assign n48866 = n44602 & n47634;
  assign n47636 = ~n48880;
  assign n48873 = n48881 & n48882;
  assign n48857 = ~n48883;
  assign n48862 = ~n48884;
  assign n47582 = ~n48885;
  assign n48871 = ~n48890;
  assign n48886 = n48905 & n48906;
  assign n48826 = n48850 & n48851;
  assign n48828 = ~n48852;
  assign n48843 = n48853 & n316;
  assign n48797 = n48862 & n48863;
  assign n47663 = ~n48866;
  assign n48854 = n48871 & n48872;
  assign n48833 = ~n48873;
  assign n48860 = n48886 ^ n46011;
  assign n48887 = n48886 & n48891;
  assign n48809 = n48826 ^ n48827;
  assign n48829 = ~n48826;
  assign n48811 = ~n48843;
  assign n48831 = n48854 ^ n48855;
  assign n48847 = n48797 & n48815;
  assign n48845 = ~n48797;
  assign n44445 = n48859 ^ n48860;
  assign n48856 = ~n48854;
  assign n48864 = ~n48887;
  assign n48792 = n316 ^ n48809;
  assign n48820 = n48828 & n48829;
  assign n48794 = n48830 ^ n48831;
  assign n48838 = n44445 & n47584;
  assign n48840 = n48845 & n48846;
  assign n48817 = ~n48847;
  assign n48841 = n44445 & n47454;
  assign n48842 = n44445 & n46011;
  assign n48844 = n48856 & n48857;
  assign n44528 = ~n44445;
  assign n48848 = n48864 & n48865;
  assign n48779 = n48791 ^ n48792;
  assign n48767 = n48792 & n48791;
  assign n48812 = n48794 & n840;
  assign n48810 = ~n48820;
  assign n48813 = ~n48794;
  assign n47586 = ~n48838;
  assign n48825 = n44528 & n48839;
  assign n48800 = ~n48840;
  assign n48821 = ~n48841;
  assign n47543 = ~n48842;
  assign n48832 = ~n48844;
  assign n47516 = n48848 ^ n48849;
  assign n45539 = n46551 ^ n48779;
  assign n48780 = n48779 & n46549;
  assign n48723 = n48779 & n46551;
  assign n48793 = n48810 & n48811;
  assign n48796 = ~n48812;
  assign n48804 = n48813 & n315;
  assign n48773 = n48821 & n48822;
  assign n47614 = ~n48825;
  assign n48814 = n48832 & n48833;
  assign n48823 = n47516 & n47468;
  assign n48824 = n47516 & n48834;
  assign n44492 = ~n47516;
  assign n48766 = n45539 & n47590;
  assign n45535 = ~n45539;
  assign n47616 = ~n48780;
  assign n48781 = n48793 ^ n48794;
  assign n48795 = ~n48793;
  assign n48783 = ~n48804;
  assign n48798 = n48814 ^ n48815;
  assign n48808 = n48773 & n48787;
  assign n48806 = ~n48773;
  assign n48816 = ~n48814;
  assign n48818 = ~n48823;
  assign n47492 = ~n48824;
  assign n45536 = n423 ^ n45535;
  assign n48762 = ~n48766;
  assign n48768 = n315 ^ n48781;
  assign n48790 = n48795 & n48796;
  assign n48770 = n48797 ^ n48798;
  assign n48803 = n48806 & n48807;
  assign n48789 = ~n48808;
  assign n48805 = n48816 & n48817;
  assign n48801 = n48818 & n48819;
  assign n48748 = n48762 & n48763;
  assign n48764 = n48767 ^ n48768;
  assign n48738 = n48768 & n48767;
  assign n48784 = n48770 & n792;
  assign n48782 = ~n48790;
  assign n48785 = ~n48770;
  assign n48747 = n48801 ^ n48802;
  assign n48776 = ~n48803;
  assign n48799 = ~n48805;
  assign n48733 = n48748 ^ n48749;
  assign n48750 = ~n48748;
  assign n48754 = n48764 & n46432;
  assign n48755 = ~n48764;
  assign n48741 = ~n48738;
  assign n48769 = n48782 & n48783;
  assign n48772 = ~n48784;
  assign n48777 = n48785 & n314;
  assign n48786 = n48799 & n48800;
  assign n47180 = n455 ^ n48733;
  assign n48619 = n48733 & n455;
  assign n48666 = n48750 & n48751;
  assign n48727 = ~n48754;
  assign n48752 = n48755 & n46439;
  assign n48756 = n48769 ^ n48770;
  assign n48771 = ~n48769;
  assign n48758 = ~n48777;
  assign n48774 = n48786 ^ n48787;
  assign n48788 = ~n48786;
  assign n48440 = ~n47180;
  assign n48737 = ~n48752;
  assign n48739 = n314 ^ n48756;
  assign n48765 = n48771 & n48772;
  assign n48743 = n48773 ^ n48774;
  assign n48778 = n48788 & n48789;
  assign n48734 = n48737 & n48723;
  assign n48735 = n48737 & n48727;
  assign n48704 = n48738 ^ n48739;
  assign n48740 = ~n48739;
  assign n48759 = n48743 & n746;
  assign n48757 = ~n48765;
  assign n48760 = ~n48743;
  assign n48775 = ~n48778;
  assign n48728 = n48704 & n46335;
  assign n48726 = ~n48734;
  assign n48724 = ~n48735;
  assign n48729 = ~n48704;
  assign n48718 = n48740 & n48741;
  assign n48742 = n48757 & n48758;
  assign n48745 = ~n48759;
  assign n48753 = n48760 & n313;
  assign n48761 = n48775 & n48776;
  assign n45509 = n48723 ^ n48724;
  assign n48715 = n48726 & n48727;
  assign n48716 = ~n48728;
  assign n48725 = n48729 & n46371;
  assign n48722 = ~n48718;
  assign n48730 = n48742 ^ n48743;
  assign n48744 = ~n48742;
  assign n48732 = ~n48753;
  assign n48746 = n312 ^ n48761;
  assign n48705 = n48715 ^ n46371;
  assign n45520 = ~n45509;
  assign n48717 = ~n48715;
  assign n48707 = ~n48725;
  assign n48719 = n313 ^ n48730;
  assign n48736 = n48744 & n48745;
  assign n48721 = n48746 ^ n48747;
  assign n45367 = n48704 ^ n48705;
  assign n48712 = n45520 & n47494;
  assign n48713 = n45520 & n46439;
  assign n48714 = n48716 & n48717;
  assign n48681 = n48718 ^ n48719;
  assign n48710 = n48719 & n48722;
  assign n48731 = ~n48736;
  assign n48692 = n45367 & n47435;
  assign n48693 = n45367 & n46335;
  assign n45365 = ~n45367;
  assign n48708 = n48681 & n46303;
  assign n48701 = ~n48712;
  assign n47518 = ~n48713;
  assign n48706 = ~n48714;
  assign n48709 = ~n48681;
  assign n48720 = n48731 & n48732;
  assign n48684 = ~n48692;
  assign n47484 = ~n48693;
  assign n48694 = n48701 & n48702;
  assign n48696 = n48706 & n48707;
  assign n48698 = ~n48708;
  assign n48703 = n48709 & n46262;
  assign n48711 = n48720 ^ n48721;
  assign n48634 = n48684 & n48685;
  assign n48689 = n48694 & n48695;
  assign n48680 = n48696 ^ n46303;
  assign n48687 = ~n48694;
  assign n48697 = ~n48696;
  assign n48683 = ~n48703;
  assign n48660 = n48710 ^ n48711;
  assign n48677 = n48634 & n48654;
  assign n48675 = ~n48634;
  assign n45280 = n48680 ^ n48681;
  assign n48686 = n48687 & n48688;
  assign n48679 = ~n48689;
  assign n48690 = n48697 & n48698;
  assign n48700 = n48660 & n46224;
  assign n48699 = ~n48660;
  assign n48669 = n48675 & n48676;
  assign n48657 = ~n48677;
  assign n45282 = ~n45280;
  assign n48678 = n48679 & n48666;
  assign n48671 = ~n48686;
  assign n48682 = ~n48690;
  assign n48691 = n48699 & n46182;
  assign n48674 = ~n48700;
  assign n48642 = ~n48669;
  assign n48663 = n45282 & n47383;
  assign n48664 = n45282 & n46303;
  assign n48670 = ~n48678;
  assign n48665 = n48671 & n48679;
  assign n48672 = n48682 & n48683;
  assign n48662 = ~n48691;
  assign n48655 = ~n48663;
  assign n47432 = ~n48664;
  assign n48658 = n48665 ^ n48666;
  assign n48667 = n48670 & n48671;
  assign n48659 = n48672 ^ n46224;
  assign n48673 = ~n48672;
  assign n48604 = n48655 & n48656;
  assign n48652 = n48658 & n454;
  assign n45179 = n48659 ^ n48660;
  assign n48651 = ~n48658;
  assign n48653 = ~n48667;
  assign n48668 = n48673 & n48674;
  assign n48645 = n48604 & n48624;
  assign n48643 = ~n48604;
  assign n48649 = n48651 & n18650;
  assign n48621 = ~n48652;
  assign n45188 = ~n45179;
  assign n48635 = n48653 ^ n48654;
  assign n48650 = n48657 & n48653;
  assign n48661 = ~n48668;
  assign n48597 = n48634 ^ n48635;
  assign n48636 = n48643 & n48644;
  assign n48638 = n45188 & n47306;
  assign n48627 = ~n48645;
  assign n48639 = n45188 & n46224;
  assign n48637 = ~n48649;
  assign n48641 = ~n48650;
  assign n48646 = n48661 & n48662;
  assign n48617 = n48597 & n453;
  assign n48616 = ~n48597;
  assign n48607 = ~n48636;
  assign n48633 = n48637 & n48619;
  assign n48618 = n48637 & n48621;
  assign n48625 = ~n48638;
  assign n47354 = ~n48639;
  assign n48623 = n48641 & n48642;
  assign n48630 = n48646 ^ n46091;
  assign n48647 = ~n48646;
  assign n48613 = n48616 & n18542;
  assign n48582 = ~n48617;
  assign n47122 = n48618 ^ n48619;
  assign n48605 = n48623 ^ n48624;
  assign n48569 = n48625 & n48626;
  assign n45088 = n48629 ^ n48630;
  assign n48620 = ~n48633;
  assign n48628 = ~n48623;
  assign n48640 = n48647 & n48648;
  assign n48561 = n48604 ^ n48605;
  assign n48599 = ~n48613;
  assign n48610 = n48569 & n48588;
  assign n47153 = ~n47122;
  assign n48608 = ~n48569;
  assign n48614 = n48620 & n48621;
  assign n45090 = ~n45088;
  assign n48622 = n48627 & n48628;
  assign n48631 = ~n48640;
  assign n48585 = n48561 & n18500;
  assign n48586 = ~n48561;
  assign n48600 = n48608 & n48609;
  assign n48592 = ~n48610;
  assign n48601 = n45090 & n47248;
  assign n48602 = n45090 & n46111;
  assign n48596 = ~n48614;
  assign n48606 = ~n48622;
  assign n48615 = n48631 & n48632;
  assign n48565 = ~n48585;
  assign n48580 = n48586 & n452;
  assign n48575 = n48596 ^ n48597;
  assign n48595 = n48599 & n48596;
  assign n48572 = ~n48600;
  assign n48589 = ~n48601;
  assign n47308 = ~n48602;
  assign n48587 = n48606 & n48607;
  assign n48612 = n48615 & n46037;
  assign n48611 = ~n48615;
  assign n48557 = n453 ^ n48575;
  assign n48545 = ~n48580;
  assign n48570 = n48587 ^ n48588;
  assign n48533 = n48589 & n48590;
  assign n48581 = ~n48595;
  assign n48591 = ~n48587;
  assign n48603 = n48611 & n45997;
  assign n48594 = ~n48612;
  assign n47096 = n48557 ^ n47122;
  assign n48530 = n48569 ^ n48570;
  assign n48559 = ~n48557;
  assign n48574 = n48533 & n48577;
  assign n48576 = n48581 & n48582;
  assign n48573 = ~n48533;
  assign n48583 = n48591 & n48592;
  assign n48593 = n48594 & n48598;
  assign n48579 = ~n48603;
  assign n48364 = ~n47096;
  assign n48550 = n48530 & n18450;
  assign n48519 = n48559 & n47153;
  assign n48551 = ~n48530;
  assign n48566 = n48573 & n48553;
  assign n48555 = ~n48574;
  assign n48560 = ~n48576;
  assign n48571 = ~n48583;
  assign n48578 = ~n48593;
  assign n48584 = n48579 & n48594;
  assign n48531 = ~n48550;
  assign n48546 = n48551 & n451;
  assign n48522 = ~n48519;
  assign n48539 = n48560 ^ n48561;
  assign n48558 = n48565 & n48560;
  assign n48536 = ~n48566;
  assign n48552 = n48571 & n48572;
  assign n48562 = n48578 & n48579;
  assign n48567 = ~n48584;
  assign n48520 = n452 ^ n48539;
  assign n48506 = ~n48546;
  assign n48534 = n48552 ^ n48553;
  assign n48544 = ~n48558;
  assign n48540 = n48562 ^ n45936;
  assign n48554 = ~n48552;
  assign n44966 = n48567 ^ n48568;
  assign n48563 = ~n48562;
  assign n47060 = n48519 ^ n48520;
  assign n48521 = ~n48520;
  assign n48489 = n48533 ^ n48534;
  assign n44862 = n48540 ^ n48541;
  assign n48529 = n48544 & n48545;
  assign n48547 = n48554 & n48555;
  assign n48548 = n44966 & n47232;
  assign n48549 = n44966 & n46037;
  assign n48556 = n48563 & n48564;
  assign n44980 = ~n44966;
  assign n48332 = ~n47060;
  assign n48484 = n48521 & n48522;
  assign n48512 = n48489 & n450;
  assign n48504 = n48529 ^ n48530;
  assign n48511 = ~n48489;
  assign n48524 = n44862 & n47202;
  assign n48525 = n44862 & n45963;
  assign n44902 = ~n44862;
  assign n48532 = ~n48529;
  assign n48535 = ~n48547;
  assign n48537 = ~n48548;
  assign n47265 = ~n48549;
  assign n48542 = ~n48556;
  assign n48485 = n451 ^ n48504;
  assign n48487 = ~n48484;
  assign n48507 = n48511 & n18410;
  assign n48468 = ~n48512;
  assign n48508 = ~n48524;
  assign n47222 = ~n48525;
  assign n48523 = n48531 & n48532;
  assign n48513 = n48535 & n48536;
  assign n48494 = n48537 & n48538;
  assign n48526 = n48542 & n48543;
  assign n47022 = n48484 ^ n48485;
  assign n48486 = ~n48485;
  assign n48490 = ~n48507;
  assign n48434 = n48508 & n48509;
  assign n48495 = n48513 ^ n48514;
  assign n48505 = ~n48523;
  assign n48517 = n48494 & n48514;
  assign n48498 = n48526 ^ n45909;
  assign n48501 = ~n48513;
  assign n48515 = ~n48494;
  assign n48527 = ~n48526;
  assign n48285 = ~n47022;
  assign n48446 = n48486 & n48487;
  assign n48451 = n48494 ^ n48495;
  assign n48493 = n48434 & n48496;
  assign n48492 = ~n48434;
  assign n44822 = n48498 ^ n48499;
  assign n48488 = n48505 & n48506;
  assign n48510 = n48515 & n48516;
  assign n48500 = ~n48517;
  assign n48518 = n48527 & n48528;
  assign n48449 = ~n48446;
  assign n48472 = n48451 & n18389;
  assign n48466 = n48488 ^ n48489;
  assign n48473 = ~n48451;
  assign n48476 = n48492 & n48463;
  assign n48458 = ~n48493;
  assign n48477 = n44822 & n47150;
  assign n48478 = n44822 & n45909;
  assign n44778 = ~n44822;
  assign n48491 = ~n48488;
  assign n48497 = n48500 & n48501;
  assign n48480 = ~n48510;
  assign n48502 = ~n48518;
  assign n48447 = n450 ^ n48466;
  assign n48453 = ~n48472;
  assign n48469 = n48473 & n449;
  assign n48437 = ~n48476;
  assign n48470 = ~n48477;
  assign n47183 = ~n48478;
  assign n48475 = n48490 & n48491;
  assign n48479 = ~n48497;
  assign n48481 = n48502 & n48503;
  assign n46993 = n48446 ^ n48447;
  assign n48448 = ~n48447;
  assign n48427 = ~n48469;
  assign n48395 = n48470 & n48471;
  assign n48467 = ~n48475;
  assign n48462 = n48479 & n48480;
  assign n48460 = n48481 ^ n45853;
  assign n48482 = ~n48481;
  assign n48244 = ~n46993;
  assign n48405 = n48448 & n48449;
  assign n48456 = n48395 & n48419;
  assign n48454 = ~n48395;
  assign n44697 = n48460 ^ n48461;
  assign n48435 = n48462 ^ n48463;
  assign n48450 = n48467 & n48468;
  assign n48459 = ~n48462;
  assign n48474 = n48482 & n48483;
  assign n48408 = ~n48405;
  assign n48410 = n48434 ^ n48435;
  assign n48428 = n48450 ^ n48451;
  assign n48438 = n48454 & n48455;
  assign n48421 = ~n48456;
  assign n48439 = n44697 & n47110;
  assign n48441 = n44697 & n47180;
  assign n48442 = n44697 & n45853;
  assign n44747 = ~n44697;
  assign n48452 = ~n48450;
  assign n48457 = n48458 & n48459;
  assign n48464 = ~n48474;
  assign n48417 = n48410 & n448;
  assign n48406 = n449 ^ n48428;
  assign n48416 = ~n48410;
  assign n48400 = ~n48438;
  assign n48429 = ~n48439;
  assign n48431 = n44747 & n48440;
  assign n47185 = ~n48441;
  assign n47148 = ~n48442;
  assign n48433 = n48452 & n48453;
  assign n48436 = ~n48457;
  assign n48443 = n48464 & n48465;
  assign n48200 = n48405 ^ n48406;
  assign n48414 = n48416 & n18335;
  assign n48407 = ~n48406;
  assign n48379 = ~n48417;
  assign n48359 = n48429 & n48430;
  assign n47206 = ~n48431;
  assign n48426 = ~n48433;
  assign n48418 = n48436 & n48437;
  assign n48423 = n48443 ^ n45788;
  assign n48444 = ~n48443;
  assign n46953 = ~n48200;
  assign n48370 = n48407 & n48408;
  assign n48412 = n48359 & n48413;
  assign n48397 = ~n48414;
  assign n48396 = n48418 ^ n48419;
  assign n48411 = ~n48359;
  assign n44611 = n48422 ^ n48423;
  assign n48409 = n48426 & n48427;
  assign n48420 = ~n48418;
  assign n48432 = n48444 & n48445;
  assign n48352 = n48395 ^ n48396;
  assign n48390 = n48409 ^ n48410;
  assign n48401 = n48411 & n48381;
  assign n48383 = ~n48412;
  assign n44651 = ~n44611;
  assign n48398 = ~n48409;
  assign n48415 = n48420 & n48421;
  assign n48424 = ~n48432;
  assign n48371 = n448 ^ n48390;
  assign n48376 = n48352 & n18294;
  assign n48377 = ~n48352;
  assign n48391 = n48397 & n48398;
  assign n48362 = ~n48401;
  assign n48392 = n44651 & n47075;
  assign n48393 = n44651 & n45788;
  assign n48399 = ~n48415;
  assign n48402 = n48424 & n48425;
  assign n48157 = n48370 ^ n48371;
  assign n48309 = n48371 & n48370;
  assign n48358 = ~n48376;
  assign n48373 = n48377 & n463;
  assign n48378 = ~n48391;
  assign n48384 = ~n48392;
  assign n47090 = ~n48393;
  assign n48380 = n48399 & n48400;
  assign n48386 = n48402 ^ n45763;
  assign n48403 = ~n48402;
  assign n46912 = ~n48157;
  assign n48337 = ~n48373;
  assign n48374 = n48378 & n48379;
  assign n48360 = n48380 ^ n48381;
  assign n48321 = n48384 & n48385;
  assign n44523 = n48386 ^ n48387;
  assign n48382 = ~n48380;
  assign n48394 = n48403 & n48404;
  assign n48320 = n48359 ^ n48360;
  assign n48365 = n44523 & n47096;
  assign n48366 = n48321 & n48372;
  assign n48351 = ~n48374;
  assign n48363 = ~n48321;
  assign n44566 = ~n44523;
  assign n48375 = n48382 & n48383;
  assign n48388 = ~n48394;
  assign n48339 = n48320 & n462;
  assign n48333 = n48351 ^ n48352;
  assign n48338 = ~n48320;
  assign n48350 = n48358 & n48351;
  assign n48353 = n48363 & n48341;
  assign n48354 = n44566 & n48364;
  assign n47117 = ~n48365;
  assign n48355 = n44566 & n47025;
  assign n48343 = ~n48366;
  assign n48356 = n44566 & n45763;
  assign n48361 = ~n48375;
  assign n48367 = n48388 & n48389;
  assign n48310 = n463 ^ n48333;
  assign n48334 = n48338 & n18263;
  assign n48296 = ~n48339;
  assign n48336 = ~n48350;
  assign n48324 = ~n48353;
  assign n47098 = ~n48354;
  assign n48344 = ~n48355;
  assign n47059 = ~n48356;
  assign n48340 = n48361 & n48362;
  assign n48347 = n48367 ^ n45723;
  assign n48368 = ~n48367;
  assign n48116 = n48309 ^ n48310;
  assign n48274 = n48310 & n48309;
  assign n48317 = ~n48334;
  assign n48319 = n48336 & n48337;
  assign n48322 = n48340 ^ n48341;
  assign n48280 = n48344 & n48345;
  assign n44455 = n48346 ^ n48347;
  assign n48342 = ~n48340;
  assign n48357 = n48368 & n48369;
  assign n46872 = ~n48116;
  assign n48294 = n48319 ^ n48320;
  assign n48277 = n48321 ^ n48322;
  assign n48326 = n48280 & n48331;
  assign n48327 = n44455 & n48332;
  assign n48318 = ~n48319;
  assign n48325 = ~n48280;
  assign n44489 = ~n44455;
  assign n48335 = n48342 & n48343;
  assign n48348 = ~n48357;
  assign n48275 = n462 ^ n48294;
  assign n48298 = n48277 & n461;
  assign n48297 = ~n48277;
  assign n48311 = n48317 & n48318;
  assign n48312 = n48325 & n48300;
  assign n48313 = n44489 & n47060;
  assign n48314 = n44489 & n46987;
  assign n48304 = ~n48326;
  assign n47084 = ~n48327;
  assign n48315 = n44489 & n45710;
  assign n48323 = ~n48335;
  assign n48328 = n48348 & n48349;
  assign n48076 = n48274 ^ n48275;
  assign n48233 = n48275 & n48274;
  assign n48292 = n48297 & n18218;
  assign n48255 = ~n48298;
  assign n48295 = ~n48311;
  assign n48283 = ~n48312;
  assign n47065 = ~n48313;
  assign n48301 = ~n48314;
  assign n47030 = ~n48315;
  assign n48299 = n48323 & n48324;
  assign n48305 = n48328 ^ n45690;
  assign n48329 = ~n48328;
  assign n46828 = ~n48076;
  assign n48279 = ~n48292;
  assign n48276 = n48295 & n48296;
  assign n48281 = n48299 ^ n48300;
  assign n48231 = n48301 & n48302;
  assign n44387 = n48305 ^ n48306;
  assign n48303 = ~n48299;
  assign n48316 = n48329 & n48330;
  assign n48253 = n48276 ^ n48277;
  assign n48236 = n48280 ^ n48281;
  assign n48286 = n44387 & n47022;
  assign n48287 = n48231 & n48291;
  assign n48278 = ~n48276;
  assign n48284 = ~n48231;
  assign n44401 = ~n44387;
  assign n48293 = n48303 & n48304;
  assign n48307 = ~n48316;
  assign n48234 = n461 ^ n48253;
  assign n48257 = n48236 & n460;
  assign n48256 = ~n48236;
  assign n48268 = n48278 & n48279;
  assign n48269 = n48284 & n48259;
  assign n48270 = n44401 & n48285;
  assign n47048 = ~n48286;
  assign n48271 = n44401 & n46969;
  assign n48263 = ~n48287;
  assign n48272 = n44401 & n45690;
  assign n48282 = ~n48293;
  assign n48288 = n48307 & n48308;
  assign n46787 = n48233 ^ n48234;
  assign n48186 = n48234 & n48233;
  assign n48251 = n48256 & n18199;
  assign n48214 = ~n48257;
  assign n48254 = ~n48268;
  assign n48240 = ~n48269;
  assign n47027 = ~n48270;
  assign n48260 = ~n48271;
  assign n46991 = ~n48272;
  assign n48258 = n48282 & n48283;
  assign n48265 = n48288 ^ n45633;
  assign n48289 = ~n48288;
  assign n48041 = ~n46787;
  assign n48189 = ~n48186;
  assign n48238 = ~n48251;
  assign n48235 = n48254 & n48255;
  assign n48232 = n48258 ^ n48259;
  assign n48194 = n48260 & n48261;
  assign n44327 = n48264 ^ n48265;
  assign n48262 = ~n48258;
  assign n48273 = n48289 & n48290;
  assign n48191 = n48231 ^ n48232;
  assign n48212 = n48235 ^ n48236;
  assign n48243 = n44327 & n46993;
  assign n48245 = n44327 & n46938;
  assign n48246 = n48194 & n48218;
  assign n48247 = n44327 & n45633;
  assign n48237 = ~n48235;
  assign n48241 = ~n48194;
  assign n44362 = ~n44327;
  assign n48252 = n48262 & n48263;
  assign n48266 = ~n48273;
  assign n48187 = n460 ^ n48212;
  assign n48216 = n48191 & n459;
  assign n48215 = ~n48191;
  assign n48227 = n48237 & n48238;
  assign n48228 = n48241 & n48242;
  assign n46995 = ~n48243;
  assign n48229 = n44362 & n48244;
  assign n48225 = ~n48245;
  assign n48220 = ~n48246;
  assign n46957 = ~n48247;
  assign n48239 = ~n48252;
  assign n48248 = n48266 & n48267;
  assign n46746 = n48186 ^ n48187;
  assign n48188 = ~n48187;
  assign n48209 = n48215 & n18144;
  assign n48170 = ~n48216;
  assign n48151 = n48225 & n48226;
  assign n48213 = ~n48227;
  assign n48197 = ~n48228;
  assign n47009 = ~n48229;
  assign n48217 = n48239 & n48240;
  assign n48221 = n48248 ^ n45601;
  assign n48249 = ~n48248;
  assign n48001 = ~n46746;
  assign n48144 = n48188 & n48189;
  assign n48193 = ~n48209;
  assign n48208 = n48151 & n48210;
  assign n48190 = n48213 & n48214;
  assign n48195 = n48217 ^ n48218;
  assign n48207 = ~n48151;
  assign n44270 = n48221 ^ n48222;
  assign n48219 = ~n48217;
  assign n48230 = n48249 & n48250;
  assign n48168 = n48190 ^ n48191;
  assign n48148 = n48194 ^ n48195;
  assign n48198 = n48207 & n48174;
  assign n48199 = n44270 & n46866;
  assign n48176 = ~n48208;
  assign n48201 = n44270 & n46953;
  assign n48202 = n44270 & n45601;
  assign n48192 = ~n48190;
  assign n44302 = ~n44270;
  assign n48211 = n48219 & n48220;
  assign n48223 = ~n48230;
  assign n48145 = n459 ^ n48168;
  assign n48171 = n48148 & n18124;
  assign n48172 = ~n48148;
  assign n48183 = n48192 & n48193;
  assign n48154 = ~n48198;
  assign n48181 = ~n48199;
  assign n48184 = n44302 & n48200;
  assign n46955 = ~n48201;
  assign n46917 = ~n48202;
  assign n48196 = ~n48211;
  assign n48203 = n48223 & n48224;
  assign n46703 = n48144 ^ n48145;
  assign n48146 = ~n48145;
  assign n48150 = ~n48171;
  assign n48165 = n48172 & n458;
  assign n48110 = n48181 & n48182;
  assign n48169 = ~n48183;
  assign n46975 = ~n48184;
  assign n48173 = n48196 & n48197;
  assign n48177 = n48203 ^ n48204;
  assign n48205 = ~n48203;
  assign n47961 = ~n46703;
  assign n48104 = n48146 & n48144;
  assign n48128 = ~n48165;
  assign n48164 = n48110 & n48166;
  assign n48147 = n48169 & n48170;
  assign n48152 = n48173 ^ n48174;
  assign n48163 = ~n48110;
  assign n44202 = n45547 ^ n48177;
  assign n48178 = n48177 & n45489;
  assign n48175 = ~n48173;
  assign n48185 = n48205 & n48206;
  assign n48126 = n48147 ^ n48148;
  assign n48107 = n48151 ^ n48152;
  assign n48155 = n48163 & n48132;
  assign n48156 = n44202 & n46849;
  assign n48134 = ~n48164;
  assign n48158 = n44202 & n46912;
  assign n48149 = ~n48147;
  assign n44253 = ~n44202;
  assign n48167 = n48175 & n48176;
  assign n46868 = ~n48178;
  assign n48179 = ~n48185;
  assign n48105 = n458 ^ n48126;
  assign n48130 = n48107 & n457;
  assign n48129 = ~n48107;
  assign n48141 = n48149 & n48150;
  assign n48113 = ~n48155;
  assign n48139 = ~n48156;
  assign n48142 = n44253 & n48157;
  assign n46915 = ~n48158;
  assign n48153 = ~n48167;
  assign n48159 = n48179 & n48180;
  assign n46666 = n48104 ^ n48105;
  assign n48062 = n48105 & n48104;
  assign n48124 = n48129 & n18059;
  assign n48088 = ~n48130;
  assign n48092 = n48139 & n48140;
  assign n48127 = ~n48141;
  assign n46936 = ~n48142;
  assign n48131 = n48153 & n48154;
  assign n48135 = n48159 ^ n48160;
  assign n48161 = ~n48159;
  assign n47909 = ~n46666;
  assign n48109 = ~n48124;
  assign n48123 = n48092 & n48070;
  assign n48106 = n48127 & n48128;
  assign n48111 = n48131 ^ n48132;
  assign n48121 = ~n48092;
  assign n44162 = n45503 ^ n48135;
  assign n48136 = n48135 & n45465;
  assign n48133 = ~n48131;
  assign n48143 = n48161 & n48162;
  assign n48086 = n48106 ^ n48107;
  assign n48066 = n48110 ^ n48111;
  assign n48114 = n48121 & n48122;
  assign n48115 = n44162 & n46813;
  assign n48093 = ~n48123;
  assign n48117 = n44162 & n46872;
  assign n48108 = ~n48106;
  assign n44191 = ~n44162;
  assign n48125 = n48133 & n48134;
  assign n46833 = ~n48136;
  assign n48137 = ~n48143;
  assign n48063 = n457 ^ n48086;
  assign n48090 = n48066 & n456;
  assign n48089 = ~n48066;
  assign n48101 = n48108 & n48109;
  assign n48072 = ~n48114;
  assign n48099 = ~n48115;
  assign n48102 = n44191 & n48116;
  assign n46874 = ~n48117;
  assign n48112 = ~n48125;
  assign n48118 = n48137 & n48138;
  assign n46620 = n48062 ^ n48063;
  assign n48064 = ~n48063;
  assign n48083 = n48089 & n18051;
  assign n48046 = ~n48090;
  assign n48050 = n48099 & n48100;
  assign n48087 = ~n48101;
  assign n46897 = ~n48102;
  assign n48091 = n48112 & n48113;
  assign n48096 = n48118 ^ n45411;
  assign n48119 = ~n48118;
  assign n47883 = ~n46620;
  assign n48027 = n48064 & n48062;
  assign n48068 = ~n48083;
  assign n48082 = n48050 & n48084;
  assign n48065 = n48087 & n48088;
  assign n48069 = n48091 ^ n48092;
  assign n48081 = ~n48050;
  assign n44132 = n48095 ^ n48096;
  assign n48094 = ~n48091;
  assign n48103 = n48119 & n48120;
  assign n48044 = n48065 ^ n48066;
  assign n48008 = n48069 ^ n48070;
  assign n48073 = n48081 & n48032;
  assign n48051 = ~n48082;
  assign n48074 = n44132 & n46772;
  assign n48075 = n44132 & n46828;
  assign n48077 = n44132 & n45411;
  assign n48067 = ~n48065;
  assign n44172 = ~n44132;
  assign n48085 = n48093 & n48094;
  assign n48097 = ~n48103;
  assign n48028 = n456 ^ n48044;
  assign n48047 = n48008 & n17983;
  assign n48048 = ~n48008;
  assign n48059 = n48067 & n48068;
  assign n48034 = ~n48073;
  assign n48057 = ~n48074;
  assign n46830 = ~n48075;
  assign n48060 = n44172 & n48076;
  assign n46792 = ~n48077;
  assign n48071 = ~n48085;
  assign n48078 = n48097 & n48098;
  assign n46599 = n48027 ^ n48028;
  assign n48029 = ~n48028;
  assign n48025 = ~n48047;
  assign n48042 = n48048 & n471;
  assign n47989 = n48057 & n48058;
  assign n48045 = ~n48059;
  assign n46856 = ~n48060;
  assign n48049 = n48071 & n48072;
  assign n48054 = n48078 ^ n45343;
  assign n48079 = ~n48078;
  assign n47841 = ~n46599;
  assign n47981 = n48029 & n48027;
  assign n48006 = ~n48042;
  assign n48030 = n48045 & n48046;
  assign n48031 = n48049 ^ n48050;
  assign n47998 = ~n47989;
  assign n44096 = n48053 ^ n48054;
  assign n48052 = ~n48049;
  assign n48061 = n48079 & n48080;
  assign n47984 = ~n47981;
  assign n48007 = n471 ^ n48030;
  assign n47986 = n48031 ^ n48032;
  assign n48035 = n44096 & n46699;
  assign n48036 = n44096 & n48041;
  assign n48037 = n44096 & n45343;
  assign n48026 = ~n48030;
  assign n44115 = ~n44096;
  assign n48043 = n48051 & n48052;
  assign n48055 = ~n48061;
  assign n47982 = n48007 ^ n48008;
  assign n48010 = n47986 & n470;
  assign n48009 = ~n47986;
  assign n48022 = n48025 & n48026;
  assign n48019 = ~n48035;
  assign n46790 = ~n48036;
  assign n46751 = ~n48037;
  assign n48023 = n44115 & n46787;
  assign n48033 = ~n48043;
  assign n48038 = n48055 & n48056;
  assign n46545 = n47981 ^ n47982;
  assign n47983 = ~n47982;
  assign n48002 = n48009 & n17956;
  assign n47965 = ~n48010;
  assign n47931 = n48019 & n48020;
  assign n48005 = ~n48022;
  assign n46811 = ~n48023;
  assign n48011 = n48033 & n48034;
  assign n48015 = n48038 ^ n45328;
  assign n48039 = ~n48038;
  assign n47798 = ~n46545;
  assign n47941 = n47983 & n47984;
  assign n47987 = ~n48002;
  assign n48000 = n47931 & n48003;
  assign n47985 = n48005 & n48006;
  assign n47990 = n48011 ^ n48012;
  assign n47999 = ~n47931;
  assign n44061 = n48015 ^ n48016;
  assign n48014 = n48011 & n48021;
  assign n48013 = ~n48011;
  assign n48024 = n48039 & n48040;
  assign n47963 = n47985 ^ n47986;
  assign n47944 = n47989 ^ n47990;
  assign n47992 = n47999 & n47958;
  assign n47960 = ~n48000;
  assign n47993 = n44061 & n48001;
  assign n47988 = ~n47985;
  assign n44063 = ~n44061;
  assign n48004 = n48013 & n48012;
  assign n47997 = ~n48014;
  assign n48017 = ~n48024;
  assign n47942 = n470 ^ n47963;
  assign n47967 = n47944 & n469;
  assign n47966 = ~n47944;
  assign n47976 = n47987 & n47988;
  assign n47934 = ~n47992;
  assign n47977 = n44063 & n46688;
  assign n46770 = ~n47993;
  assign n47978 = n44063 & n46746;
  assign n47979 = n44063 & n45328;
  assign n47991 = n47997 & n47998;
  assign n47975 = ~n48004;
  assign n47994 = n48017 & n48018;
  assign n46458 = n47941 ^ n47942;
  assign n47901 = n47942 & n47941;
  assign n47962 = n47966 & n17901;
  assign n47926 = ~n47967;
  assign n47964 = ~n47976;
  assign n47968 = ~n47977;
  assign n46749 = ~n47978;
  assign n46707 = ~n47979;
  assign n47974 = ~n47991;
  assign n47971 = n47994 ^ n45157;
  assign n47995 = ~n47994;
  assign n47746 = ~n46458;
  assign n47945 = ~n47962;
  assign n47943 = n47964 & n47965;
  assign n47893 = n47968 & n47969;
  assign n44003 = n47970 ^ n47971;
  assign n47957 = n47974 & n47975;
  assign n47980 = n47995 & n47996;
  assign n47924 = n47943 ^ n47944;
  assign n47932 = n47957 ^ n47958;
  assign n47950 = n47893 & n47918;
  assign n47951 = n44003 & n46616;
  assign n47952 = n44003 & n47961;
  assign n47953 = n44003 & n45258;
  assign n47946 = ~n47943;
  assign n47948 = ~n47893;
  assign n44028 = ~n44003;
  assign n47959 = ~n47957;
  assign n47972 = ~n47980;
  assign n47902 = n469 ^ n47924;
  assign n47904 = n47931 ^ n47932;
  assign n47937 = n47945 & n47946;
  assign n47938 = n47948 & n47949;
  assign n47920 = ~n47950;
  assign n47935 = ~n47951;
  assign n47939 = n44028 & n46703;
  assign n46705 = ~n47952;
  assign n46662 = ~n47953;
  assign n47947 = n47959 & n47960;
  assign n47954 = n47972 & n47973;
  assign n46395 = n47901 ^ n47902;
  assign n47862 = n47902 & n47901;
  assign n47916 = n47904 & n468;
  assign n47915 = ~n47904;
  assign n47848 = n47935 & n47936;
  assign n47925 = ~n47937;
  assign n47898 = ~n47938;
  assign n46730 = ~n47939;
  assign n47933 = ~n47947;
  assign n47928 = n47954 ^ n45113;
  assign n47955 = ~n47954;
  assign n47718 = ~n46395;
  assign n47861 = ~n47862;
  assign n47905 = n47915 & n17859;
  assign n47874 = ~n47916;
  assign n47922 = n47848 & n47923;
  assign n47903 = n47925 & n47926;
  assign n47921 = ~n47848;
  assign n43964 = n47927 ^ n47928;
  assign n47917 = n47933 & n47934;
  assign n47940 = n47955 & n47956;
  assign n47885 = n47903 ^ n47904;
  assign n47891 = ~n47905;
  assign n47894 = n47917 ^ n47918;
  assign n47907 = n47921 & n47878;
  assign n47880 = ~n47922;
  assign n47908 = n43964 & n46565;
  assign n47910 = n43964 & n45113;
  assign n47911 = n43964 & n46666;
  assign n47892 = ~n47903;
  assign n43989 = ~n43964;
  assign n47919 = ~n47917;
  assign n47929 = ~n47940;
  assign n47863 = n468 ^ n47885;
  assign n47886 = n47891 & n47892;
  assign n47851 = n47893 ^ n47894;
  assign n47855 = ~n47907;
  assign n47895 = ~n47908;
  assign n47899 = n43989 & n47909;
  assign n46624 = ~n47910;
  assign n46668 = ~n47911;
  assign n47906 = n47919 & n47920;
  assign n47912 = n47929 & n47930;
  assign n46325 = n47862 ^ n47863;
  assign n47860 = ~n47863;
  assign n47875 = n47851 & n17816;
  assign n47873 = ~n47886;
  assign n47876 = ~n47851;
  assign n47812 = n47895 & n47896;
  assign n46685 = ~n47899;
  assign n47897 = ~n47906;
  assign n47887 = n47912 ^ n45056;
  assign n47913 = ~n47912;
  assign n47660 = ~n46325;
  assign n47806 = n47860 & n47861;
  assign n47850 = n47873 & n47874;
  assign n47853 = ~n47875;
  assign n47864 = n47876 & n467;
  assign n47882 = n47812 & n47884;
  assign n47881 = ~n47812;
  assign n43922 = n47887 ^ n47888;
  assign n47877 = n47897 & n47898;
  assign n47900 = n47913 & n47914;
  assign n47832 = n47850 ^ n47851;
  assign n47809 = ~n47806;
  assign n47852 = ~n47850;
  assign n47831 = ~n47864;
  assign n47849 = n47877 ^ n47878;
  assign n47866 = n47881 & n47836;
  assign n47838 = ~n47882;
  assign n47867 = n43922 & n46512;
  assign n47868 = n43922 & n47883;
  assign n47869 = n43922 & n45056;
  assign n43944 = ~n43922;
  assign n47879 = ~n47877;
  assign n47889 = ~n47900;
  assign n47807 = n467 ^ n47832;
  assign n47811 = n47848 ^ n47849;
  assign n47843 = n47852 & n47853;
  assign n47815 = ~n47866;
  assign n47856 = ~n47867;
  assign n46622 = ~n47868;
  assign n46567 = ~n47869;
  assign n47858 = n43944 & n46620;
  assign n47865 = n47879 & n47880;
  assign n47870 = n47889 & n47890;
  assign n47625 = n47806 ^ n47807;
  assign n47808 = ~n47807;
  assign n47834 = n47811 & n466;
  assign n47830 = ~n47843;
  assign n47833 = ~n47811;
  assign n47770 = n47856 & n47857;
  assign n46648 = ~n47858;
  assign n47854 = ~n47865;
  assign n47845 = n47870 ^ n44891;
  assign n47871 = ~n47870;
  assign n46243 = ~n47625;
  assign n47764 = n47808 & n47809;
  assign n47810 = n47830 & n47831;
  assign n47820 = n47833 & n17747;
  assign n47788 = ~n47834;
  assign n47840 = n47770 & n47842;
  assign n47839 = ~n47770;
  assign n43869 = n47844 ^ n47845;
  assign n47835 = n47854 & n47855;
  assign n47859 = n47871 & n47872;
  assign n47786 = n47810 ^ n47811;
  assign n47804 = ~n47810;
  assign n47805 = ~n47820;
  assign n47813 = n47835 ^ n47836;
  assign n47822 = n47839 & n47792;
  assign n47823 = n43869 & n46422;
  assign n47794 = ~n47840;
  assign n47824 = n43869 & n47841;
  assign n47825 = n43869 & n44891;
  assign n43929 = ~n43869;
  assign n47837 = ~n47835;
  assign n47846 = ~n47859;
  assign n47765 = n466 ^ n47786;
  assign n47799 = n47804 & n47805;
  assign n47767 = n47812 ^ n47813;
  assign n47775 = ~n47822;
  assign n47816 = ~n47823;
  assign n47818 = n43929 & n46599;
  assign n46573 = ~n47824;
  assign n46521 = ~n47825;
  assign n47821 = n47837 & n47838;
  assign n47826 = n47846 & n47847;
  assign n46164 = n47764 ^ n47765;
  assign n47727 = n47765 & n47764;
  assign n47790 = n47767 & n465;
  assign n47787 = ~n47799;
  assign n47789 = ~n47767;
  assign n47756 = n47816 & n47817;
  assign n46601 = ~n47818;
  assign n47814 = ~n47821;
  assign n47800 = n47826 ^ n47827;
  assign n47828 = ~n47826;
  assign n47572 = ~n46164;
  assign n47730 = ~n47727;
  assign n47766 = n47787 & n47788;
  assign n47778 = n47789 & n17696;
  assign n47753 = ~n47790;
  assign n47797 = n47756 & n47736;
  assign n47795 = ~n47756;
  assign n43846 = n44851 ^ n47800;
  assign n47791 = n47814 & n47815;
  assign n47801 = n47800 & n44946;
  assign n47819 = n47828 & n47829;
  assign n47751 = n47766 ^ n47767;
  assign n47769 = ~n47778;
  assign n47768 = ~n47766;
  assign n47771 = n47791 ^ n47792;
  assign n47780 = n47795 & n47796;
  assign n47758 = ~n47797;
  assign n47781 = n43846 & n46435;
  assign n47782 = n43846 & n47798;
  assign n43852 = ~n43846;
  assign n47793 = ~n47791;
  assign n46465 = ~n47801;
  assign n47802 = ~n47819;
  assign n47728 = n465 ^ n47751;
  assign n47759 = n47768 & n47769;
  assign n47732 = n47770 ^ n47771;
  assign n47738 = ~n47780;
  assign n47772 = ~n47781;
  assign n46518 = ~n47782;
  assign n47776 = n43852 & n46545;
  assign n47779 = n47793 & n47794;
  assign n47783 = n47802 & n47803;
  assign n46085 = n47727 ^ n47728;
  assign n47729 = ~n47728;
  assign n47754 = n47732 & n464;
  assign n47752 = ~n47759;
  assign n47750 = ~n47732;
  assign n47713 = n47772 & n47773;
  assign n46547 = ~n47776;
  assign n47774 = ~n47779;
  assign n47761 = n47783 ^ n44768;
  assign n47784 = ~n47783;
  assign n47682 = n47729 & n47730;
  assign n47743 = n47750 & n17666;
  assign n47731 = n47752 & n47753;
  assign n47710 = ~n47754;
  assign n47694 = ~n47713;
  assign n43792 = n47760 ^ n47761;
  assign n47755 = n47774 & n47775;
  assign n47777 = n47784 & n47785;
  assign n47708 = n47731 ^ n47732;
  assign n47733 = ~n47731;
  assign n47734 = ~n47743;
  assign n47735 = n47755 ^ n47756;
  assign n47745 = n43792 & n46458;
  assign n43830 = ~n43792;
  assign n47757 = ~n47755;
  assign n47762 = ~n47777;
  assign n47683 = n464 ^ n47708;
  assign n47720 = n47733 & n47734;
  assign n47667 = n47735 ^ n47736;
  assign n47739 = n43830 & n46361;
  assign n46492 = ~n47745;
  assign n47740 = n43830 & n44768;
  assign n47741 = n43830 & n47746;
  assign n47744 = n47757 & n47758;
  assign n47747 = n47762 & n47763;
  assign n47664 = n47682 ^ n47683;
  assign n47684 = ~n47683;
  assign n47711 = n47667 & n17570;
  assign n47709 = ~n47720;
  assign n47712 = ~n47667;
  assign n47721 = ~n47739;
  assign n46392 = ~n47740;
  assign n46461 = ~n47741;
  assign n47737 = ~n47744;
  assign n47723 = n47747 ^ n44786;
  assign n47748 = ~n47747;
  assign n43600 = n47664 ^ n45539;
  assign n47665 = ~n47664;
  assign n47637 = n47684 & n47682;
  assign n47685 = n47709 & n47710;
  assign n47687 = ~n47711;
  assign n47698 = n47712 & n479;
  assign n47627 = n47721 & n47722;
  assign n43789 = n47723 ^ n47724;
  assign n47714 = n47737 & n47738;
  assign n47742 = n47748 & n47749;
  assign n43602 = ~n43600;
  assign n47567 = n47665 & n45539;
  assign n47654 = n47665 & n45535;
  assign n47640 = ~n47637;
  assign n47666 = n479 ^ n47685;
  assign n47686 = ~n47685;
  assign n47669 = ~n47698;
  assign n47688 = n47713 ^ n47714;
  assign n47701 = n47627 & n47716;
  assign n47702 = n43789 & n47718;
  assign n47703 = n43789 & n44786;
  assign n47704 = n43789 & n46240;
  assign n47717 = n47714 & n47719;
  assign n47699 = ~n47627;
  assign n43750 = ~n43789;
  assign n47715 = ~n47714;
  assign n47725 = ~n47742;
  assign n47631 = n43602 & n46551;
  assign n46575 = ~n47654;
  assign n47638 = n47666 ^ n47667;
  assign n47677 = n47686 & n47687;
  assign n47642 = n47688 ^ n47689;
  assign n47695 = n47699 & n47649;
  assign n47651 = ~n47701;
  assign n46398 = ~n47702;
  assign n47696 = n43750 & n46395;
  assign n46337 = ~n47703;
  assign n47690 = ~n47704;
  assign n47700 = n47715 & n47689;
  assign n47693 = ~n47717;
  assign n47705 = n47725 & n47726;
  assign n47615 = ~n47631;
  assign n47626 = n47637 ^ n47638;
  assign n47639 = ~n47638;
  assign n47671 = n47642 & n478;
  assign n47668 = ~n47677;
  assign n47670 = ~n47642;
  assign n47577 = n47690 & n47691;
  assign n47692 = n47693 & n47694;
  assign n47630 = ~n47695;
  assign n46429 = ~n47696;
  assign n47676 = ~n47700;
  assign n47679 = n47705 ^ n44689;
  assign n47706 = ~n47705;
  assign n47587 = n47615 & n47616;
  assign n47617 = n47626 & n45509;
  assign n47618 = ~n47626;
  assign n47593 = n47639 & n47640;
  assign n47641 = n47668 & n47669;
  assign n47655 = n47670 & n17477;
  assign n47621 = ~n47671;
  assign n47674 = n47577 & n47602;
  assign n47672 = ~n47577;
  assign n43709 = n47678 ^ n47679;
  assign n47675 = ~n47692;
  assign n47697 = n47706 & n47707;
  assign n47565 = n47587 ^ n47588;
  assign n47589 = ~n47587;
  assign n47592 = ~n47617;
  assign n47609 = n47618 & n45520;
  assign n47619 = n47641 ^ n47642;
  assign n47643 = ~n47641;
  assign n47644 = ~n47655;
  assign n47656 = n47672 & n47673;
  assign n47604 = ~n47674;
  assign n47657 = n43709 & n46161;
  assign n47658 = n43709 & n46325;
  assign n47659 = n43709 & n44689;
  assign n47648 = n47675 & n47676;
  assign n43753 = ~n43709;
  assign n47680 = ~n47697;
  assign n45676 = n103 ^ n47565;
  assign n47367 = n47565 & n103;
  assign n47445 = n47589 & n47590;
  assign n47591 = n47592 & n47567;
  assign n47574 = ~n47609;
  assign n47594 = n478 ^ n47619;
  assign n47632 = n47643 & n47644;
  assign n47628 = n47648 ^ n47649;
  assign n47580 = ~n47656;
  assign n47646 = ~n47657;
  assign n46327 = ~n47658;
  assign n46260 = ~n47659;
  assign n47652 = n43753 & n47660;
  assign n47650 = ~n47648;
  assign n47661 = n47680 & n47681;
  assign n45706 = ~n45676;
  assign n47573 = ~n47591;
  assign n47566 = n47592 & n47574;
  assign n47519 = n47593 ^ n47594;
  assign n47536 = n47594 & n47593;
  assign n47596 = n47627 ^ n47628;
  assign n47620 = ~n47632;
  assign n47527 = n47646 & n47647;
  assign n47645 = n47650 & n47651;
  assign n46369 = ~n47652;
  assign n47633 = n47661 ^ n44602;
  assign n47662 = ~n47661;
  assign n43547 = n47566 ^ n47567;
  assign n47546 = n47573 & n47574;
  assign n47568 = n47519 & n45365;
  assign n47569 = ~n47519;
  assign n47539 = ~n47536;
  assign n47600 = n47596 & n477;
  assign n47595 = n47620 & n47621;
  assign n47599 = ~n47596;
  assign n47624 = n47527 & n47552;
  assign n47622 = ~n47527;
  assign n43672 = n47633 ^ n47634;
  assign n47629 = ~n47645;
  assign n47653 = n47662 & n47663;
  assign n47533 = n43547 & n46432;
  assign n47534 = n43547 & n45509;
  assign n47520 = n47546 ^ n45367;
  assign n43551 = ~n43547;
  assign n47545 = ~n47546;
  assign n47544 = ~n47568;
  assign n47557 = n47569 & n45367;
  assign n47570 = n47595 ^ n47596;
  assign n47597 = n47599 & n17431;
  assign n47548 = ~n47600;
  assign n47576 = ~n47595;
  assign n47610 = n47622 & n47623;
  assign n47554 = ~n47624;
  assign n47611 = n43672 & n47625;
  assign n47601 = n47629 & n47630;
  assign n43698 = ~n43672;
  assign n47635 = ~n47653;
  assign n43521 = n47519 ^ n47520;
  assign n47517 = ~n47533;
  assign n46463 = ~n47534;
  assign n47535 = n47544 & n47545;
  assign n47522 = ~n47557;
  assign n47537 = n477 ^ n47570;
  assign n47575 = ~n47597;
  assign n47578 = n47601 ^ n47602;
  assign n47530 = ~n47610;
  assign n47605 = n43698 & n46082;
  assign n47606 = n43698 & n44602;
  assign n46291 = ~n47611;
  assign n47607 = n43698 & n46243;
  assign n47603 = ~n47601;
  assign n47612 = n47635 & n47636;
  assign n47495 = n43521 & n46371;
  assign n47496 = n43521 & n45365;
  assign n43510 = ~n43521;
  assign n47508 = n47517 & n47518;
  assign n47521 = ~n47535;
  assign n47469 = n47536 ^ n47537;
  assign n47538 = ~n47537;
  assign n47571 = n47575 & n47576;
  assign n47524 = n47577 ^ n47578;
  assign n47598 = n47603 & n47604;
  assign n47581 = ~n47605;
  assign n46178 = ~n47606;
  assign n46246 = ~n47607;
  assign n47583 = n47612 ^ n44528;
  assign n47613 = ~n47612;
  assign n47483 = ~n47495;
  assign n46400 = ~n47496;
  assign n47497 = n47508 & n47509;
  assign n47493 = ~n47508;
  assign n47498 = n47521 & n47522;
  assign n47514 = n47469 & n45282;
  assign n47513 = ~n47469;
  assign n47473 = n47538 & n47539;
  assign n47549 = n47524 & n17352;
  assign n47547 = ~n47571;
  assign n47550 = ~n47524;
  assign n47479 = n47581 & n47582;
  assign n43642 = n47583 ^ n47584;
  assign n47579 = ~n47598;
  assign n47608 = n47613 & n47614;
  assign n47403 = n47483 & n47484;
  assign n47486 = n47493 & n47494;
  assign n47472 = ~n47497;
  assign n47470 = n47498 ^ n45280;
  assign n47487 = ~n47498;
  assign n47510 = n47513 & n45280;
  assign n47464 = ~n47514;
  assign n47523 = n47547 & n47548;
  assign n47526 = ~n47549;
  assign n47540 = n47550 & n476;
  assign n47560 = n47479 & n47505;
  assign n47561 = n43642 & n46063;
  assign n47562 = n43642 & n44528;
  assign n47563 = n43642 & n47572;
  assign n47551 = n47579 & n47580;
  assign n47558 = ~n47479;
  assign n43648 = ~n43642;
  assign n47585 = ~n47608;
  assign n47458 = n47403 & n47465;
  assign n47457 = ~n47403;
  assign n43481 = n47469 ^ n47470;
  assign n47471 = n47472 & n47445;
  assign n47460 = ~n47486;
  assign n47488 = ~n47510;
  assign n47499 = n47523 ^ n47524;
  assign n47525 = ~n47523;
  assign n47501 = ~n47540;
  assign n47528 = n47551 ^ n47552;
  assign n47555 = n47558 & n47559;
  assign n47507 = ~n47560;
  assign n47542 = ~n47561;
  assign n46099 = ~n47562;
  assign n47556 = n43648 & n46164;
  assign n46167 = ~n47563;
  assign n47553 = ~n47551;
  assign n47564 = n47585 & n47586;
  assign n47441 = n47457 & n47435;
  assign n47429 = ~n47458;
  assign n47442 = n43481 & n46262;
  assign n47443 = n43481 & n45280;
  assign n43493 = ~n43481;
  assign n47459 = ~n47471;
  assign n47444 = n47460 & n47472;
  assign n47485 = n47487 & n47488;
  assign n47474 = n476 ^ n47499;
  assign n47515 = n47525 & n47526;
  assign n47476 = n47527 ^ n47528;
  assign n47426 = n47542 & n47543;
  assign n47541 = n47553 & n47554;
  assign n47482 = ~n47555;
  assign n46209 = ~n47556;
  assign n47532 = n47564 ^ n47516;
  assign n47402 = ~n47441;
  assign n47431 = ~n47442;
  assign n46330 = ~n47443;
  assign n47433 = n47444 ^ n47445;
  assign n47434 = n47459 & n47460;
  assign n47407 = n47473 ^ n47474;
  assign n47463 = ~n47485;
  assign n47420 = n47474 & n47473;
  assign n47502 = n47476 & n17233;
  assign n47500 = ~n47515;
  assign n47503 = ~n47476;
  assign n47437 = ~n47426;
  assign n43634 = n47531 ^ n47532;
  assign n47529 = ~n47541;
  assign n47355 = n47431 & n47432;
  assign n47417 = n47433 & n102;
  assign n47404 = n47434 ^ n47435;
  assign n47416 = ~n47433;
  assign n47430 = ~n47434;
  assign n47446 = n47407 & n45188;
  assign n47461 = n47463 & n47464;
  assign n47447 = ~n47407;
  assign n47475 = n47500 & n47501;
  assign n47478 = ~n47502;
  assign n47489 = n47503 & n475;
  assign n47511 = n43634 & n45973;
  assign n47512 = n43634 & n47516;
  assign n47504 = n47529 & n47530;
  assign n44569 = ~n43634;
  assign n47343 = n47403 ^ n47404;
  assign n47406 = n47355 & n47411;
  assign n47405 = ~n47355;
  assign n47412 = n47416 & n14810;
  assign n47364 = ~n47417;
  assign n47415 = n47429 & n47430;
  assign n47393 = ~n47446;
  assign n47438 = n47447 & n45179;
  assign n47418 = ~n47461;
  assign n47448 = n47475 ^ n47476;
  assign n47477 = ~n47475;
  assign n47450 = ~n47489;
  assign n47480 = n47504 ^ n47505;
  assign n47491 = ~n47511;
  assign n46015 = ~n47512;
  assign n47506 = ~n47504;
  assign n47381 = n47343 & n101;
  assign n47380 = ~n47343;
  assign n47390 = n47405 & n47383;
  assign n47384 = ~n47406;
  assign n47391 = ~n47412;
  assign n47401 = ~n47415;
  assign n47408 = n47418 ^ n45179;
  assign n47419 = ~n47438;
  assign n47421 = n475 ^ n47448;
  assign n47466 = n47477 & n47478;
  assign n47423 = n47479 ^ n47480;
  assign n47467 = n47491 & n47492;
  assign n47490 = n47506 & n47507;
  assign n47365 = n47380 & n14752;
  assign n47319 = ~n47381;
  assign n47358 = ~n47390;
  assign n47387 = n47391 & n47367;
  assign n47366 = n47391 & n47364;
  assign n47382 = n47401 & n47402;
  assign n43438 = n47407 ^ n47408;
  assign n47413 = n47418 & n47419;
  assign n47344 = n47420 ^ n47421;
  assign n47374 = n47421 & n47420;
  assign n47451 = n47423 & n17168;
  assign n47449 = ~n47466;
  assign n47452 = ~n47423;
  assign n47360 = n47467 ^ n47468;
  assign n47481 = ~n47490;
  assign n47339 = ~n47365;
  assign n47338 = n47366 ^ n47367;
  assign n47356 = n47382 ^ n47383;
  assign n47363 = ~n47387;
  assign n47385 = ~n47382;
  assign n43453 = ~n43438;
  assign n47395 = n47344 & n45090;
  assign n47392 = ~n47413;
  assign n47394 = ~n47344;
  assign n47422 = n47449 & n47450;
  assign n47425 = ~n47451;
  assign n47439 = n47452 & n474;
  assign n47453 = n47481 & n47482;
  assign n46932 = n47338 ^ n45676;
  assign n47291 = n47355 ^ n47356;
  assign n47341 = ~n47338;
  assign n47342 = n47363 & n47364;
  assign n47368 = n47384 & n47385;
  assign n47369 = n43453 & n46182;
  assign n47370 = n43453 & n45179;
  assign n47371 = n47392 & n47393;
  assign n47388 = n47394 & n45088;
  assign n47347 = ~n47395;
  assign n47396 = n47422 ^ n47423;
  assign n47424 = ~n47422;
  assign n47398 = ~n47439;
  assign n47427 = n47453 ^ n47454;
  assign n47456 = n47453 & n47462;
  assign n47455 = ~n47453;
  assign n47329 = n47291 & n100;
  assign n45646 = ~n46932;
  assign n47328 = ~n47291;
  assign n47296 = n47341 & n45706;
  assign n47317 = n47342 ^ n47343;
  assign n47340 = ~n47342;
  assign n47357 = ~n47368;
  assign n47353 = ~n47369;
  assign n46253 = ~n47370;
  assign n47345 = n47371 ^ n45088;
  assign n47372 = ~n47371;
  assign n47373 = ~n47388;
  assign n47375 = n474 ^ n47396;
  assign n47414 = n47424 & n47425;
  assign n47377 = n47426 ^ n47427;
  assign n47440 = n47455 & n47454;
  assign n47436 = ~n47456;
  assign n47297 = n101 ^ n47317;
  assign n47316 = n47328 & n14710;
  assign n47275 = ~n47329;
  assign n47335 = n47339 & n47340;
  assign n43407 = n47344 ^ n47345;
  assign n47331 = n47353 & n47354;
  assign n47330 = n47357 & n47358;
  assign n47361 = n47372 & n47373;
  assign n47300 = n47374 ^ n47375;
  assign n47326 = n47375 & n47374;
  assign n47400 = n47377 & n473;
  assign n47397 = ~n47414;
  assign n47399 = ~n47377;
  assign n47428 = n47436 & n47437;
  assign n47410 = ~n47440;
  assign n45609 = n47296 ^ n47297;
  assign n47244 = n47297 & n47296;
  assign n47298 = ~n47316;
  assign n47305 = n47330 ^ n47331;
  assign n47320 = n43407 & n46091;
  assign n47321 = n43407 & n45088;
  assign n47318 = ~n47335;
  assign n47333 = n47331 & n47336;
  assign n43441 = ~n43407;
  assign n47313 = ~n47330;
  assign n47332 = ~n47331;
  assign n47349 = n47300 & n44966;
  assign n47346 = ~n47361;
  assign n47348 = ~n47300;
  assign n47334 = ~n47326;
  assign n47376 = n47397 & n47398;
  assign n47389 = n47399 & n17141;
  assign n47352 = ~n47400;
  assign n47409 = ~n47428;
  assign n46894 = ~n45609;
  assign n47255 = ~n47244;
  assign n47257 = n47305 ^ n47306;
  assign n47312 = n47318 & n47319;
  assign n47307 = ~n47320;
  assign n46144 = ~n47321;
  assign n47322 = n47332 & n47306;
  assign n47314 = ~n47333;
  assign n47323 = n47346 & n47347;
  assign n47337 = n47348 & n44980;
  assign n47302 = ~n47349;
  assign n47350 = n47376 ^ n47377;
  assign n47378 = ~n47376;
  assign n47379 = ~n47389;
  assign n47386 = n47409 & n47410;
  assign n47284 = n47257 & n99;
  assign n47283 = ~n47257;
  assign n47272 = n47307 & n47308;
  assign n47290 = ~n47312;
  assign n47309 = n47313 & n47314;
  assign n47294 = ~n47322;
  assign n47299 = n47323 ^ n44980;
  assign n47324 = ~n47323;
  assign n47325 = ~n47337;
  assign n47327 = n473 ^ n47350;
  assign n47362 = n47378 & n47379;
  assign n47359 = n472 ^ n47386;
  assign n47276 = n47283 & n14678;
  assign n47239 = ~n47284;
  assign n47268 = n47290 ^ n47291;
  assign n47286 = n47272 & n47292;
  assign n47289 = n47298 & n47290;
  assign n47285 = ~n47272;
  assign n43374 = n47299 ^ n47300;
  assign n47293 = ~n47309;
  assign n47315 = n47324 & n47325;
  assign n47258 = n47326 ^ n47327;
  assign n47311 = n47327 & n47334;
  assign n47288 = n47359 ^ n47360;
  assign n47351 = ~n47362;
  assign n47245 = n100 ^ n47268;
  assign n47253 = ~n47276;
  assign n47277 = n47285 & n47248;
  assign n47278 = n43374 & n45997;
  assign n47270 = ~n47286;
  assign n47279 = n43374 & n44980;
  assign n47274 = ~n47289;
  assign n47271 = n47293 & n47294;
  assign n43380 = ~n43374;
  assign n47303 = n47258 & n44862;
  assign n47301 = ~n47315;
  assign n47304 = ~n47258;
  assign n47310 = n47351 & n47352;
  assign n45593 = n47244 ^ n47245;
  assign n47216 = n47245 & n47255;
  assign n47247 = n47271 ^ n47272;
  assign n47256 = n47274 & n47275;
  assign n47250 = ~n47277;
  assign n47264 = ~n47278;
  assign n46067 = ~n47279;
  assign n47269 = ~n47271;
  assign n47280 = n47301 & n47302;
  assign n47262 = ~n47303;
  assign n47295 = n47304 & n44902;
  assign n47287 = n47310 ^ n47311;
  assign n46857 = ~n45593;
  assign n47220 = n47247 ^ n47248;
  assign n47237 = n47256 ^ n47257;
  assign n47210 = n47264 & n47265;
  assign n47254 = ~n47256;
  assign n47263 = n47269 & n47270;
  assign n47259 = n47280 ^ n44862;
  assign n47214 = n47287 ^ n47288;
  assign n47282 = ~n47280;
  assign n47281 = ~n47295;
  assign n47217 = n99 ^ n47237;
  assign n47230 = n47220 & n98;
  assign n47229 = ~n47220;
  assign n47243 = n47210 & n47251;
  assign n47246 = n47253 & n47254;
  assign n47242 = ~n47210;
  assign n43321 = n47258 ^ n47259;
  assign n47249 = ~n47263;
  assign n47266 = n47214 & n44822;
  assign n47267 = ~n47214;
  assign n47273 = n47281 & n47282;
  assign n45526 = n47216 ^ n47217;
  assign n47218 = ~n47217;
  assign n47225 = n47229 & n14640;
  assign n47191 = ~n47230;
  assign n47240 = n47242 & n47232;
  assign n47228 = ~n47243;
  assign n47238 = ~n47246;
  assign n47231 = n47249 & n47250;
  assign n43343 = ~n43321;
  assign n47224 = ~n47266;
  assign n47260 = n47267 & n44778;
  assign n47261 = ~n47273;
  assign n46814 = ~n45526;
  assign n47176 = n47218 & n47216;
  assign n47208 = ~n47225;
  assign n47211 = n47231 ^ n47232;
  assign n47219 = n47238 & n47239;
  assign n47213 = ~n47240;
  assign n47233 = n43343 & n45936;
  assign n47234 = n43343 & n44902;
  assign n47227 = ~n47231;
  assign n47241 = ~n47260;
  assign n47252 = n47261 & n47262;
  assign n47169 = n47210 ^ n47211;
  assign n47200 = n47219 ^ n47220;
  assign n47226 = n47227 & n47228;
  assign n47209 = ~n47219;
  assign n47221 = ~n47233;
  assign n45991 = ~n47234;
  assign n47236 = ~n47252;
  assign n47177 = n98 ^ n47200;
  assign n47193 = n47169 & n97;
  assign n47192 = ~n47169;
  assign n47207 = n47208 & n47209;
  assign n47174 = n47221 & n47222;
  assign n47212 = ~n47226;
  assign n47215 = n47236 ^ n44822;
  assign n47235 = n47236 & n47241;
  assign n45496 = n47176 ^ n47177;
  assign n47178 = ~n47177;
  assign n47186 = n47192 & n14600;
  assign n47155 = ~n47193;
  assign n47190 = ~n47207;
  assign n47203 = n47174 & n47195;
  assign n47194 = n47212 & n47213;
  assign n47201 = ~n47174;
  assign n43281 = n47214 ^ n47215;
  assign n47223 = ~n47235;
  assign n46773 = ~n45496;
  assign n47125 = n47178 & n47176;
  assign n47173 = ~n47186;
  assign n47187 = n47190 & n47191;
  assign n47175 = n47194 ^ n47195;
  assign n47196 = n47201 & n47202;
  assign n47189 = ~n47203;
  assign n47197 = n43281 & n45883;
  assign n47198 = n43281 & n44778;
  assign n47188 = ~n47194;
  assign n43312 = ~n43281;
  assign n47204 = n47223 & n47224;
  assign n47137 = n47174 ^ n47175;
  assign n47168 = ~n47187;
  assign n47181 = n47188 & n47189;
  assign n47171 = ~n47196;
  assign n47182 = ~n47197;
  assign n45931 = ~n47198;
  assign n47179 = n47204 ^ n44747;
  assign n47205 = ~n47204;
  assign n47156 = n47137 & n14563;
  assign n47145 = n47168 ^ n47169;
  assign n47157 = ~n47137;
  assign n47167 = n47168 & n47173;
  assign n43241 = n47179 ^ n47180;
  assign n47170 = ~n47181;
  assign n47128 = n47182 & n47183;
  assign n47199 = n47205 & n47206;
  assign n47126 = n97 ^ n47145;
  assign n47139 = ~n47156;
  assign n47146 = n47157 & n96;
  assign n47163 = n47128 & n47166;
  assign n47154 = ~n47167;
  assign n47161 = n43241 & n45842;
  assign n47162 = n43241 & n44747;
  assign n47149 = n47170 & n47171;
  assign n43276 = ~n43241;
  assign n47160 = ~n47128;
  assign n47184 = ~n47199;
  assign n45415 = n47125 ^ n47126;
  assign n47099 = n47126 & n47125;
  assign n47120 = ~n47146;
  assign n47129 = n47149 ^ n47150;
  assign n47136 = n47154 & n47155;
  assign n47158 = n47160 & n47150;
  assign n47147 = ~n47161;
  assign n45870 = ~n47162;
  assign n47152 = ~n47149;
  assign n47151 = ~n47163;
  assign n47172 = n47184 & n47185;
  assign n46725 = ~n45415;
  assign n47102 = ~n47099;
  assign n47104 = n47128 ^ n47129;
  assign n47118 = n47136 ^ n47137;
  assign n47138 = ~n47136;
  assign n47087 = n47147 & n47148;
  assign n47142 = n47151 & n47152;
  assign n47133 = ~n47158;
  assign n47165 = n47172 & n44611;
  assign n47164 = ~n47172;
  assign n47100 = n96 ^ n47118;
  assign n47113 = n47104 & n111;
  assign n47112 = ~n47104;
  assign n47127 = n47138 & n47139;
  assign n47131 = n47087 & n47140;
  assign n47130 = ~n47087;
  assign n47132 = ~n47142;
  assign n47159 = n47164 & n44651;
  assign n47144 = ~n47165;
  assign n46689 = n47099 ^ n47100;
  assign n47101 = ~n47100;
  assign n47107 = n47112 & n14517;
  assign n47079 = ~n47113;
  assign n47119 = ~n47127;
  assign n47123 = n47130 & n47110;
  assign n47114 = ~n47131;
  assign n47124 = n47132 & n47133;
  assign n47143 = n47144 & n47153;
  assign n47135 = ~n47159;
  assign n45346 = ~n46689;
  assign n47066 = n47101 & n47102;
  assign n47092 = ~n47107;
  assign n47103 = n47119 & n47120;
  assign n47094 = ~n47123;
  assign n47109 = ~n47124;
  assign n47134 = ~n47143;
  assign n47141 = n47135 & n47144;
  assign n47085 = n47103 ^ n47104;
  assign n47088 = n47109 ^ n47110;
  assign n47091 = ~n47103;
  assign n47108 = n47109 & n47114;
  assign n47115 = n47134 & n47135;
  assign n47121 = ~n47141;
  assign n47067 = n111 ^ n47085;
  assign n47053 = n47087 ^ n47088;
  assign n47086 = n47091 & n47092;
  assign n47093 = ~n47108;
  assign n47095 = n47115 ^ n44523;
  assign n43201 = n47121 ^ n47122;
  assign n47116 = ~n47115;
  assign n45275 = n47066 ^ n47067;
  assign n47018 = n47067 & n47066;
  assign n47070 = n47053 & n14497;
  assign n47071 = ~n47053;
  assign n47078 = ~n47086;
  assign n47080 = n47093 & n47094;
  assign n43165 = n47095 ^ n47096;
  assign n47105 = n43201 & n45809;
  assign n47106 = n43201 & n44611;
  assign n47111 = n47116 & n47117;
  assign n43234 = ~n43201;
  assign n46649 = ~n45275;
  assign n47028 = ~n47018;
  assign n47056 = ~n47070;
  assign n47068 = n47071 & n110;
  assign n47052 = n47078 & n47079;
  assign n47055 = n47080 ^ n47075;
  assign n47063 = ~n47080;
  assign n43187 = ~n43165;
  assign n47089 = ~n47105;
  assign n45829 = ~n47106;
  assign n47097 = ~n47111;
  assign n47035 = n47052 ^ n47053;
  assign n47039 = ~n47068;
  assign n47057 = ~n47052;
  assign n47072 = n43187 & n45748;
  assign n47073 = n43187 & n44523;
  assign n47054 = n47089 & n47090;
  assign n47082 = n47097 & n47098;
  assign n47019 = n110 ^ n47035;
  assign n47014 = n47054 ^ n47055;
  assign n47050 = n47056 & n47057;
  assign n47058 = ~n47072;
  assign n45783 = ~n47073;
  assign n47076 = n47054 & n47081;
  assign n47061 = n47082 ^ n44455;
  assign n47074 = ~n47054;
  assign n47083 = ~n47082;
  assign n45202 = n47018 ^ n47019;
  assign n46978 = n47019 & n47028;
  assign n47037 = n47014 & n109;
  assign n47036 = ~n47014;
  assign n47038 = ~n47050;
  assign n47002 = n47058 & n47059;
  assign n43124 = n47060 ^ n47061;
  assign n47069 = n47074 & n47075;
  assign n47062 = ~n47076;
  assign n47077 = n47083 & n47084;
  assign n46596 = ~n45202;
  assign n46977 = ~n46978;
  assign n47031 = n47036 & n14444;
  assign n47001 = ~n47037;
  assign n47032 = n47038 & n47039;
  assign n47041 = n47002 & n47049;
  assign n47042 = n43124 & n45723;
  assign n47043 = n43124 & n44455;
  assign n47040 = ~n47002;
  assign n43156 = ~n43124;
  assign n47051 = n47062 & n47063;
  assign n47045 = ~n47069;
  assign n47064 = ~n47077;
  assign n47017 = ~n47031;
  assign n47013 = ~n47032;
  assign n47033 = n47040 & n47025;
  assign n47020 = ~n47041;
  assign n47029 = ~n47042;
  assign n45743 = ~n47043;
  assign n47044 = ~n47051;
  assign n47046 = n47064 & n47065;
  assign n46996 = n47013 ^ n47014;
  assign n47012 = n47013 & n47017;
  assign n46964 = n47029 & n47030;
  assign n47005 = ~n47033;
  assign n47024 = n47044 & n47045;
  assign n47023 = n47046 ^ n44387;
  assign n47047 = ~n47046;
  assign n46979 = n109 ^ n46996;
  assign n47000 = ~n47012;
  assign n47011 = n46964 & n47015;
  assign n47010 = ~n46964;
  assign n43081 = n47022 ^ n47023;
  assign n47003 = n47024 ^ n47025;
  assign n47021 = ~n47024;
  assign n47034 = n47047 & n47048;
  assign n45119 = n46978 ^ n46979;
  assign n46976 = ~n46979;
  assign n46982 = n47000 & n47001;
  assign n46983 = n47002 ^ n47003;
  assign n47006 = n47010 & n46987;
  assign n46988 = ~n47011;
  assign n43113 = ~n43081;
  assign n47016 = n47020 & n47021;
  assign n47026 = ~n47034;
  assign n46552 = ~n45119;
  assign n46942 = n46976 & n46977;
  assign n46963 = n46982 ^ n46983;
  assign n46985 = n46983 & n108;
  assign n46962 = ~n46982;
  assign n46984 = ~n46983;
  assign n46967 = ~n47006;
  assign n46997 = n43113 & n45672;
  assign n46998 = n43113 & n44387;
  assign n47004 = ~n47016;
  assign n47007 = n47026 & n47027;
  assign n46943 = n108 ^ n46963;
  assign n46980 = n46984 & n14397;
  assign n46947 = ~n46985;
  assign n46990 = ~n46997;
  assign n45705 = ~n46998;
  assign n46986 = n47004 & n47005;
  assign n46992 = n47007 ^ n44362;
  assign n47008 = ~n47007;
  assign n45083 = n46942 ^ n46943;
  assign n46880 = n46943 & n46942;
  assign n46961 = ~n46980;
  assign n46965 = n46986 ^ n46987;
  assign n46923 = n46990 & n46991;
  assign n43038 = n46992 ^ n46993;
  assign n46989 = ~n46986;
  assign n46999 = n47008 & n47009;
  assign n46495 = ~n45083;
  assign n46883 = ~n46880;
  assign n46958 = n46961 & n46962;
  assign n46926 = n46964 ^ n46965;
  assign n46970 = n43038 & n45629;
  assign n46971 = n46923 & n46949;
  assign n46972 = n43038 & n44362;
  assign n46968 = ~n46923;
  assign n43072 = ~n43038;
  assign n46981 = n46988 & n46989;
  assign n46994 = ~n46999;
  assign n46945 = n46926 & n107;
  assign n46944 = ~n46926;
  assign n46946 = ~n46958;
  assign n46959 = n46968 & n46969;
  assign n46956 = ~n46970;
  assign n46950 = ~n46971;
  assign n45645 = ~n46972;
  assign n46966 = ~n46981;
  assign n46973 = n46994 & n46995;
  assign n46940 = n46944 & n14377;
  assign n46905 = ~n46945;
  assign n46925 = n46946 & n46947;
  assign n46888 = n46956 & n46957;
  assign n46928 = ~n46959;
  assign n46948 = n46966 & n46967;
  assign n46952 = n46973 ^ n44302;
  assign n46974 = ~n46973;
  assign n46903 = n46925 ^ n46926;
  assign n46921 = ~n46940;
  assign n46922 = ~n46925;
  assign n46939 = n46888 & n46909;
  assign n46924 = n46948 ^ n46949;
  assign n46937 = ~n46888;
  assign n43024 = n46952 ^ n46953;
  assign n46951 = ~n46948;
  assign n46960 = n46974 & n46975;
  assign n46881 = n107 ^ n46903;
  assign n46918 = n46921 & n46922;
  assign n46885 = n46923 ^ n46924;
  assign n46929 = n46937 & n46938;
  assign n46930 = n43024 & n45646;
  assign n46931 = n43024 & n45563;
  assign n46910 = ~n46939;
  assign n46933 = n43024 & n44302;
  assign n42998 = ~n43024;
  assign n46941 = n46950 & n46951;
  assign n46954 = ~n46960;
  assign n44960 = n46880 ^ n46881;
  assign n46882 = ~n46881;
  assign n46906 = n46885 & n14316;
  assign n46904 = ~n46918;
  assign n46907 = ~n46885;
  assign n46891 = ~n46929;
  assign n45649 = ~n46930;
  assign n46916 = ~n46931;
  assign n46919 = n42998 & n46932;
  assign n45608 = ~n46933;
  assign n46927 = ~n46941;
  assign n46934 = n46954 & n46955;
  assign n46437 = ~n44960;
  assign n46838 = n46882 & n46883;
  assign n46884 = n46904 & n46905;
  assign n46886 = ~n46906;
  assign n46900 = n46907 & n106;
  assign n46844 = n46916 & n46917;
  assign n45667 = ~n46919;
  assign n46908 = n46927 & n46928;
  assign n46913 = n46934 ^ n44202;
  assign n46935 = ~n46934;
  assign n46860 = n46884 ^ n46885;
  assign n46887 = ~n46884;
  assign n46862 = ~n46900;
  assign n46899 = n46844 & n46901;
  assign n46889 = n46908 ^ n46909;
  assign n46898 = ~n46844;
  assign n42966 = n46912 ^ n46913;
  assign n46911 = ~n46908;
  assign n46920 = n46935 & n46936;
  assign n46839 = n106 ^ n46860;
  assign n46875 = n46886 & n46887;
  assign n46841 = n46888 ^ n46889;
  assign n46892 = n46898 & n46866;
  assign n46893 = n42966 & n45609;
  assign n46869 = ~n46899;
  assign n42959 = ~n42966;
  assign n46902 = n46910 & n46911;
  assign n46914 = ~n46920;
  assign n44877 = n46838 ^ n46839;
  assign n46797 = n46839 & n46838;
  assign n46863 = n46841 & n14279;
  assign n46861 = ~n46875;
  assign n46864 = ~n46841;
  assign n46847 = ~n46892;
  assign n45636 = ~n46893;
  assign n46876 = n42959 & n45547;
  assign n46877 = n42959 & n46894;
  assign n46878 = n42959 & n44253;
  assign n46890 = ~n46902;
  assign n46895 = n46914 & n46915;
  assign n46366 = ~n44877;
  assign n46840 = n46861 & n46862;
  assign n46843 = ~n46863;
  assign n46858 = n46864 & n105;
  assign n46867 = ~n46876;
  assign n45614 = ~n46877;
  assign n45567 = ~n46878;
  assign n46865 = n46890 & n46891;
  assign n46871 = n46895 ^ n44191;
  assign n46896 = ~n46895;
  assign n46820 = n46840 ^ n46841;
  assign n46842 = ~n46840;
  assign n46819 = ~n46858;
  assign n46845 = n46865 ^ n46866;
  assign n46824 = n46867 & n46868;
  assign n42883 = n46871 ^ n46872;
  assign n46870 = ~n46865;
  assign n46879 = n46896 & n46897;
  assign n46798 = n105 ^ n46820;
  assign n46834 = n46842 & n46843;
  assign n46831 = n46844 ^ n46845;
  assign n46850 = n42883 & n45503;
  assign n46851 = n46824 & n46802;
  assign n46852 = n42883 & n46857;
  assign n46853 = n42883 & n44191;
  assign n46848 = ~n46824;
  assign n42952 = ~n42883;
  assign n46859 = n46869 & n46870;
  assign n46873 = ~n46879;
  assign n44793 = n46797 ^ n46798;
  assign n46753 = n46798 & n46797;
  assign n46822 = n46831 & n104;
  assign n46818 = ~n46834;
  assign n46821 = ~n46831;
  assign n46835 = n46848 & n46849;
  assign n46832 = ~n46850;
  assign n46826 = ~n46851;
  assign n45572 = ~n46852;
  assign n46836 = n42952 & n45593;
  assign n45533 = ~n46853;
  assign n46846 = ~n46859;
  assign n46854 = n46873 & n46874;
  assign n46287 = ~n44793;
  assign n46775 = n46818 & n46819;
  assign n46816 = n46821 & n14245;
  assign n46780 = ~n46822;
  assign n46760 = n46832 & n46833;
  assign n46804 = ~n46835;
  assign n45595 = ~n46836;
  assign n46823 = n46846 & n46847;
  assign n46827 = n46854 ^ n44172;
  assign n46855 = ~n46854;
  assign n46799 = ~n46775;
  assign n46800 = ~n46816;
  assign n46815 = n46760 & n46784;
  assign n46801 = n46823 ^ n46824;
  assign n46812 = ~n46760;
  assign n42867 = n46827 ^ n46828;
  assign n46825 = ~n46823;
  assign n46837 = n46855 & n46856;
  assign n46793 = n46799 & n46800;
  assign n46794 = n46800 & n46780;
  assign n46737 = n46801 ^ n46802;
  assign n46805 = n46812 & n46813;
  assign n46806 = n42867 & n46814;
  assign n46807 = n42867 & n45443;
  assign n46786 = ~n46815;
  assign n46808 = n42867 & n44172;
  assign n42913 = ~n42867;
  assign n46817 = n46825 & n46826;
  assign n46829 = ~n46837;
  assign n46781 = n46737 & n14200;
  assign n46779 = ~n46793;
  assign n46776 = ~n46794;
  assign n46782 = ~n46737;
  assign n46763 = ~n46805;
  assign n45528 = ~n46806;
  assign n46791 = ~n46807;
  assign n46795 = n42913 & n45526;
  assign n45467 = ~n46808;
  assign n46803 = ~n46817;
  assign n46809 = n46829 & n46830;
  assign n46754 = n46775 ^ n46776;
  assign n46757 = n46779 & n46780;
  assign n46759 = ~n46781;
  assign n46777 = n46782 & n119;
  assign n46743 = n46791 & n46792;
  assign n45552 = ~n46795;
  assign n46783 = n46803 & n46804;
  assign n46788 = n46809 ^ n44096;
  assign n46810 = ~n46809;
  assign n44713 = n46753 ^ n46754;
  assign n46711 = n46754 & n46753;
  assign n46736 = n119 ^ n46757;
  assign n46758 = ~n46757;
  assign n46739 = ~n46777;
  assign n46774 = n46743 & n46720;
  assign n46761 = n46783 ^ n46784;
  assign n46771 = ~n46743;
  assign n42827 = n46787 ^ n46788;
  assign n46785 = ~n46783;
  assign n46796 = n46810 & n46811;
  assign n46712 = n46736 ^ n46737;
  assign n46205 = ~n44713;
  assign n46714 = ~n46711;
  assign n46752 = n46758 & n46759;
  assign n46716 = n46760 ^ n46761;
  assign n46764 = n46771 & n46772;
  assign n46765 = n42827 & n46773;
  assign n46766 = n42827 & n45391;
  assign n46745 = ~n46774;
  assign n46767 = n42827 & n44115;
  assign n42873 = ~n42827;
  assign n46778 = n46785 & n46786;
  assign n46789 = ~n46796;
  assign n44625 = n46711 ^ n46712;
  assign n46713 = ~n46712;
  assign n46740 = n46716 & n14171;
  assign n46738 = ~n46752;
  assign n46741 = ~n46716;
  assign n46722 = ~n46764;
  assign n45473 = ~n46765;
  assign n46755 = n42873 & n45496;
  assign n46750 = ~n46766;
  assign n45422 = ~n46767;
  assign n46762 = ~n46778;
  assign n46768 = n46789 & n46790;
  assign n46140 = ~n44625;
  assign n46046 = n46713 & n46714;
  assign n46715 = n46738 & n46739;
  assign n46718 = ~n46740;
  assign n46733 = n46741 & n118;
  assign n46677 = n46750 & n46751;
  assign n45498 = ~n46755;
  assign n46742 = n46762 & n46763;
  assign n46747 = n46768 ^ n44061;
  assign n46769 = ~n46768;
  assign n46686 = ~n46046;
  assign n46695 = n46715 ^ n46716;
  assign n46717 = ~n46715;
  assign n46694 = ~n46733;
  assign n46732 = n46677 & n46734;
  assign n46719 = n46742 ^ n46743;
  assign n46731 = ~n46677;
  assign n42788 = n46746 ^ n46747;
  assign n46744 = ~n46742;
  assign n46756 = n46769 & n46770;
  assign n46009 = n118 ^ n46695;
  assign n46708 = n46717 & n46718;
  assign n46654 = n46719 ^ n46720;
  assign n46723 = n46731 & n46699;
  assign n46724 = n42788 & n45272;
  assign n46701 = ~n46732;
  assign n46726 = n42788 & n45415;
  assign n46727 = n42788 & n44061;
  assign n42832 = ~n42788;
  assign n46735 = n46744 & n46745;
  assign n46748 = ~n46756;
  assign n46629 = n46009 & n46686;
  assign n46696 = n46654 & n14111;
  assign n46693 = ~n46708;
  assign n46697 = ~n46654;
  assign n46680 = ~n46723;
  assign n46706 = ~n46724;
  assign n46709 = n42832 & n46725;
  assign n45417 = ~n46726;
  assign n45357 = ~n46727;
  assign n46721 = ~n46735;
  assign n46728 = n46748 & n46749;
  assign n46632 = ~n46629;
  assign n46674 = n46693 & n46694;
  assign n46676 = ~n46696;
  assign n46691 = n46697 & n117;
  assign n46637 = n46706 & n46707;
  assign n45448 = ~n46709;
  assign n46698 = n46721 & n46722;
  assign n46702 = n46728 ^ n44028;
  assign n46729 = ~n46728;
  assign n46653 = n117 ^ n46674;
  assign n46675 = ~n46674;
  assign n46656 = ~n46691;
  assign n46690 = n46637 & n46660;
  assign n46678 = n46698 ^ n46699;
  assign n46687 = ~n46637;
  assign n42744 = n46702 ^ n46703;
  assign n46700 = ~n46698;
  assign n46710 = n46729 & n46730;
  assign n46630 = n46653 ^ n46654;
  assign n46669 = n46675 & n46676;
  assign n46634 = n46677 ^ n46678;
  assign n46681 = n46687 & n46688;
  assign n46682 = n42744 & n46689;
  assign n46663 = ~n46690;
  assign n42777 = ~n42744;
  assign n46692 = n46700 & n46701;
  assign n46704 = ~n46710;
  assign n46609 = n46629 ^ n46630;
  assign n46631 = ~n46630;
  assign n46658 = n46634 & n116;
  assign n46655 = ~n46669;
  assign n46657 = ~n46634;
  assign n46640 = ~n46681;
  assign n45384 = ~n46682;
  assign n46670 = n42777 & n45157;
  assign n46671 = n42777 & n45346;
  assign n46672 = n42777 & n44028;
  assign n46679 = ~n46692;
  assign n46683 = n46704 & n46705;
  assign n42460 = n46609 ^ n43600;
  assign n46610 = ~n46609;
  assign n46585 = n46631 & n46632;
  assign n46633 = n46655 & n46656;
  assign n46651 = n46657 & n14072;
  assign n46613 = ~n46658;
  assign n46661 = ~n46670;
  assign n45349 = ~n46671;
  assign n45285 = ~n46672;
  assign n46659 = n46679 & n46680;
  assign n46665 = n46683 ^ n43989;
  assign n46684 = ~n46683;
  assign n46584 = n42460 & n45539;
  assign n42462 = ~n42460;
  assign n46501 = n46610 & n43602;
  assign n46604 = n46610 & n43600;
  assign n46583 = ~n46585;
  assign n46611 = n46633 ^ n46634;
  assign n46635 = ~n46633;
  assign n46636 = ~n46651;
  assign n46638 = n46659 ^ n46660;
  assign n46591 = n46661 & n46662;
  assign n42748 = n46665 ^ n46666;
  assign n46664 = ~n46659;
  assign n46673 = n46684 & n46685;
  assign n46574 = ~n46584;
  assign n45558 = ~n46604;
  assign n46586 = n116 ^ n46611;
  assign n46625 = n46635 & n46636;
  assign n46588 = n46637 ^ n46638;
  assign n46642 = n42748 & n46649;
  assign n46643 = n46591 & n46650;
  assign n46644 = n42748 & n45174;
  assign n46645 = n42748 & n43989;
  assign n46641 = ~n46591;
  assign n42706 = ~n42748;
  assign n46652 = n46663 & n46664;
  assign n46667 = ~n46673;
  assign n46548 = n46574 & n46575;
  assign n46576 = n46585 ^ n46586;
  assign n46582 = ~n46586;
  assign n46608 = n46588 & n14061;
  assign n46612 = ~n46625;
  assign n46614 = ~n46588;
  assign n46626 = n46641 & n46616;
  assign n45278 = ~n46642;
  assign n46618 = ~n46643;
  assign n46623 = ~n46644;
  assign n46627 = n42706 & n45275;
  assign n45212 = ~n46645;
  assign n46639 = ~n46652;
  assign n46646 = n46667 & n46668;
  assign n46519 = n46548 ^ n46549;
  assign n46550 = ~n46548;
  assign n46558 = n46576 & n43547;
  assign n46557 = ~n46576;
  assign n46530 = n46582 & n46583;
  assign n46590 = ~n46608;
  assign n46587 = n46612 & n46613;
  assign n46605 = n46614 & n115;
  assign n46536 = n46623 & n46624;
  assign n46594 = ~n46626;
  assign n45318 = ~n46627;
  assign n46615 = n46639 & n46640;
  assign n46619 = n46646 ^ n43944;
  assign n46647 = ~n46646;
  assign n44105 = n263 ^ n46519;
  assign n46251 = n46519 & n263;
  assign n46374 = n46550 & n46551;
  assign n46554 = n46557 & n43551;
  assign n46503 = ~n46558;
  assign n46533 = ~n46530;
  assign n46559 = n46587 ^ n46588;
  assign n46589 = ~n46587;
  assign n46561 = ~n46605;
  assign n46603 = n46536 & n46606;
  assign n46592 = n46615 ^ n46616;
  assign n46602 = ~n46536;
  assign n42660 = n46619 ^ n46620;
  assign n46617 = ~n46615;
  assign n46628 = n46647 & n46648;
  assign n44135 = ~n44105;
  assign n46529 = ~n46554;
  assign n46531 = n115 ^ n46559;
  assign n46577 = n46589 & n46590;
  assign n46535 = n46591 ^ n46592;
  assign n46595 = n46602 & n46565;
  assign n46569 = ~n46603;
  assign n46597 = n42660 & n45202;
  assign n42695 = ~n42660;
  assign n46607 = n46617 & n46618;
  assign n46621 = ~n46628;
  assign n46522 = n46529 & n46501;
  assign n46500 = n46529 & n46503;
  assign n46445 = n46530 ^ n46531;
  assign n46532 = ~n46531;
  assign n46563 = n46535 & n114;
  assign n46560 = ~n46577;
  assign n46562 = ~n46535;
  assign n46539 = ~n46595;
  assign n46578 = n42695 & n45040;
  assign n46579 = n42695 & n46596;
  assign n45245 = ~n46597;
  assign n46580 = n42695 & n43944;
  assign n46593 = ~n46607;
  assign n46598 = n46621 & n46622;
  assign n42355 = n46500 ^ n46501;
  assign n46505 = n46445 & n43510;
  assign n46502 = ~n46522;
  assign n46504 = ~n46445;
  assign n46475 = n46532 & n46533;
  assign n46534 = n46560 & n46561;
  assign n46555 = n46562 & n14006;
  assign n46508 = ~n46563;
  assign n46566 = ~n46578;
  assign n45205 = ~n46579;
  assign n45117 = ~n46580;
  assign n46564 = n46593 & n46594;
  assign n46570 = n46598 ^ n46599;
  assign n46600 = ~n46598;
  assign n46472 = n42355 & n45520;
  assign n46473 = n42355 & n43551;
  assign n42364 = ~n42355;
  assign n46474 = n46502 & n46503;
  assign n46496 = n46504 & n43521;
  assign n46470 = ~n46505;
  assign n46478 = ~n46475;
  assign n46506 = n46534 ^ n46535;
  assign n46527 = ~n46534;
  assign n46528 = ~n46555;
  assign n46537 = n46564 ^ n46565;
  assign n46483 = n46566 & n46567;
  assign n42595 = n43869 ^ n46570;
  assign n46571 = n46570 & n43929;
  assign n46568 = ~n46564;
  assign n46581 = n46600 & n46601;
  assign n46462 = ~n46472;
  assign n45458 = ~n46473;
  assign n46446 = n46474 ^ n43521;
  assign n46471 = ~n46474;
  assign n46448 = ~n46496;
  assign n46476 = n114 ^ n46506;
  assign n46523 = n46527 & n46528;
  assign n46480 = n46536 ^ n46537;
  assign n46541 = n42595 & n46552;
  assign n46542 = n42595 & n45000;
  assign n46543 = n46483 & n46553;
  assign n46540 = ~n46483;
  assign n42667 = ~n42595;
  assign n46556 = n46568 & n46569;
  assign n45042 = ~n46571;
  assign n46572 = ~n46581;
  assign n42287 = n46445 ^ n46446;
  assign n46438 = n46462 & n46463;
  assign n46466 = n46470 & n46471;
  assign n46381 = n46475 ^ n46476;
  assign n46477 = ~n46476;
  assign n46510 = n46480 & n113;
  assign n46507 = ~n46523;
  assign n46509 = ~n46480;
  assign n46524 = n46540 & n46512;
  assign n45121 = ~n46541;
  assign n46525 = n42667 & n45119;
  assign n46520 = ~n46542;
  assign n46514 = ~n46543;
  assign n46538 = ~n46556;
  assign n46544 = n46572 & n46573;
  assign n46409 = n42287 & n45367;
  assign n46410 = n42287 & n43510;
  assign n46430 = n46438 & n46439;
  assign n42305 = ~n42287;
  assign n46431 = ~n46438;
  assign n46450 = n46381 & n43481;
  assign n46447 = ~n46466;
  assign n46449 = ~n46381;
  assign n46415 = n46477 & n46478;
  assign n46479 = n46507 & n46508;
  assign n46497 = n46509 & n13964;
  assign n46444 = ~n46510;
  assign n46455 = n46520 & n46521;
  assign n46486 = ~n46524;
  assign n45165 = ~n46525;
  assign n46511 = n46538 & n46539;
  assign n46515 = n46544 ^ n46545;
  assign n46546 = ~n46544;
  assign n46399 = ~n46409;
  assign n45398 = ~n46410;
  assign n46402 = ~n46430;
  assign n46411 = n46431 & n46432;
  assign n46412 = n46447 & n46448;
  assign n46440 = n46449 & n43493;
  assign n46383 = ~n46450;
  assign n46433 = ~n46415;
  assign n46451 = n46479 ^ n46480;
  assign n46481 = ~n46479;
  assign n46482 = ~n46497;
  assign n46494 = n46455 & n46498;
  assign n46484 = n46511 ^ n46512;
  assign n46493 = ~n46455;
  assign n42622 = n46515 ^ n43846;
  assign n46516 = n46515 & n43852;
  assign n46513 = ~n46511;
  assign n46526 = n46546 & n46547;
  assign n46292 = n46399 & n46400;
  assign n46401 = n46402 & n46374;
  assign n46377 = ~n46411;
  assign n46380 = n46412 ^ n43493;
  assign n46413 = ~n46412;
  assign n46414 = ~n46440;
  assign n46416 = n113 ^ n46451;
  assign n46467 = n46481 & n46482;
  assign n46418 = n46483 ^ n46484;
  assign n46487 = n46493 & n46422;
  assign n46456 = ~n46494;
  assign n46488 = n42622 & n44851;
  assign n46489 = n42622 & n46495;
  assign n42555 = ~n42622;
  assign n46499 = n46513 & n46514;
  assign n44974 = ~n46516;
  assign n46517 = ~n46526;
  assign n46372 = n46292 & n46335;
  assign n46370 = ~n46292;
  assign n42228 = n46380 ^ n46381;
  assign n46376 = ~n46401;
  assign n46373 = n46377 & n46402;
  assign n46403 = n46413 & n46414;
  assign n46310 = n46415 ^ n46416;
  assign n46351 = n46416 & n46433;
  assign n46453 = n46418 & n112;
  assign n46443 = ~n46467;
  assign n46452 = ~n46418;
  assign n46424 = ~n46487;
  assign n46464 = ~n46488;
  assign n45048 = ~n46489;
  assign n46468 = n42555 & n45083;
  assign n46485 = ~n46499;
  assign n46490 = n46517 & n46518;
  assign n46345 = n46370 & n46371;
  assign n46346 = n42228 & n45282;
  assign n46338 = ~n46372;
  assign n46347 = n42228 & n43493;
  assign n46339 = n46373 ^ n46374;
  assign n46375 = n46376 & n46377;
  assign n42261 = ~n42228;
  assign n46382 = ~n46403;
  assign n46417 = n46443 & n46444;
  assign n46441 = n46452 & n13918;
  assign n46386 = ~n46453;
  assign n46390 = n46464 & n46465;
  assign n45085 = ~n46468;
  assign n46454 = n46485 & n46486;
  assign n46459 = n46490 ^ n43792;
  assign n46491 = ~n46490;
  assign n46333 = n46339 & n262;
  assign n46302 = ~n46345;
  assign n46329 = ~n46346;
  assign n45324 = ~n46347;
  assign n46332 = ~n46339;
  assign n46334 = ~n46375;
  assign n46348 = n46382 & n46383;
  assign n46384 = n46417 ^ n46418;
  assign n46420 = ~n46417;
  assign n46419 = ~n46441;
  assign n46436 = n46390 & n46357;
  assign n46421 = n46454 ^ n46455;
  assign n46434 = ~n46390;
  assign n42509 = n46458 ^ n46459;
  assign n46457 = ~n46454;
  assign n46469 = n46491 & n46492;
  assign n46220 = n46329 & n46330;
  assign n46309 = n46332 & n11627;
  assign n46255 = ~n46333;
  assign n46293 = n46334 ^ n46335;
  assign n46331 = n46338 & n46334;
  assign n46311 = n46348 ^ n43438;
  assign n46350 = n46348 & n43438;
  assign n46349 = ~n46348;
  assign n46352 = n112 ^ n46384;
  assign n46404 = n46419 & n46420;
  assign n46315 = n46421 ^ n46422;
  assign n46425 = n46434 & n46435;
  assign n46393 = ~n46436;
  assign n46426 = n42509 & n46437;
  assign n42582 = ~n42509;
  assign n46442 = n46456 & n46457;
  assign n46460 = ~n46469;
  assign n46190 = n46292 ^ n46293;
  assign n46296 = n46220 & n46303;
  assign n46294 = ~n46220;
  assign n46295 = ~n46309;
  assign n42189 = n46310 ^ n46311;
  assign n46301 = ~n46331;
  assign n46340 = n46349 & n43453;
  assign n46328 = ~n46350;
  assign n46211 = n46351 ^ n46352;
  assign n46272 = n46352 & n46351;
  assign n46388 = n46315 & n127;
  assign n46385 = ~n46404;
  assign n46387 = ~n46315;
  assign n46359 = ~n46425;
  assign n46405 = n42582 & n44855;
  assign n46406 = n42582 & n43792;
  assign n46407 = n42582 & n44960;
  assign n45006 = ~n46426;
  assign n46423 = ~n46442;
  assign n46427 = n46460 & n46461;
  assign n46249 = n46190 & n261;
  assign n46248 = ~n46190;
  assign n46268 = n46294 & n46262;
  assign n46269 = n46295 & n46251;
  assign n46250 = n46295 & n46255;
  assign n46270 = n42189 & n45188;
  assign n46263 = ~n46296;
  assign n46271 = n42189 & n43438;
  assign n46261 = n46301 & n46302;
  assign n42216 = ~n42189;
  assign n46312 = n46328 & n46310;
  assign n46313 = n46211 & n43441;
  assign n46298 = ~n46340;
  assign n46308 = ~n46211;
  assign n46275 = ~n46272;
  assign n46353 = n46385 & n46386;
  assign n46378 = n46387 & n13893;
  assign n46317 = ~n46388;
  assign n46391 = ~n46405;
  assign n44893 = ~n46406;
  assign n44963 = ~n46407;
  assign n46389 = n46423 & n46424;
  assign n46396 = n46427 ^ n43789;
  assign n46428 = ~n46427;
  assign n46229 = n46248 & n11492;
  assign n46170 = ~n46249;
  assign n46210 = n46250 ^ n46251;
  assign n46221 = n46261 ^ n46262;
  assign n46223 = ~n46268;
  assign n46254 = ~n46269;
  assign n46252 = ~n46270;
  assign n45226 = ~n46271;
  assign n46264 = ~n46261;
  assign n46304 = n46308 & n43407;
  assign n46297 = ~n46312;
  assign n46258 = ~n46313;
  assign n46314 = n127 ^ n46353;
  assign n46355 = ~n46353;
  assign n46354 = ~n46378;
  assign n46356 = n46389 ^ n46390;
  assign n46280 = n46391 & n46392;
  assign n42489 = n46395 ^ n46396;
  assign n46394 = ~n46389;
  assign n46408 = n46428 & n46429;
  assign n44080 = n46210 ^ n44105;
  assign n46132 = n46220 ^ n46221;
  assign n46106 = n46210 & n44105;
  assign n46213 = ~n46229;
  assign n46141 = n46252 & n46253;
  assign n46230 = n46254 & n46255;
  assign n46247 = n46263 & n46264;
  assign n46256 = n46297 & n46298;
  assign n46217 = ~n46304;
  assign n46273 = n46314 ^ n46315;
  assign n46341 = n46354 & n46355;
  assign n46277 = n46356 ^ n46357;
  assign n46362 = n42489 & n44685;
  assign n46363 = n46280 & n46321;
  assign n46364 = n42489 & n44877;
  assign n46365 = n42489 & n43750;
  assign n46360 = ~n46280;
  assign n42536 = ~n42489;
  assign n46379 = n46393 & n46394;
  assign n46397 = ~n46408;
  assign n46180 = n46132 & n260;
  assign n45313 = ~n44080;
  assign n46179 = ~n46132;
  assign n46110 = ~n46106;
  assign n46215 = n46141 & n46224;
  assign n46214 = ~n46141;
  assign n46189 = ~n46230;
  assign n46222 = ~n46247;
  assign n46212 = n46256 ^ n43407;
  assign n46257 = ~n46256;
  assign n46135 = n46272 ^ n46273;
  assign n46274 = ~n46273;
  assign n46318 = n46277 & n13832;
  assign n46316 = ~n46341;
  assign n46319 = ~n46277;
  assign n46342 = n46360 & n46361;
  assign n46336 = ~n46362;
  assign n46323 = ~n46363;
  assign n44879 = ~n46364;
  assign n44811 = ~n46365;
  assign n46343 = n42536 & n46366;
  assign n46358 = ~n46379;
  assign n46367 = n46397 & n46398;
  assign n46168 = n46179 & n11437;
  assign n46089 = ~n46180;
  assign n46151 = n46189 ^ n46190;
  assign n42142 = n46211 ^ n46212;
  assign n46188 = n46213 & n46189;
  assign n46191 = n46214 & n46182;
  assign n46184 = ~n46215;
  assign n46181 = n46222 & n46223;
  assign n46231 = n46257 & n46258;
  assign n46233 = n46135 & n43374;
  assign n46232 = ~n46135;
  assign n46192 = n46274 & n46275;
  assign n46276 = n46316 & n46317;
  assign n46278 = ~n46318;
  assign n46305 = n46319 & n126;
  assign n46198 = n46336 & n46337;
  assign n46283 = ~n46342;
  assign n44924 = ~n46343;
  assign n46320 = n46358 & n46359;
  assign n46324 = n46367 ^ n43753;
  assign n46368 = ~n46367;
  assign n46107 = n261 ^ n46151;
  assign n46129 = ~n46168;
  assign n46142 = n46181 ^ n46182;
  assign n46172 = n42142 & n43441;
  assign n46173 = n42142 & n45090;
  assign n46169 = ~n46188;
  assign n46146 = ~n46191;
  assign n42167 = ~n42142;
  assign n46183 = ~n46181;
  assign n46216 = ~n46231;
  assign n46225 = n46232 & n43380;
  assign n46137 = ~n46233;
  assign n46234 = n46276 ^ n46277;
  assign n46279 = ~n46276;
  assign n46236 = ~n46305;
  assign n46300 = n46198 & n46306;
  assign n46281 = n46320 ^ n46321;
  assign n46299 = ~n46198;
  assign n42513 = n46324 ^ n46325;
  assign n46322 = ~n46320;
  assign n46344 = n46368 & n46369;
  assign n45241 = n46106 ^ n46107;
  assign n46053 = n46141 ^ n46142;
  assign n46109 = ~n46107;
  assign n46131 = n46169 & n46170;
  assign n45129 = ~n46172;
  assign n46143 = ~n46173;
  assign n46171 = n46183 & n46184;
  assign n46174 = n46216 & n46217;
  assign n46176 = ~n46225;
  assign n46193 = n126 ^ n46234;
  assign n46265 = n46278 & n46279;
  assign n46195 = n46280 ^ n46281;
  assign n46284 = n46299 & n46240;
  assign n46242 = ~n46300;
  assign n46285 = n42513 & n44668;
  assign n46286 = n42513 & n44793;
  assign n46288 = n42513 & n43753;
  assign n42439 = ~n42513;
  assign n46307 = n46322 & n46323;
  assign n46326 = ~n46344;
  assign n44040 = ~n45241;
  assign n46101 = n46053 & n259;
  assign n46050 = n46109 & n46110;
  assign n46100 = ~n46053;
  assign n46087 = n46131 ^ n46132;
  assign n46056 = n46143 & n46144;
  assign n46130 = ~n46131;
  assign n46145 = ~n46171;
  assign n46134 = n46174 ^ n43380;
  assign n46175 = ~n46174;
  assign n46058 = n46192 ^ n46193;
  assign n46112 = n46193 & n46192;
  assign n46237 = n46195 & n13776;
  assign n46235 = ~n46265;
  assign n46238 = ~n46195;
  assign n46201 = ~n46284;
  assign n46259 = ~n46285;
  assign n44796 = ~n46286;
  assign n46266 = n42439 & n46287;
  assign n44712 = ~n46288;
  assign n46282 = ~n46307;
  assign n46289 = n46326 & n46327;
  assign n46051 = n260 ^ n46087;
  assign n46090 = n46100 & n11347;
  assign n46017 = ~n46101;
  assign n46103 = n46056 & n46111;
  assign n46108 = n46129 & n46130;
  assign n46102 = ~n46056;
  assign n42097 = n46134 ^ n46135;
  assign n46133 = n46145 & n46146;
  assign n46152 = n46175 & n46176;
  assign n46154 = n46058 & n43343;
  assign n46153 = ~n46058;
  assign n46115 = ~n46112;
  assign n46194 = n46235 & n46236;
  assign n46196 = ~n46237;
  assign n46226 = n46238 & n125;
  assign n46120 = n46259 & n46260;
  assign n44841 = ~n46266;
  assign n46239 = n46282 & n46283;
  assign n46244 = n46289 ^ n43672;
  assign n46290 = ~n46289;
  assign n43998 = n46050 ^ n46051;
  assign n45978 = n46051 & n46050;
  assign n46054 = ~n46090;
  assign n46092 = n46102 & n46091;
  assign n46093 = n42097 & n44966;
  assign n46071 = ~n46103;
  assign n46094 = n42097 & n43380;
  assign n46088 = ~n46108;
  assign n42117 = ~n42097;
  assign n46072 = ~n46133;
  assign n46136 = ~n46152;
  assign n46147 = n46153 & n43321;
  assign n46061 = ~n46154;
  assign n46155 = n46194 ^ n46195;
  assign n46197 = ~n46194;
  assign n46157 = ~n46226;
  assign n46219 = n46120 & n46227;
  assign n46199 = n46239 ^ n46240;
  assign n46218 = ~n46120;
  assign n42386 = n46243 ^ n46244;
  assign n46241 = ~n46239;
  assign n46267 = n46290 & n46291;
  assign n45162 = ~n43998;
  assign n45977 = ~n45978;
  assign n46065 = n46071 & n46072;
  assign n46052 = n46088 & n46089;
  assign n46057 = n46072 ^ n46091;
  assign n46036 = ~n46092;
  assign n46066 = ~n46093;
  assign n45010 = ~n46094;
  assign n46095 = n46136 & n46137;
  assign n46097 = ~n46147;
  assign n46113 = n125 ^ n46155;
  assign n46185 = n46196 & n46197;
  assign n46117 = n46198 ^ n46199;
  assign n46202 = n46218 & n46161;
  assign n46203 = n42386 & n44513;
  assign n46163 = ~n46219;
  assign n46204 = n42386 & n43672;
  assign n46206 = n42386 & n44713;
  assign n42443 = ~n42386;
  assign n46228 = n46241 & n46242;
  assign n46245 = ~n46267;
  assign n46018 = n46052 ^ n46053;
  assign n45981 = n46056 ^ n46057;
  assign n46035 = ~n46065;
  assign n45960 = n46066 & n46067;
  assign n46055 = ~n46052;
  assign n46059 = n46095 ^ n43321;
  assign n46096 = ~n46095;
  assign n45984 = n46112 ^ n46113;
  assign n46114 = ~n46113;
  assign n46159 = n46117 & n124;
  assign n46156 = ~n46185;
  assign n46158 = ~n46117;
  assign n46123 = ~n46202;
  assign n46177 = ~n46203;
  assign n44624 = ~n46204;
  assign n46186 = n42443 & n46205;
  assign n44716 = ~n46206;
  assign n46200 = ~n46228;
  assign n46207 = n46245 & n46246;
  assign n45979 = n259 ^ n46018;
  assign n46019 = n45981 & n11226;
  assign n46020 = ~n45981;
  assign n45996 = n46035 & n46036;
  assign n46028 = n45960 & n46037;
  assign n46034 = n46054 & n46055;
  assign n46027 = ~n45960;
  assign n42062 = n46058 ^ n46059;
  assign n46073 = n46096 & n46097;
  assign n46075 = n45984 & n43312;
  assign n46074 = ~n45984;
  assign n46032 = n46114 & n46115;
  assign n46116 = n46156 & n46157;
  assign n46148 = n46158 & n13745;
  assign n46078 = ~n46159;
  assign n46044 = n46177 & n46178;
  assign n44758 = ~n46186;
  assign n46160 = n46200 & n46201;
  assign n46165 = n46207 ^ n43642;
  assign n46208 = ~n46207;
  assign n45081 = n45978 ^ n45979;
  assign n45976 = ~n45979;
  assign n45961 = n45996 ^ n45997;
  assign n45982 = ~n46019;
  assign n45995 = n46020 & n258;
  assign n45998 = ~n45996;
  assign n46021 = n46027 & n45997;
  assign n46022 = n42062 & n44862;
  assign n45999 = ~n46028;
  assign n46023 = n42062 & n43321;
  assign n46016 = ~n46034;
  assign n42075 = ~n42062;
  assign n46060 = ~n46073;
  assign n46068 = n46074 & n43281;
  assign n46025 = ~n46075;
  assign n46039 = ~n46032;
  assign n46076 = n46116 ^ n46117;
  assign n46119 = ~n46116;
  assign n46118 = ~n46148;
  assign n46139 = n46044 & n46149;
  assign n46121 = n46160 ^ n46161;
  assign n46138 = ~n46044;
  assign n42333 = n46164 ^ n46165;
  assign n46162 = ~n46160;
  assign n46187 = n46208 & n46209;
  assign n45096 = ~n45081;
  assign n45923 = n45960 ^ n45961;
  assign n45918 = n45976 & n45977;
  assign n45948 = ~n45995;
  assign n45989 = n45998 & n45999;
  assign n45980 = n46016 & n46017;
  assign n45959 = ~n46021;
  assign n45990 = ~n46022;
  assign n44927 = ~n46023;
  assign n46024 = n46060 & n46061;
  assign n45987 = ~n46068;
  assign n46033 = n124 ^ n46076;
  assign n46104 = n46118 & n46119;
  assign n46041 = n46120 ^ n46121;
  assign n46124 = n46138 & n46082;
  assign n46125 = n42333 & n44445;
  assign n46084 = ~n46139;
  assign n46126 = n42333 & n46140;
  assign n46127 = n42333 & n43648;
  assign n42393 = ~n42333;
  assign n46150 = n46162 & n46163;
  assign n46166 = ~n46187;
  assign n45934 = n45923 & n257;
  assign n45933 = ~n45923;
  assign n45921 = ~n45918;
  assign n45946 = n45980 ^ n45981;
  assign n45958 = ~n45989;
  assign n45905 = n45990 & n45991;
  assign n45983 = ~n45980;
  assign n45985 = n46024 ^ n43281;
  assign n45924 = n46032 ^ n46033;
  assign n46026 = ~n46024;
  assign n46038 = ~n46033;
  assign n46080 = n46041 & n123;
  assign n46077 = ~n46104;
  assign n46079 = ~n46041;
  assign n46048 = ~n46124;
  assign n46098 = ~n46125;
  assign n46105 = n42393 & n44625;
  assign n44690 = ~n46126;
  assign n44555 = ~n46127;
  assign n46122 = ~n46150;
  assign n46128 = n46166 & n46167;
  assign n45928 = n45933 & n11154;
  assign n45879 = ~n45934;
  assign n45919 = n258 ^ n45946;
  assign n45935 = n45958 & n45959;
  assign n45956 = n45905 & n45963;
  assign n45962 = n45982 & n45983;
  assign n45955 = ~n45905;
  assign n42018 = n45984 ^ n45985;
  assign n46000 = n46025 & n46026;
  assign n46002 = n45924 & n43241;
  assign n46001 = ~n45924;
  assign n45964 = n46038 & n46039;
  assign n46040 = n46077 & n46078;
  assign n46069 = n46079 & n13696;
  assign n46005 = ~n46080;
  assign n45970 = n46098 & n46099;
  assign n44643 = ~n46105;
  assign n46081 = n46122 & n46123;
  assign n46086 = n46128 ^ n43634;
  assign n43935 = n45918 ^ n45919;
  assign n45903 = ~n45928;
  assign n45920 = ~n45919;
  assign n45906 = n45935 ^ n45936;
  assign n45938 = ~n45935;
  assign n45949 = n45955 & n45936;
  assign n45937 = ~n45956;
  assign n45950 = n42018 & n44822;
  assign n45951 = n42018 & n43312;
  assign n45947 = ~n45962;
  assign n42040 = ~n42018;
  assign n45986 = ~n46000;
  assign n45992 = n46001 & n43276;
  assign n45927 = ~n46002;
  assign n45988 = ~n45964;
  assign n46003 = n46040 ^ n46041;
  assign n46042 = ~n46040;
  assign n46043 = ~n46069;
  assign n46064 = n45970 & n46011;
  assign n46045 = n46081 ^ n46082;
  assign n46062 = ~n45970;
  assign n42337 = n46085 ^ n46086;
  assign n46083 = ~n46081;
  assign n45017 = ~n43935;
  assign n45857 = n45905 ^ n45906;
  assign n45867 = n45920 & n45921;
  assign n45929 = n45937 & n45938;
  assign n45922 = n45947 & n45948;
  assign n45908 = ~n45949;
  assign n45930 = ~n45950;
  assign n44866 = ~n45951;
  assign n45952 = n45986 & n45987;
  assign n45954 = ~n45992;
  assign n45965 = n123 ^ n46003;
  assign n46029 = n46042 & n46043;
  assign n45967 = n46044 ^ n46045;
  assign n46008 = n46046 ^ n42337;
  assign n46049 = n46062 & n46063;
  assign n46013 = ~n46064;
  assign n44570 = ~n42337;
  assign n46070 = n46083 & n46084;
  assign n45881 = n45857 & n256;
  assign n45880 = ~n45857;
  assign n45893 = n45922 ^ n45923;
  assign n45907 = ~n45929;
  assign n45860 = n45930 & n45931;
  assign n45904 = ~n45922;
  assign n45925 = n45952 ^ n43241;
  assign n45953 = ~n45952;
  assign n45872 = n45964 ^ n45965;
  assign n45910 = n45965 & n45988;
  assign n44605 = n46008 ^ n46009;
  assign n46007 = n45967 & n122;
  assign n46004 = ~n46029;
  assign n46006 = ~n45967;
  assign n45975 = ~n46049;
  assign n46030 = n44570 & n44492;
  assign n46031 = n44570 & n43634;
  assign n46047 = ~n46070;
  assign n45874 = n45880 & n11085;
  assign n45838 = ~n45881;
  assign n45868 = n257 ^ n45893;
  assign n45899 = n45903 & n45904;
  assign n45882 = n45907 & n45908;
  assign n45901 = n45860 & n45909;
  assign n45900 = ~n45860;
  assign n41980 = n45924 ^ n45925;
  assign n45939 = n45953 & n45954;
  assign n45966 = n46004 & n46005;
  assign n45993 = n46006 & n13622;
  assign n45942 = ~n46007;
  assign n46014 = ~n46030;
  assign n44531 = ~n46031;
  assign n46010 = n46047 & n46048;
  assign n44919 = n45867 ^ n45868;
  assign n45815 = n45868 & n45867;
  assign n45859 = ~n45874;
  assign n45861 = n45882 ^ n45883;
  assign n45878 = ~n45899;
  assign n45884 = ~n45882;
  assign n45894 = n45900 & n45883;
  assign n45885 = ~n45901;
  assign n41991 = ~n41980;
  assign n45926 = ~n45939;
  assign n45940 = n45966 ^ n45967;
  assign n45968 = ~n45966;
  assign n45969 = ~n45993;
  assign n45971 = n46010 ^ n46011;
  assign n45972 = n46014 & n46015;
  assign n46012 = ~n46010;
  assign n43875 = ~n44919;
  assign n45818 = n45860 ^ n45861;
  assign n45856 = n45878 & n45879;
  assign n45875 = n45884 & n45885;
  assign n45863 = ~n45894;
  assign n45886 = n41991 & n44697;
  assign n45887 = n41991 & n43276;
  assign n45895 = n45926 & n45927;
  assign n45911 = n122 ^ n45940;
  assign n45957 = n45968 & n45969;
  assign n45913 = n45970 ^ n45971;
  assign n45917 = n45972 ^ n45973;
  assign n45994 = n46012 & n46013;
  assign n45840 = n45818 & n271;
  assign n45839 = ~n45818;
  assign n45836 = n45856 ^ n45857;
  assign n45858 = ~n45856;
  assign n45862 = ~n45875;
  assign n45869 = ~n45886;
  assign n44782 = ~n45887;
  assign n45871 = n45895 ^ n43234;
  assign n45898 = n45895 & n43234;
  assign n45896 = ~n45895;
  assign n45897 = n45910 ^ n45911;
  assign n45864 = n45911 & n45910;
  assign n45943 = n45913 & n13583;
  assign n45941 = ~n45957;
  assign n45944 = ~n45913;
  assign n45974 = ~n45994;
  assign n45816 = n256 ^ n45836;
  assign n45827 = n45839 & n10976;
  assign n45799 = ~n45840;
  assign n45852 = n45858 & n45859;
  assign n45841 = n45862 & n45863;
  assign n45821 = n45869 & n45870;
  assign n41952 = n45871 ^ n45872;
  assign n45888 = n45896 & n43201;
  assign n45889 = n45897 & n43165;
  assign n45876 = ~n45898;
  assign n45811 = ~n45897;
  assign n45912 = n45941 & n45942;
  assign n45915 = ~n45943;
  assign n45932 = n45944 & n121;
  assign n45945 = n45974 & n45975;
  assign n43836 = n45815 ^ n45816;
  assign n45774 = n45816 & n45815;
  assign n45820 = ~n45827;
  assign n45822 = n45841 ^ n45842;
  assign n45837 = ~n45852;
  assign n45831 = ~n45841;
  assign n45849 = n41952 & n44651;
  assign n45850 = n45821 & n45853;
  assign n45851 = n41952 & n43234;
  assign n45848 = ~n45821;
  assign n41920 = ~n41952;
  assign n45873 = n45876 & n45872;
  assign n45855 = ~n45888;
  assign n45834 = ~n45889;
  assign n45877 = n45811 & n43187;
  assign n45890 = n45912 ^ n45913;
  assign n45914 = ~n45912;
  assign n45892 = ~n45932;
  assign n45916 = n120 ^ n45945;
  assign n44857 = ~n43836;
  assign n45777 = ~n45774;
  assign n45779 = n45821 ^ n45822;
  assign n45817 = n45837 & n45838;
  assign n45843 = n45848 & n45842;
  assign n45828 = ~n45849;
  assign n45830 = ~n45850;
  assign n44701 = ~n45851;
  assign n45854 = ~n45873;
  assign n45814 = ~n45877;
  assign n45865 = n121 ^ n45890;
  assign n45902 = n45914 & n45915;
  assign n45824 = n45916 ^ n45917;
  assign n45801 = n45779 & n270;
  assign n45800 = ~n45779;
  assign n45797 = n45817 ^ n45818;
  assign n45819 = ~n45817;
  assign n45766 = n45828 & n45829;
  assign n45825 = n45830 & n45831;
  assign n45807 = ~n45843;
  assign n45832 = n45854 & n45855;
  assign n45771 = n45864 ^ n45865;
  assign n45866 = ~n45865;
  assign n45891 = ~n45902;
  assign n45775 = n271 ^ n45797;
  assign n45786 = n45800 & n10896;
  assign n45760 = ~n45801;
  assign n45805 = n45819 & n45820;
  assign n45810 = n45766 & n45788;
  assign n45808 = ~n45766;
  assign n45806 = ~n45825;
  assign n45812 = n45832 ^ n43165;
  assign n45833 = ~n45832;
  assign n45844 = n45771 & n43124;
  assign n45845 = ~n45771;
  assign n45847 = n45866 & n45864;
  assign n45846 = n45891 & n45892;
  assign n43796 = n45774 ^ n45775;
  assign n45776 = ~n45775;
  assign n45781 = ~n45786;
  assign n45798 = ~n45805;
  assign n45787 = n45806 & n45807;
  assign n45804 = n45808 & n45809;
  assign n45790 = ~n45810;
  assign n41905 = n45811 ^ n45812;
  assign n45826 = n45833 & n45834;
  assign n45773 = ~n45844;
  assign n45835 = n45845 & n43156;
  assign n45823 = n45846 ^ n45847;
  assign n44773 = ~n43796;
  assign n45735 = n45776 & n45777;
  assign n45767 = n45787 ^ n45788;
  assign n45778 = n45798 & n45799;
  assign n45791 = n41905 & n44566;
  assign n45792 = n41905 & n43165;
  assign n45789 = ~n45787;
  assign n45769 = ~n45804;
  assign n41931 = ~n41905;
  assign n45731 = n45823 ^ n45824;
  assign n45813 = ~n45826;
  assign n45795 = ~n45835;
  assign n45739 = n45766 ^ n45767;
  assign n45758 = n45778 ^ n45779;
  assign n45780 = ~n45778;
  assign n45784 = n45789 & n45790;
  assign n45782 = ~n45791;
  assign n44607 = ~n45792;
  assign n45803 = n45731 & n43113;
  assign n45793 = n45813 & n45814;
  assign n45802 = ~n45731;
  assign n45736 = n270 ^ n45758;
  assign n45750 = n45739 & n10806;
  assign n45751 = ~n45739;
  assign n45765 = n45780 & n45781;
  assign n45726 = n45782 & n45783;
  assign n45768 = ~n45784;
  assign n45770 = n45793 ^ n43156;
  assign n45796 = n45802 & n43081;
  assign n45734 = ~n45803;
  assign n45794 = ~n45793;
  assign n43777 = n45735 ^ n45736;
  assign n45737 = ~n45736;
  assign n45740 = ~n45750;
  assign n45745 = n45751 & n269;
  assign n45762 = n45726 & n45763;
  assign n45759 = ~n45765;
  assign n45761 = ~n45726;
  assign n45764 = n45768 & n45769;
  assign n41862 = n45770 ^ n45771;
  assign n45785 = n45794 & n45795;
  assign n45757 = ~n45796;
  assign n44670 = ~n43777;
  assign n45698 = n45737 & n45735;
  assign n45721 = ~n45745;
  assign n45738 = n45759 & n45760;
  assign n45752 = n45761 & n45748;
  assign n45753 = n41862 & n44489;
  assign n45746 = ~n45762;
  assign n45754 = n41862 & n43156;
  assign n45747 = ~n45764;
  assign n41871 = ~n41862;
  assign n45772 = ~n45785;
  assign n45697 = ~n45698;
  assign n45719 = n45738 ^ n45739;
  assign n45744 = n45746 & n45747;
  assign n45727 = n45747 ^ n45748;
  assign n45741 = ~n45738;
  assign n45729 = ~n45752;
  assign n45742 = ~n45753;
  assign n44527 = ~n45754;
  assign n45755 = n45772 & n45773;
  assign n45699 = n269 ^ n45719;
  assign n45701 = n45726 ^ n45727;
  assign n45730 = n45740 & n45741;
  assign n45685 = n45742 & n45743;
  assign n45728 = ~n45744;
  assign n45732 = n45755 ^ n43081;
  assign n45756 = ~n45755;
  assign n43717 = n45698 ^ n45699;
  assign n45696 = ~n45699;
  assign n45707 = n45701 & n10723;
  assign n45708 = ~n45701;
  assign n45709 = n45728 & n45729;
  assign n45724 = n45685 & n45710;
  assign n45720 = ~n45730;
  assign n45722 = ~n45685;
  assign n41829 = n45731 ^ n45732;
  assign n45749 = n45756 & n45757;
  assign n44603 = ~n43717;
  assign n45661 = n45696 & n45697;
  assign n45693 = ~n45707;
  assign n45702 = n45708 & n268;
  assign n45686 = n45709 ^ n45710;
  assign n45712 = ~n45709;
  assign n45700 = n45720 & n45721;
  assign n45714 = n45722 & n45723;
  assign n45711 = ~n45724;
  assign n45715 = n41829 & n44401;
  assign n45716 = n41829 & n43081;
  assign n41804 = ~n41829;
  assign n45733 = ~n45749;
  assign n45641 = n45685 ^ n45686;
  assign n45669 = ~n45661;
  assign n45680 = n45700 ^ n45701;
  assign n45678 = ~n45702;
  assign n45703 = n45711 & n45712;
  assign n45692 = ~n45700;
  assign n45689 = ~n45714;
  assign n45704 = ~n45715;
  assign n44435 = ~n45716;
  assign n45725 = n45733 & n45734;
  assign n45670 = n45641 & n10627;
  assign n45662 = n268 ^ n45680;
  assign n45668 = ~n45641;
  assign n45687 = n45692 & n45693;
  assign n45688 = ~n45703;
  assign n45651 = n45704 & n45705;
  assign n45718 = n45725 & n43072;
  assign n45717 = ~n45725;
  assign n43703 = n45661 ^ n45662;
  assign n45663 = n45668 & n267;
  assign n45620 = n45662 & n45669;
  assign n45657 = ~n45670;
  assign n45677 = ~n45687;
  assign n45671 = n45688 & n45689;
  assign n45682 = n45651 & n45690;
  assign n45681 = ~n45651;
  assign n45713 = n45717 & n43038;
  assign n45695 = ~n45718;
  assign n45623 = ~n45620;
  assign n45643 = ~n45663;
  assign n45652 = n45671 ^ n45672;
  assign n45659 = n45677 & n45678;
  assign n45674 = ~n45671;
  assign n45679 = n45681 & n45672;
  assign n45673 = ~n45682;
  assign n45694 = n45695 & n45706;
  assign n45684 = ~n45713;
  assign n45625 = n45651 ^ n45652;
  assign n45640 = n267 ^ n45659;
  assign n45658 = ~n45659;
  assign n45664 = n45673 & n45674;
  assign n45654 = ~n45679;
  assign n45683 = ~n45694;
  assign n45691 = n45684 & n45695;
  assign n45621 = n45640 ^ n45641;
  assign n45638 = n45625 & n266;
  assign n45637 = ~n45625;
  assign n45650 = n45657 & n45658;
  assign n45653 = ~n45664;
  assign n45665 = n45683 & n45684;
  assign n45675 = ~n45691;
  assign n45602 = n45620 ^ n45621;
  assign n45622 = ~n45621;
  assign n45632 = n45637 & n10589;
  assign n45597 = ~n45638;
  assign n45642 = ~n45650;
  assign n45639 = n45653 & n45654;
  assign n45647 = n45665 ^ n43024;
  assign n41772 = n45675 ^ n45676;
  assign n45666 = ~n45665;
  assign n41413 = n45602 ^ n42460;
  assign n45603 = ~n45602;
  assign n45578 = n45622 & n45623;
  assign n45615 = ~n45632;
  assign n45618 = n45639 ^ n45633;
  assign n45624 = n45642 & n45643;
  assign n45612 = ~n45639;
  assign n41732 = n45646 ^ n45647;
  assign n45655 = n41772 & n44327;
  assign n45656 = n41772 & n43072;
  assign n45660 = n45666 & n45667;
  assign n41801 = ~n41772;
  assign n41415 = ~n41413;
  assign n45507 = n45603 & n42460;
  assign n45598 = n45603 & n42462;
  assign n45581 = ~n45578;
  assign n45604 = n45624 ^ n45625;
  assign n45616 = ~n45624;
  assign n41756 = ~n41732;
  assign n45644 = ~n45655;
  assign n44385 = ~n45656;
  assign n45648 = ~n45660;
  assign n45573 = n41415 & n43602;
  assign n43615 = ~n45598;
  assign n45579 = n266 ^ n45604;
  assign n45606 = n45615 & n45616;
  assign n45626 = n41756 & n44270;
  assign n45627 = n41756 & n42998;
  assign n45617 = n45644 & n45645;
  assign n45634 = n45648 & n45649;
  assign n45557 = ~n45573;
  assign n45564 = n45578 ^ n45579;
  assign n45580 = ~n45579;
  assign n45596 = ~n45606;
  assign n45575 = n45617 ^ n45618;
  assign n45607 = ~n45626;
  assign n44308 = ~n45627;
  assign n45630 = n45617 & n45633;
  assign n45610 = n45634 ^ n42966;
  assign n45628 = ~n45617;
  assign n45635 = ~n45634;
  assign n45534 = n45557 & n45558;
  assign n45559 = n45564 & n42355;
  assign n45560 = ~n45564;
  assign n45530 = n45580 & n45581;
  assign n45574 = n45596 & n45597;
  assign n45599 = n45575 & n10522;
  assign n45600 = ~n45575;
  assign n45540 = n45607 & n45608;
  assign n41674 = n45609 ^ n45610;
  assign n45619 = n45628 & n45629;
  assign n45611 = ~n45630;
  assign n45631 = n45635 & n45636;
  assign n45519 = n45534 ^ n45535;
  assign n45144 = n45534 ^ n45536;
  assign n45538 = ~n45534;
  assign n45511 = ~n45559;
  assign n45553 = n45560 & n42364;
  assign n45554 = n45574 ^ n45575;
  assign n45576 = ~n45574;
  assign n45577 = ~n45599;
  assign n45587 = n45600 & n265;
  assign n45589 = n45540 & n45601;
  assign n45588 = ~n45540;
  assign n41713 = ~n41674;
  assign n45605 = n45611 & n45612;
  assign n45591 = ~n45619;
  assign n45613 = ~n45631;
  assign n45399 = n45519 & n423;
  assign n45170 = ~n45144;
  assign n45508 = n45538 & n45539;
  assign n45537 = ~n45553;
  assign n45531 = n265 ^ n45554;
  assign n45565 = n45576 & n45577;
  assign n45556 = ~n45587;
  assign n45582 = n45588 & n45563;
  assign n45583 = n41713 & n44202;
  assign n45568 = ~n45589;
  assign n45584 = n41713 & n42966;
  assign n45590 = ~n45605;
  assign n45592 = n45613 & n45614;
  assign n45486 = n45399 & n422;
  assign n45485 = ~n45399;
  assign n45432 = n45508 ^ n45509;
  assign n45513 = n45508 & n45520;
  assign n45512 = ~n45508;
  assign n45452 = n45530 ^ n45531;
  assign n45529 = n45537 & n45507;
  assign n45506 = n45537 & n45511;
  assign n45453 = n45531 & n45530;
  assign n45555 = ~n45565;
  assign n45545 = ~n45582;
  assign n45566 = ~n45583;
  assign n44260 = ~n45584;
  assign n45585 = n45590 & n45591;
  assign n45569 = n45592 ^ n45593;
  assign n45594 = ~n45592;
  assign n45476 = n45485 & n7609;
  assign n45386 = ~n45486;
  assign n41299 = n45506 ^ n45507;
  assign n45499 = n45512 & n45509;
  assign n45500 = n45452 & n42287;
  assign n45403 = ~n45513;
  assign n45501 = ~n45452;
  assign n45510 = ~n45529;
  assign n45514 = n45555 & n45556;
  assign n45522 = n45566 & n45567;
  assign n41654 = n42883 ^ n45569;
  assign n45570 = n45569 & n42952;
  assign n45562 = ~n45585;
  assign n45586 = n45594 & n45595;
  assign n45418 = ~n45476;
  assign n45478 = n41299 & n42364;
  assign n45477 = n41299 & n43547;
  assign n41313 = ~n41299;
  assign n45433 = ~n45499;
  assign n45450 = ~n45500;
  assign n45487 = n45501 & n42305;
  assign n45479 = n45510 & n45511;
  assign n45491 = ~n45514;
  assign n45548 = n45522 & n45489;
  assign n45549 = n41654 & n44162;
  assign n45546 = ~n45522;
  assign n41666 = ~n41654;
  assign n45541 = n45562 ^ n45563;
  assign n45561 = n45568 & n45562;
  assign n44225 = ~n45570;
  assign n45571 = ~n45586;
  assign n45457 = ~n45477;
  assign n43561 = ~n45478;
  assign n45451 = n45479 ^ n42305;
  assign n45474 = ~n45487;
  assign n45475 = ~n45479;
  assign n45515 = n45540 ^ n45541;
  assign n45542 = n45546 & n45547;
  assign n45524 = ~n45548;
  assign n45532 = ~n45549;
  assign n45544 = ~n45561;
  assign n45550 = n45571 & n45572;
  assign n41250 = n45451 ^ n45452;
  assign n45431 = n45457 & n45458;
  assign n45459 = n45474 & n45475;
  assign n45480 = n45514 ^ n45515;
  assign n45516 = n45515 & n10470;
  assign n45438 = n45532 & n45533;
  assign n45517 = ~n45515;
  assign n45493 = ~n45542;
  assign n45521 = n45544 & n45545;
  assign n45525 = n45550 ^ n42913;
  assign n45551 = ~n45550;
  assign n45423 = n41250 & n43521;
  assign n45424 = n41250 & n42305;
  assign n45400 = n45431 ^ n45432;
  assign n41204 = ~n41250;
  assign n45434 = ~n45431;
  assign n45449 = ~n45459;
  assign n45454 = n264 ^ n45480;
  assign n45490 = ~n45516;
  assign n45504 = n45438 & n45465;
  assign n45505 = n45517 & n264;
  assign n45488 = n45521 ^ n45522;
  assign n45502 = ~n45438;
  assign n41602 = n45525 ^ n45526;
  assign n45523 = ~n45521;
  assign n45543 = n45551 & n45552;
  assign n45363 = n45399 ^ n45400;
  assign n45401 = n45418 & n45400;
  assign n45397 = ~n45423;
  assign n43533 = ~n45424;
  assign n45425 = n45433 & n45434;
  assign n45419 = n45449 & n45450;
  assign n45388 = n45453 ^ n45454;
  assign n45369 = n45454 & n45453;
  assign n45405 = n45488 ^ n45489;
  assign n45481 = n45490 & n45491;
  assign n45494 = n45502 & n45503;
  assign n45468 = ~n45504;
  assign n45463 = ~n45505;
  assign n41643 = ~n41602;
  assign n45518 = n45523 & n45524;
  assign n45527 = ~n45543;
  assign n45332 = n422 ^ n45363;
  assign n45333 = n45397 & n45398;
  assign n45385 = ~n45401;
  assign n45387 = n45419 ^ n42261;
  assign n45402 = ~n45425;
  assign n45394 = ~n45419;
  assign n45426 = n45388 & n42228;
  assign n45427 = ~n45388;
  assign n45460 = n45405 & n10418;
  assign n45461 = ~n45405;
  assign n45462 = ~n45481;
  assign n45441 = ~n45494;
  assign n45482 = n41643 & n44132;
  assign n45483 = n41643 & n42913;
  assign n45492 = ~n45518;
  assign n45495 = n45527 & n45528;
  assign n43425 = n45332 ^ n45144;
  assign n45221 = n45332 & n45144;
  assign n45293 = n45385 & n45386;
  assign n41141 = n45387 ^ n45388;
  assign n45353 = ~n45333;
  assign n45364 = n45402 & n45403;
  assign n45360 = ~n45426;
  assign n45420 = n45427 & n42261;
  assign n45435 = ~n45460;
  assign n45455 = n45461 & n279;
  assign n45437 = n45462 & n45463;
  assign n45466 = ~n45482;
  assign n44184 = ~n45483;
  assign n45464 = n45492 & n45493;
  assign n45470 = n45495 ^ n45496;
  assign n45497 = ~n45495;
  assign n45061 = ~n43425;
  assign n45224 = ~n45221;
  assign n45351 = n45293 & n7523;
  assign n45354 = n41141 & n43481;
  assign n45355 = n41141 & n42261;
  assign n45350 = ~n45293;
  assign n45334 = n45364 ^ n45365;
  assign n41159 = ~n41141;
  assign n45368 = n45364 & n45365;
  assign n45366 = ~n45364;
  assign n45393 = ~n45420;
  assign n45404 = n279 ^ n45437;
  assign n45407 = ~n45455;
  assign n45436 = ~n45437;
  assign n45439 = n45464 ^ n45465;
  assign n45375 = n45466 & n45467;
  assign n41563 = n42827 ^ n45470;
  assign n45471 = n45470 & n42873;
  assign n45469 = ~n45464;
  assign n45484 = n45497 & n45498;
  assign n45294 = n45333 ^ n45334;
  assign n45335 = n45350 & n421;
  assign n45295 = ~n45351;
  assign n45323 = ~n45354;
  assign n43504 = ~n45355;
  assign n45358 = n45366 & n45367;
  assign n45352 = ~n45368;
  assign n45389 = n45393 & n45394;
  assign n45370 = n45404 ^ n45405;
  assign n45428 = n45435 & n45436;
  assign n45372 = n45438 ^ n45439;
  assign n45444 = n41563 & n44096;
  assign n45445 = n45375 & n45411;
  assign n45442 = ~n45375;
  assign n41605 = ~n41563;
  assign n45456 = n45468 & n45469;
  assign n44127 = ~n45471;
  assign n45472 = ~n45484;
  assign n45262 = n45293 ^ n45294;
  assign n45296 = ~n45294;
  assign n45246 = n45323 & n45324;
  assign n45264 = ~n45335;
  assign n45336 = n45352 & n45353;
  assign n45320 = ~n45358;
  assign n45288 = n45369 ^ n45370;
  assign n45359 = ~n45389;
  assign n45297 = n45370 & n45369;
  assign n45408 = n45372 & n10398;
  assign n45406 = ~n45428;
  assign n45409 = ~n45372;
  assign n45429 = n45442 & n45443;
  assign n45421 = ~n45444;
  assign n45413 = ~n45445;
  assign n45440 = ~n45456;
  assign n45446 = n45472 & n45473;
  assign n45222 = n421 ^ n45262;
  assign n45286 = n45295 & n45296;
  assign n45254 = ~n45246;
  assign n45319 = ~n45336;
  assign n45337 = n45288 & n42189;
  assign n45325 = n45359 & n45360;
  assign n45338 = ~n45288;
  assign n45302 = ~n45297;
  assign n45371 = n45406 & n45407;
  assign n45373 = ~n45408;
  assign n45395 = n45409 & n278;
  assign n45307 = n45421 & n45422;
  assign n45378 = ~n45429;
  assign n45410 = n45440 & n45441;
  assign n45414 = n45446 ^ n42832;
  assign n45447 = ~n45446;
  assign n43393 = n45221 ^ n45222;
  assign n45223 = ~n45222;
  assign n45263 = ~n45286;
  assign n45279 = n45319 & n45320;
  assign n45287 = n45325 ^ n42216;
  assign n45261 = ~n45337;
  assign n45326 = n45338 & n42216;
  assign n45300 = ~n45325;
  assign n45339 = n45371 ^ n45372;
  assign n45374 = ~n45371;
  assign n45331 = ~n45395;
  assign n45392 = n45307 & n45343;
  assign n45376 = n45410 ^ n45411;
  assign n45390 = ~n45307;
  assign n41524 = n45414 ^ n45415;
  assign n45412 = ~n45410;
  assign n45430 = n45447 & n45448;
  assign n44968 = ~n43393;
  assign n45122 = n45223 & n45224;
  assign n45252 = n45263 & n45264;
  assign n45247 = n45279 ^ n45280;
  assign n45283 = n45279 & n45280;
  assign n41041 = n45287 ^ n45288;
  assign n45281 = ~n45279;
  assign n45299 = ~n45326;
  assign n45298 = n278 ^ n45339;
  assign n45361 = n45373 & n45374;
  assign n45304 = n45375 ^ n45376;
  assign n45379 = n45390 & n45391;
  assign n45380 = n41524 & n44063;
  assign n45344 = ~n45392;
  assign n45381 = n41524 & n42832;
  assign n41566 = ~n41524;
  assign n45396 = n45412 & n45413;
  assign n45416 = ~n45430;
  assign n45125 = ~n45122;
  assign n45206 = n45246 ^ n45247;
  assign n45177 = ~n45252;
  assign n45255 = n41041 & n43453;
  assign n45256 = n41041 & n42216;
  assign n45265 = n45281 & n45282;
  assign n45253 = ~n45283;
  assign n41084 = ~n41041;
  assign n45190 = n45297 ^ n45298;
  assign n45289 = n45299 & n45300;
  assign n45301 = ~n45298;
  assign n45340 = n45304 & n10372;
  assign n45330 = ~n45361;
  assign n45341 = ~n45304;
  assign n45310 = ~n45379;
  assign n45356 = ~n45380;
  assign n44071 = ~n45381;
  assign n45377 = ~n45396;
  assign n45382 = n45416 & n45417;
  assign n45166 = n45177 ^ n45206;
  assign n45207 = n45206 & n7437;
  assign n45208 = ~n45206;
  assign n45248 = n45253 & n45254;
  assign n45225 = ~n45255;
  assign n43471 = ~n45256;
  assign n45214 = ~n45265;
  assign n45209 = ~n45190;
  assign n45260 = ~n45289;
  assign n45219 = n45301 & n45302;
  assign n45303 = n45330 & n45331;
  assign n45305 = ~n45340;
  assign n45327 = n45341 & n277;
  assign n45234 = n45356 & n45357;
  assign n45342 = n45377 & n45378;
  assign n45347 = n45382 ^ n42744;
  assign n45383 = ~n45382;
  assign n45123 = n420 ^ n45166;
  assign n45176 = ~n45207;
  assign n45186 = n45208 & n420;
  assign n45135 = n45225 & n45226;
  assign n45213 = ~n45248;
  assign n45227 = n45260 & n45261;
  assign n45249 = ~n45219;
  assign n45266 = n45303 ^ n45304;
  assign n45306 = ~n45303;
  assign n45268 = ~n45327;
  assign n45322 = n45234 & n45328;
  assign n45308 = n45342 ^ n45343;
  assign n45321 = ~n45234;
  assign n41515 = n45346 ^ n45347;
  assign n45345 = ~n45342;
  assign n45362 = n45383 & n45384;
  assign n43362 = n45122 ^ n45123;
  assign n45124 = ~n45123;
  assign n45167 = n45176 & n45177;
  assign n45134 = ~n45186;
  assign n45189 = n45135 & n45179;
  assign n45187 = ~n45135;
  assign n45178 = n45213 & n45214;
  assign n45191 = n45227 ^ n42142;
  assign n45229 = n45227 & n42167;
  assign n45228 = ~n45227;
  assign n45220 = n277 ^ n45266;
  assign n45290 = n45305 & n45306;
  assign n45231 = n45307 ^ n45308;
  assign n45311 = n45321 & n45272;
  assign n45312 = n41515 & n44003;
  assign n45274 = ~n45322;
  assign n45314 = n41515 & n44080;
  assign n45315 = n41515 & n42744;
  assign n41483 = ~n41515;
  assign n45329 = n45344 & n45345;
  assign n45348 = ~n45362;
  assign n44881 = ~n43362;
  assign n45018 = n45124 & n45125;
  assign n45133 = ~n45167;
  assign n45136 = n45178 ^ n45179;
  assign n45180 = n45187 & n45188;
  assign n45169 = ~n45189;
  assign n40967 = n45190 ^ n45191;
  assign n45168 = ~n45178;
  assign n45093 = n45219 ^ n45220;
  assign n45215 = n45228 & n42142;
  assign n45210 = ~n45229;
  assign n45148 = n45220 & n45249;
  assign n45269 = n45231 & n10334;
  assign n45267 = ~n45290;
  assign n45270 = ~n45231;
  assign n45237 = ~n45311;
  assign n45284 = ~n45312;
  assign n45291 = n41483 & n45313;
  assign n44082 = ~n45314;
  assign n44037 = ~n45315;
  assign n45309 = ~n45329;
  assign n45316 = n45348 & n45349;
  assign n45097 = n45133 & n45134;
  assign n45098 = n45135 ^ n45136;
  assign n43486 = n45144 ^ n40967;
  assign n45143 = n45168 & n45169;
  assign n45145 = n40967 & n43407;
  assign n45146 = n40967 & n45170;
  assign n45147 = n40967 & n42167;
  assign n45127 = ~n45180;
  assign n41011 = ~n40967;
  assign n45193 = n45093 & n42117;
  assign n45194 = n45209 & n45210;
  assign n45192 = ~n45093;
  assign n45172 = ~n45215;
  assign n45151 = ~n45148;
  assign n45230 = n45267 & n45268;
  assign n45233 = ~n45269;
  assign n45257 = n45270 & n276;
  assign n45199 = n45284 & n45285;
  assign n44101 = ~n45291;
  assign n45271 = n45309 & n45310;
  assign n45276 = n45316 ^ n42748;
  assign n45317 = ~n45316;
  assign n45057 = n45097 ^ n45098;
  assign n45099 = n45098 & n7333;
  assign n45068 = ~n45097;
  assign n45100 = ~n45098;
  assign n45126 = ~n45143;
  assign n45128 = ~n45145;
  assign n45137 = n41011 & n45144;
  assign n43465 = ~n45146;
  assign n43456 = ~n45147;
  assign n45181 = n45192 & n42097;
  assign n45132 = ~n45193;
  assign n45171 = ~n45194;
  assign n45195 = n45230 ^ n45231;
  assign n45232 = ~n45230;
  assign n45185 = ~n45257;
  assign n45251 = n45199 & n45258;
  assign n45235 = n45271 ^ n45272;
  assign n45250 = ~n45199;
  assign n41433 = n45275 ^ n45276;
  assign n45273 = ~n45271;
  assign n45292 = n45317 & n45318;
  assign n45019 = n419 ^ n45057;
  assign n45067 = ~n45099;
  assign n45086 = n45100 & n419;
  assign n45087 = n45126 & n45127;
  assign n45049 = n45128 & n45129;
  assign n43488 = ~n45137;
  assign n45130 = n45171 & n45172;
  assign n45095 = ~n45181;
  assign n45149 = n276 ^ n45195;
  assign n45216 = n45232 & n45233;
  assign n45153 = n45234 ^ n45235;
  assign n45238 = n45250 & n45157;
  assign n45239 = n41433 & n43964;
  assign n45240 = n41433 & n44040;
  assign n45201 = ~n45251;
  assign n45242 = n41433 & n42706;
  assign n41486 = ~n41433;
  assign n45259 = n45273 & n45274;
  assign n45277 = ~n45292;
  assign n43327 = n45018 ^ n45019;
  assign n44906 = n45019 & n45018;
  assign n45058 = n45067 & n45068;
  assign n45027 = ~n45086;
  assign n45050 = n45087 ^ n45088;
  assign n45091 = n45049 & n45088;
  assign n45060 = ~n45087;
  assign n45089 = ~n45049;
  assign n45092 = n45130 ^ n42117;
  assign n45012 = n45148 ^ n45149;
  assign n45131 = ~n45130;
  assign n45150 = ~n45149;
  assign n45197 = n45153 & n275;
  assign n45184 = ~n45216;
  assign n45196 = ~n45153;
  assign n45159 = ~n45238;
  assign n45211 = ~n45239;
  assign n44042 = ~n45240;
  assign n45217 = n41486 & n45241;
  assign n44005 = ~n45242;
  assign n45236 = ~n45259;
  assign n45243 = n45277 & n45278;
  assign n44800 = ~n43327;
  assign n44986 = n45049 ^ n45050;
  assign n45026 = ~n45058;
  assign n45069 = n45089 & n45090;
  assign n45059 = ~n45091;
  assign n40892 = n45092 ^ n45093;
  assign n45107 = n45012 & n42075;
  assign n45108 = n45131 & n45132;
  assign n45106 = ~n45012;
  assign n45070 = n45150 & n45151;
  assign n45152 = n45184 & n45185;
  assign n45182 = n45196 & n10269;
  assign n45105 = ~n45197;
  assign n45076 = n45211 & n45212;
  assign n44067 = ~n45217;
  assign n45198 = n45236 & n45237;
  assign n45203 = n45243 ^ n42660;
  assign n45244 = ~n45243;
  assign n45007 = n44986 & n7273;
  assign n44985 = n45026 & n45027;
  assign n45008 = ~n44986;
  assign n45051 = n45059 & n45060;
  assign n45052 = n40892 & n45061;
  assign n45021 = ~n45069;
  assign n40905 = ~n40892;
  assign n45101 = n45106 & n42062;
  assign n45054 = ~n45107;
  assign n45094 = ~n45108;
  assign n45109 = n45152 ^ n45153;
  assign n45155 = ~n45152;
  assign n45154 = ~n45182;
  assign n45175 = n45076 & n45113;
  assign n45156 = n45198 ^ n45199;
  assign n45173 = ~n45076;
  assign n41443 = n45202 ^ n45203;
  assign n45200 = ~n45198;
  assign n45218 = n45244 & n45245;
  assign n44947 = n44985 ^ n44986;
  assign n44978 = ~n45007;
  assign n44987 = n45008 & n418;
  assign n44977 = ~n44985;
  assign n45020 = ~n45051;
  assign n45028 = n40905 & n43374;
  assign n43448 = ~n45052;
  assign n45029 = n40905 & n42117;
  assign n45030 = n40905 & n43425;
  assign n45053 = n45094 & n45095;
  assign n45014 = ~n45101;
  assign n45071 = n275 ^ n45109;
  assign n45138 = n45154 & n45155;
  assign n45073 = n45156 ^ n45157;
  assign n45160 = n45173 & n45174;
  assign n45115 = ~n45175;
  assign n45161 = n41443 & n43998;
  assign n41437 = ~n41443;
  assign n45183 = n45200 & n45201;
  assign n45204 = ~n45218;
  assign n44907 = n418 ^ n44947;
  assign n44964 = n44977 & n44978;
  assign n44939 = ~n44987;
  assign n44979 = n45020 & n45021;
  assign n45009 = ~n45028;
  assign n43400 = ~n45029;
  assign n43428 = ~n45030;
  assign n45011 = n45053 ^ n42075;
  assign n44928 = n45070 ^ n45071;
  assign n45055 = ~n45053;
  assign n44988 = n45071 & n45070;
  assign n45111 = n45073 & n274;
  assign n45104 = ~n45138;
  assign n45110 = ~n45073;
  assign n45079 = ~n45160;
  assign n45139 = n41437 & n43922;
  assign n45140 = n41437 & n42660;
  assign n44024 = ~n45161;
  assign n45141 = n41437 & n45162;
  assign n45158 = ~n45183;
  assign n45163 = n45204 & n45205;
  assign n43308 = n44906 ^ n44907;
  assign n44812 = n44907 & n44906;
  assign n44938 = ~n44964;
  assign n44941 = n44979 ^ n44966;
  assign n44940 = n45009 & n45010;
  assign n44943 = ~n44979;
  assign n40831 = n45011 ^ n45012;
  assign n45031 = n44928 & n42040;
  assign n45033 = n45054 & n45055;
  assign n45032 = ~n44928;
  assign n44991 = ~n44988;
  assign n45072 = n45104 & n45105;
  assign n45102 = n45110 & n10216;
  assign n45036 = ~n45111;
  assign n45116 = ~n45139;
  assign n43954 = ~n45140;
  assign n44001 = ~n45141;
  assign n45112 = n45158 & n45159;
  assign n45118 = n45163 ^ n42667;
  assign n45164 = ~n45163;
  assign n44718 = ~n43308;
  assign n44896 = n44938 & n44939;
  assign n44897 = n44940 ^ n44941;
  assign n44967 = n40831 & n43393;
  assign n44969 = n44940 & n44980;
  assign n44965 = ~n44940;
  assign n40860 = ~n40831;
  assign n44971 = ~n45031;
  assign n45022 = n45032 & n42018;
  assign n45013 = ~n45033;
  assign n45034 = n45072 ^ n45073;
  assign n45074 = ~n45072;
  assign n45075 = ~n45102;
  assign n45077 = n45112 ^ n45113;
  assign n44996 = n45116 & n45117;
  assign n41290 = n45118 ^ n45119;
  assign n45114 = ~n45112;
  assign n45142 = n45164 & n45165;
  assign n44858 = n44896 ^ n44897;
  assign n44899 = n44897 & n417;
  assign n44860 = ~n44896;
  assign n44898 = ~n44897;
  assign n44948 = n44965 & n44966;
  assign n44949 = n40860 & n43343;
  assign n43415 = ~n44967;
  assign n44950 = n40860 & n44968;
  assign n44942 = ~n44969;
  assign n44951 = n40860 & n42075;
  assign n44970 = n45013 & n45014;
  assign n44931 = ~n45022;
  assign n44989 = n274 ^ n45034;
  assign n45062 = n45074 & n45075;
  assign n44993 = n45076 ^ n45077;
  assign n45080 = n41290 & n45096;
  assign n45016 = ~n44996;
  assign n41379 = ~n41290;
  assign n45103 = n45114 & n45115;
  assign n45120 = ~n45142;
  assign n44813 = n417 ^ n44858;
  assign n44880 = n44898 & n7227;
  assign n44816 = ~n44899;
  assign n44925 = n44942 & n44943;
  assign n44901 = ~n44948;
  assign n44926 = ~n44949;
  assign n43396 = ~n44950;
  assign n43361 = ~n44951;
  assign n44929 = n44970 ^ n42018;
  assign n44972 = ~n44970;
  assign n44846 = n44988 ^ n44989;
  assign n44990 = ~n44989;
  assign n45037 = n44993 & n10199;
  assign n45035 = ~n45062;
  assign n45038 = ~n44993;
  assign n45063 = n41379 & n43869;
  assign n43981 = ~n45080;
  assign n45064 = n41379 & n45081;
  assign n45065 = n41379 & n42667;
  assign n45078 = ~n45103;
  assign n45082 = n45120 & n45121;
  assign n43247 = n44812 ^ n44813;
  assign n44814 = ~n44813;
  assign n44859 = ~n44880;
  assign n44900 = ~n44925;
  assign n44817 = n44926 & n44927;
  assign n40780 = n44928 ^ n44929;
  assign n44953 = n44846 & n41991;
  assign n44954 = n44971 & n44972;
  assign n44952 = ~n44846;
  assign n44908 = n44990 & n44991;
  assign n44992 = n45035 & n45036;
  assign n44995 = ~n45037;
  assign n45023 = n45038 & n273;
  assign n45041 = ~n45063;
  assign n43959 = ~n45064;
  assign n43946 = ~n45065;
  assign n45039 = n45078 & n45079;
  assign n45045 = n45082 ^ n45083;
  assign n45084 = ~n45082;
  assign n44646 = ~n43247;
  assign n44691 = n44814 & n44812;
  assign n44844 = n44859 & n44860;
  assign n44882 = n40780 & n43362;
  assign n44861 = n44900 & n44901;
  assign n44884 = n44817 & n44902;
  assign n44885 = n40780 & n43281;
  assign n44886 = n40780 & n42040;
  assign n44883 = ~n44817;
  assign n40761 = ~n40780;
  assign n44944 = n44952 & n41980;
  assign n44843 = ~n44953;
  assign n44930 = ~n44954;
  assign n44911 = ~n44908;
  assign n44955 = n44992 ^ n44993;
  assign n44994 = ~n44992;
  assign n44957 = ~n45023;
  assign n44997 = n45039 ^ n45040;
  assign n44933 = n45041 & n45042;
  assign n45025 = n43981 & n43959;
  assign n41327 = n45045 ^ n42622;
  assign n45044 = n45039 & n45056;
  assign n45046 = n45045 & n42555;
  assign n45043 = ~n45039;
  assign n45066 = n45084 & n45085;
  assign n44815 = ~n44844;
  assign n44818 = n44861 ^ n44862;
  assign n44868 = n40761 & n44881;
  assign n43365 = ~n44882;
  assign n44864 = ~n44861;
  assign n44869 = n44883 & n44862;
  assign n44863 = ~n44884;
  assign n44865 = ~n44885;
  assign n43325 = ~n44886;
  assign n44887 = n44930 & n44931;
  assign n44889 = ~n44944;
  assign n44909 = n273 ^ n44955;
  assign n44981 = n44994 & n44995;
  assign n44913 = n44996 ^ n44997;
  assign n45001 = n41327 & n43846;
  assign n45002 = n44933 & n44891;
  assign n45003 = n41327 & n45017;
  assign n44999 = ~n44933;
  assign n43979 = ~n45025;
  assign n41264 = ~n41327;
  assign n45024 = n45043 & n45040;
  assign n45015 = ~n45044;
  assign n43888 = ~n45046;
  assign n45047 = ~n45066;
  assign n44774 = n44815 & n44816;
  assign n44746 = n44817 ^ n44818;
  assign n44845 = n44863 & n44864;
  assign n44733 = n44865 & n44866;
  assign n43383 = ~n44868;
  assign n44820 = ~n44869;
  assign n44847 = n44887 ^ n41980;
  assign n44761 = n44908 ^ n44909;
  assign n44888 = ~n44887;
  assign n44910 = ~n44909;
  assign n44959 = n44913 & n272;
  assign n44956 = ~n44981;
  assign n44958 = ~n44913;
  assign n44982 = n44999 & n45000;
  assign n44973 = ~n45001;
  assign n44935 = ~n45002;
  assign n43916 = ~n45003;
  assign n44983 = n41264 & n43935;
  assign n44998 = n45015 & n45016;
  assign n44976 = ~n45024;
  assign n45004 = n45047 & n45048;
  assign n44731 = n44774 ^ n44746;
  assign n44776 = n44774 & n7122;
  assign n44775 = ~n44774;
  assign n44823 = n44733 & n44778;
  assign n44819 = ~n44845;
  assign n44821 = ~n44733;
  assign n40715 = n44846 ^ n44847;
  assign n44871 = n44761 & n41920;
  assign n44872 = n44888 & n44889;
  assign n44870 = ~n44761;
  assign n44830 = n44910 & n44911;
  assign n44912 = n44956 & n44957;
  assign n44945 = n44958 & n10140;
  assign n44875 = ~n44959;
  assign n44806 = n44973 & n44974;
  assign n44895 = ~n44982;
  assign n43937 = ~n44983;
  assign n44975 = ~n44998;
  assign n44961 = n45004 ^ n42509;
  assign n45005 = ~n45004;
  assign n44692 = n416 ^ n44731;
  assign n44759 = n44775 & n416;
  assign n44745 = ~n44776;
  assign n44799 = n40715 & n43327;
  assign n44777 = n44819 & n44820;
  assign n44801 = n44821 & n44822;
  assign n44779 = ~n44823;
  assign n44802 = n40715 & n43241;
  assign n44803 = n40715 & n41980;
  assign n40738 = ~n40715;
  assign n44867 = n44870 & n41952;
  assign n44797 = ~n44871;
  assign n44842 = ~n44872;
  assign n44829 = ~n44830;
  assign n44873 = n44912 ^ n44913;
  assign n44914 = ~n44912;
  assign n44915 = ~n44945;
  assign n44937 = n44806 & n44946;
  assign n44936 = ~n44806;
  assign n41195 = n44960 ^ n44961;
  assign n44932 = n44975 & n44976;
  assign n44984 = n45005 & n45006;
  assign n43227 = n44691 ^ n44692;
  assign n44693 = ~n44692;
  assign n44732 = n44745 & n44746;
  assign n44705 = ~n44759;
  assign n44734 = n44777 ^ n44778;
  assign n43329 = ~n44799;
  assign n44787 = n40738 & n44800;
  assign n44780 = ~n44777;
  assign n44736 = ~n44801;
  assign n44781 = ~n44802;
  assign n43290 = ~n44803;
  assign n44804 = n44842 & n44843;
  assign n44764 = ~n44867;
  assign n44831 = n272 ^ n44873;
  assign n44903 = n44914 & n44915;
  assign n44890 = n44932 ^ n44933;
  assign n44917 = n44936 & n44851;
  assign n44918 = n41195 & n43830;
  assign n44853 = ~n44937;
  assign n44920 = n41195 & n43875;
  assign n44921 = n41195 & n42509;
  assign n41269 = ~n41195;
  assign n44934 = ~n44932;
  assign n44962 = ~n44984;
  assign n44558 = ~n43227;
  assign n44574 = n44693 & n44691;
  assign n44704 = ~n44732;
  assign n44664 = n44733 ^ n44734;
  assign n44760 = n44779 & n44780;
  assign n44648 = n44781 & n44782;
  assign n43347 = ~n44787;
  assign n44762 = n44804 ^ n41952;
  assign n44677 = n44830 ^ n44831;
  assign n44798 = ~n44804;
  assign n44828 = ~n44831;
  assign n44792 = n44890 ^ n44891;
  assign n44874 = ~n44903;
  assign n44809 = ~n44917;
  assign n44892 = ~n44918;
  assign n44904 = n41269 & n44919;
  assign n43877 = ~n44920;
  assign n43848 = ~n44921;
  assign n44916 = n44934 & n44935;
  assign n44922 = n44962 & n44963;
  assign n44573 = ~n44574;
  assign n44663 = n44704 & n44705;
  assign n44694 = n44664 & n7117;
  assign n44695 = ~n44664;
  assign n44738 = n44648 & n44747;
  assign n44735 = ~n44760;
  assign n44737 = ~n44648;
  assign n40685 = n44761 ^ n44762;
  assign n44790 = n44797 & n44798;
  assign n44788 = n44677 & n41905;
  assign n44789 = ~n44677;
  assign n44748 = n44828 & n44829;
  assign n44848 = n44792 & n10097;
  assign n44832 = n44874 & n44875;
  assign n44849 = ~n44792;
  assign n44727 = n44892 & n44893;
  assign n43897 = ~n44904;
  assign n44894 = ~n44916;
  assign n44876 = n44922 ^ n42536;
  assign n44923 = ~n44922;
  assign n44617 = n44663 ^ n44664;
  assign n44661 = ~n44663;
  assign n44662 = ~n44694;
  assign n44674 = n44695 & n431;
  assign n44719 = n40685 & n43308;
  assign n44696 = n44735 & n44736;
  assign n44717 = n44737 & n44697;
  assign n44698 = ~n44738;
  assign n44720 = n40685 & n43201;
  assign n44721 = n40685 & n41920;
  assign n40672 = ~n40685;
  assign n44679 = ~n44788;
  assign n44783 = n44789 & n41931;
  assign n44763 = ~n44790;
  assign n44751 = ~n44748;
  assign n44791 = n287 ^ n44832;
  assign n44824 = ~n44848;
  assign n44833 = n44849 & n287;
  assign n44825 = ~n44832;
  assign n44856 = n44727 & n44768;
  assign n44854 = ~n44727;
  assign n41110 = n44876 ^ n44877;
  assign n44850 = n44894 & n44895;
  assign n44905 = n44923 & n44924;
  assign n44575 = n431 ^ n44617;
  assign n44647 = n44661 & n44662;
  assign n44619 = ~n44674;
  assign n44649 = n44696 ^ n44697;
  assign n44645 = ~n44717;
  assign n44699 = ~n44696;
  assign n44706 = n40672 & n44718;
  assign n43287 = ~n44719;
  assign n44700 = ~n44720;
  assign n43245 = ~n44721;
  assign n44722 = n44763 & n44764;
  assign n44724 = ~n44783;
  assign n44749 = n44791 ^ n44792;
  assign n44805 = n44824 & n44825;
  assign n44785 = ~n44833;
  assign n44807 = n44850 ^ n44851;
  assign n44835 = n44854 & n44855;
  assign n44836 = n41110 & n43789;
  assign n44770 = ~n44856;
  assign n44837 = n41110 & n44857;
  assign n44838 = n41110 & n42536;
  assign n41198 = ~n41110;
  assign n44852 = ~n44850;
  assign n44878 = ~n44905;
  assign n43170 = n44574 ^ n44575;
  assign n44572 = ~n44575;
  assign n44618 = ~n44647;
  assign n44577 = n44648 ^ n44649;
  assign n44675 = n44698 & n44699;
  assign n44561 = n44700 & n44701;
  assign n43310 = ~n44706;
  assign n44676 = n44722 ^ n41931;
  assign n44723 = ~n44722;
  assign n44590 = n44748 ^ n44749;
  assign n44750 = ~n44749;
  assign n44784 = ~n44805;
  assign n44740 = n44806 ^ n44807;
  assign n44730 = ~n44835;
  assign n44810 = ~n44836;
  assign n44826 = n41198 & n43836;
  assign n43839 = ~n44837;
  assign n43807 = ~n44838;
  assign n44834 = n44852 & n44853;
  assign n44839 = n44878 & n44879;
  assign n44465 = ~n43170;
  assign n44493 = n44572 & n44573;
  assign n44576 = n44618 & n44619;
  assign n44609 = n44577 & n430;
  assign n44608 = ~n44577;
  assign n44652 = n44561 & n44611;
  assign n44644 = ~n44675;
  assign n44650 = ~n44561;
  assign n40636 = n44676 ^ n44677;
  assign n44707 = n44590 & n41871;
  assign n44709 = n44723 & n44724;
  assign n44708 = ~n44590;
  assign n44653 = n44750 & n44751;
  assign n44739 = n44784 & n44785;
  assign n44766 = n44740 & n286;
  assign n44765 = ~n44740;
  assign n44638 = n44810 & n44811;
  assign n43861 = ~n44826;
  assign n44808 = ~n44834;
  assign n44794 = n44839 ^ n42513;
  assign n44840 = ~n44839;
  assign n44496 = ~n44493;
  assign n44532 = n44576 ^ n44577;
  assign n44560 = ~n44576;
  assign n44588 = n44608 & n7047;
  assign n44519 = ~n44609;
  assign n44610 = n44644 & n44645;
  assign n44627 = n40636 & n44646;
  assign n44628 = n44650 & n44651;
  assign n44629 = n40636 & n43187;
  assign n44613 = ~n44652;
  assign n44630 = n40636 & n41931;
  assign n40661 = ~n40636;
  assign n44633 = ~n44707;
  assign n44702 = n44708 & n41862;
  assign n44678 = ~n44709;
  assign n44656 = ~n44653;
  assign n44703 = n44739 ^ n44740;
  assign n44726 = ~n44739;
  assign n44752 = n44765 & n10065;
  assign n44681 = ~n44766;
  assign n44772 = n44638 & n44786;
  assign n44771 = ~n44638;
  assign n41029 = n44793 ^ n44794;
  assign n44767 = n44808 & n44809;
  assign n44827 = n44840 & n44841;
  assign n44494 = n430 ^ n44532;
  assign n44559 = ~n44588;
  assign n44562 = n44610 ^ n44611;
  assign n43249 = ~n44627;
  assign n44620 = n40661 & n43247;
  assign n44612 = ~n44610;
  assign n44564 = ~n44628;
  assign n44606 = ~n44629;
  assign n43205 = ~n44630;
  assign n44631 = n44678 & n44679;
  assign n44594 = ~n44702;
  assign n44654 = n286 ^ n44703;
  assign n44725 = ~n44752;
  assign n44728 = n44767 ^ n44768;
  assign n44754 = n44771 & n44685;
  assign n44687 = ~n44772;
  assign n44755 = n41029 & n44773;
  assign n41114 = ~n41029;
  assign n44769 = ~n44767;
  assign n44795 = ~n44827;
  assign n43127 = n44493 ^ n44494;
  assign n44495 = ~n44494;
  assign n44541 = n44559 & n44560;
  assign n44483 = n44561 ^ n44562;
  assign n44484 = n44606 & n44607;
  assign n44589 = n44612 & n44613;
  assign n43266 = ~n44620;
  assign n44591 = n44631 ^ n41862;
  assign n44497 = n44653 ^ n44654;
  assign n44632 = ~n44631;
  assign n44655 = ~n44654;
  assign n44710 = n44725 & n44726;
  assign n44635 = n44727 ^ n44728;
  assign n44641 = ~n44754;
  assign n44741 = n41114 & n43709;
  assign n44742 = n41114 & n43796;
  assign n43819 = ~n44755;
  assign n44743 = n41114 & n42439;
  assign n44753 = n44769 & n44770;
  assign n44756 = n44795 & n44796;
  assign n44396 = ~n43127;
  assign n44418 = n44495 & n44496;
  assign n44520 = n44483 & n7015;
  assign n44518 = ~n44541;
  assign n44521 = ~n44483;
  assign n44567 = n44484 & n44523;
  assign n44565 = ~n44484;
  assign n44563 = ~n44589;
  assign n40602 = n44590 ^ n44591;
  assign n44615 = n44497 & n41829;
  assign n44614 = ~n44497;
  assign n44621 = n44632 & n44633;
  assign n44546 = n44655 & n44656;
  assign n44682 = n44635 & n10044;
  assign n44680 = ~n44710;
  assign n44683 = ~n44635;
  assign n44711 = ~n44741;
  assign n43799 = ~n44742;
  assign n43763 = ~n44743;
  assign n44729 = ~n44753;
  assign n44714 = n44756 ^ n42386;
  assign n44757 = ~n44756;
  assign n44482 = n44518 & n44519;
  assign n44480 = ~n44520;
  assign n44506 = n44521 & n429;
  assign n44544 = n40602 & n43124;
  assign n44542 = n40602 & n44558;
  assign n44522 = n44563 & n44564;
  assign n44543 = n44565 & n44566;
  assign n44525 = ~n44567;
  assign n44545 = n40602 & n41871;
  assign n40607 = ~n40602;
  assign n44592 = n44614 & n41804;
  assign n44505 = ~n44615;
  assign n44593 = ~n44621;
  assign n44549 = ~n44546;
  assign n44634 = n44680 & n44681;
  assign n44637 = ~n44682;
  assign n44665 = n44683 & n285;
  assign n44688 = n44711 & n44712;
  assign n40957 = n44713 ^ n44714;
  assign n44684 = n44729 & n44730;
  assign n44744 = n44757 & n44758;
  assign n44449 = n44482 ^ n44483;
  assign n44481 = ~n44482;
  assign n44452 = ~n44506;
  assign n44485 = n44522 ^ n44523;
  assign n44533 = n40607 & n43227;
  assign n43209 = ~n44542;
  assign n44524 = ~n44522;
  assign n44487 = ~n44543;
  assign n44526 = ~n44544;
  assign n43169 = ~n44545;
  assign n44540 = ~n44592;
  assign n44578 = n44593 & n44594;
  assign n44595 = n44634 ^ n44635;
  assign n44636 = ~n44634;
  assign n44597 = ~n44665;
  assign n44639 = n44684 ^ n44685;
  assign n44669 = n44688 & n44689;
  assign n44671 = n40957 & n43777;
  assign n44667 = ~n44688;
  assign n41033 = ~n40957;
  assign n44686 = ~n44684;
  assign n44715 = ~n44744;
  assign n44419 = n429 ^ n44449;
  assign n44466 = n44480 & n44481;
  assign n44421 = n44484 ^ n44485;
  assign n44507 = n44524 & n44525;
  assign n44424 = n44526 & n44527;
  assign n43229 = ~n44533;
  assign n44535 = ~n44578;
  assign n44547 = n285 ^ n44595;
  assign n44622 = n44636 & n44637;
  assign n44616 = n44638 ^ n44639;
  assign n44657 = n44667 & n44668;
  assign n44601 = ~n44669;
  assign n44658 = n41033 & n44670;
  assign n43779 = ~n44671;
  assign n44659 = n41033 & n42443;
  assign n44660 = n41033 & n43698;
  assign n44666 = n44686 & n44687;
  assign n44672 = n44715 & n44716;
  assign n43086 = n44418 ^ n44419;
  assign n44349 = n44419 & n44418;
  assign n44453 = n44421 & n6946;
  assign n44451 = ~n44466;
  assign n44448 = ~n44421;
  assign n44490 = n44424 & n44455;
  assign n44486 = ~n44507;
  assign n44488 = ~n44424;
  assign n44498 = n44535 ^ n41829;
  assign n44534 = n44535 & n44540;
  assign n44432 = n44546 ^ n44547;
  assign n44548 = ~n44547;
  assign n44599 = n44616 & n284;
  assign n44596 = ~n44622;
  assign n44598 = ~n44616;
  assign n44553 = ~n44657;
  assign n43758 = ~n44658;
  assign n43716 = ~n44659;
  assign n44623 = ~n44660;
  assign n44640 = ~n44666;
  assign n44626 = n44672 ^ n42333;
  assign n44673 = n44672 & n44690;
  assign n44353 = ~n43086;
  assign n44352 = ~n44349;
  assign n44431 = n44448 & n428;
  assign n44420 = n44451 & n44452;
  assign n44423 = ~n44453;
  assign n44454 = n44486 & n44487;
  assign n44467 = n44488 & n44489;
  assign n44457 = ~n44490;
  assign n40552 = n44497 ^ n44498;
  assign n44508 = n44432 & n41801;
  assign n44504 = ~n44534;
  assign n44509 = ~n44432;
  assign n44462 = n44548 & n44549;
  assign n44500 = n44596 & n44597;
  assign n44579 = n44598 & n9976;
  assign n44511 = ~n44599;
  assign n44476 = n44623 & n44624;
  assign n44580 = n44553 & n44601;
  assign n40961 = n44625 ^ n44626;
  assign n44581 = n44640 & n44641;
  assign n44642 = ~n44673;
  assign n44379 = n44420 ^ n44421;
  assign n44422 = ~n44420;
  assign n44381 = ~n44431;
  assign n44425 = n44454 ^ n44455;
  assign n44459 = n40552 & n43113;
  assign n44458 = n40552 & n44465;
  assign n44456 = ~n44454;
  assign n44417 = ~n44467;
  assign n44460 = n40552 & n41804;
  assign n40573 = ~n40552;
  assign n44468 = n44504 & n44505;
  assign n44469 = ~n44508;
  assign n44499 = n44509 & n41772;
  assign n44471 = ~n44462;
  assign n44550 = ~n44500;
  assign n44551 = ~n44579;
  assign n44473 = n44580 ^ n44581;
  assign n44584 = n40961 & n42393;
  assign n44585 = n44476 & n44602;
  assign n44586 = n40961 & n43642;
  assign n44587 = n40961 & n44603;
  assign n44583 = ~n44476;
  assign n40884 = ~n40961;
  assign n44600 = ~n44581;
  assign n44604 = n44642 & n44643;
  assign n44350 = n428 ^ n44379;
  assign n44397 = n44422 & n44423;
  assign n44355 = n44424 ^ n44425;
  assign n44436 = n44456 & n44457;
  assign n44450 = n40573 & n43170;
  assign n43173 = ~n44458;
  assign n44434 = ~n44459;
  assign n43132 = ~n44460;
  assign n44433 = n44468 ^ n41772;
  assign n44470 = ~n44468;
  assign n44438 = ~n44499;
  assign n44536 = n44550 & n44551;
  assign n44537 = n44551 & n44511;
  assign n44538 = n44473 & n9936;
  assign n44539 = ~n44473;
  assign n44568 = n44583 & n44513;
  assign n43680 = ~n44584;
  assign n44515 = ~n44585;
  assign n44554 = ~n44586;
  assign n44571 = n40884 & n43717;
  assign n43720 = ~n44587;
  assign n44582 = n44600 & n44601;
  assign n43668 = n44604 ^ n44605;
  assign n44293 = n44349 ^ n44350;
  assign n44351 = ~n44350;
  assign n44382 = n44355 & n6920;
  assign n44380 = ~n44397;
  assign n44383 = ~n44355;
  assign n40523 = n44432 ^ n44433;
  assign n44347 = n44434 & n44435;
  assign n44416 = ~n44436;
  assign n43191 = ~n44450;
  assign n44461 = n44469 & n44470;
  assign n44510 = ~n44536;
  assign n44501 = ~n44537;
  assign n44475 = ~n44538;
  assign n44529 = n44539 & n283;
  assign n44412 = n44554 & n44555;
  assign n44479 = ~n44568;
  assign n44556 = n43668 & n44569;
  assign n44557 = n43668 & n44570;
  assign n43737 = ~n44571;
  assign n44552 = ~n44582;
  assign n40933 = ~n43668;
  assign n44279 = ~n44293;
  assign n44291 = n44351 & n44352;
  assign n44354 = n44380 & n44381;
  assign n44356 = ~n44382;
  assign n44365 = n44383 & n427;
  assign n44402 = n44347 & n44387;
  assign n44386 = n44416 & n44417;
  assign n44398 = n40523 & n43038;
  assign n44395 = n40523 & n43127;
  assign n44399 = n40523 & n41801;
  assign n44400 = ~n44347;
  assign n40520 = ~n40523;
  assign n44437 = ~n44461;
  assign n44463 = n44500 ^ n44501;
  assign n44472 = n44510 & n44511;
  assign n44517 = n44412 & n44528;
  assign n44441 = ~n44529;
  assign n44516 = ~n44412;
  assign n44512 = n44552 & n44553;
  assign n44530 = ~n44556;
  assign n43651 = ~n44557;
  assign n44304 = ~n44291;
  assign n44319 = n44354 ^ n44355;
  assign n44357 = ~n44354;
  assign n44321 = ~n44365;
  assign n44348 = n44386 ^ n44387;
  assign n43130 = ~n44395;
  assign n44391 = n40520 & n44396;
  assign n44384 = ~n44398;
  assign n43085 = ~n44399;
  assign n44388 = ~n44386;
  assign n44392 = n44400 & n44401;
  assign n44389 = ~n44402;
  assign n44403 = n44437 & n44438;
  assign n44366 = n44462 ^ n44463;
  assign n44406 = n44463 & n44471;
  assign n44439 = n44472 ^ n44473;
  assign n44474 = ~n44472;
  assign n44477 = n44512 ^ n44513;
  assign n44503 = n44516 & n44445;
  assign n44447 = ~n44517;
  assign n44491 = n44530 & n44531;
  assign n44514 = ~n44512;
  assign n44292 = n427 ^ n44319;
  assign n44295 = n44347 ^ n44348;
  assign n44334 = n44356 & n44357;
  assign n44298 = n44384 & n44385;
  assign n44368 = n44388 & n44389;
  assign n43155 = ~n44391;
  assign n44361 = ~n44392;
  assign n44367 = n44403 ^ n41732;
  assign n44404 = ~n44403;
  assign n44428 = n44366 & n41732;
  assign n44407 = n283 ^ n44439;
  assign n44427 = ~n44366;
  assign n44464 = n44474 & n44475;
  assign n44409 = n44476 ^ n44477;
  assign n44346 = n44491 ^ n44492;
  assign n44415 = ~n44503;
  assign n44502 = n44514 & n44515;
  assign n43020 = n44291 ^ n44292;
  assign n44240 = n44292 & n44304;
  assign n44322 = n44295 & n6878;
  assign n44320 = ~n44334;
  assign n44323 = ~n44295;
  assign n44359 = n44298 & n44362;
  assign n44358 = ~n44298;
  assign n40467 = n44366 ^ n44367;
  assign n44360 = ~n44368;
  assign n44390 = n44406 ^ n44407;
  assign n44338 = n44407 & n44406;
  assign n44426 = n44427 & n41756;
  assign n44405 = ~n44428;
  assign n44443 = n44409 & n282;
  assign n44440 = ~n44464;
  assign n44442 = ~n44409;
  assign n44478 = ~n44502;
  assign n44244 = ~n43020;
  assign n44243 = ~n44240;
  assign n44294 = n44320 & n44321;
  assign n44297 = ~n44322;
  assign n44306 = n44323 & n426;
  assign n44333 = n40467 & n44353;
  assign n44335 = n44358 & n44327;
  assign n44325 = ~n44359;
  assign n44326 = n44360 & n44361;
  assign n40489 = ~n40467;
  assign n44372 = n44390 & n41713;
  assign n44371 = ~n44390;
  assign n44393 = n44404 & n44405;
  assign n44370 = ~n44426;
  assign n44408 = n44440 & n44441;
  assign n44429 = n44442 & n9908;
  assign n44375 = ~n44443;
  assign n44444 = n44478 & n44479;
  assign n44264 = n44294 ^ n44295;
  assign n44296 = ~n44294;
  assign n44266 = ~n44306;
  assign n44299 = n44326 ^ n44327;
  assign n44328 = n40489 & n43086;
  assign n43111 = ~n44333;
  assign n44301 = ~n44335;
  assign n44329 = n40489 & n41732;
  assign n44330 = n40489 & n43024;
  assign n44324 = ~n44326;
  assign n44363 = n44371 & n41674;
  assign n44313 = ~n44372;
  assign n44369 = ~n44393;
  assign n44373 = n44408 ^ n44409;
  assign n44411 = ~n44408;
  assign n44410 = ~n44429;
  assign n44413 = n44444 ^ n44445;
  assign n44446 = ~n44444;
  assign n44241 = n426 ^ n44264;
  assign n44281 = n44296 & n44297;
  assign n44246 = n44298 ^ n44299;
  assign n44309 = n44324 & n44325;
  assign n43089 = ~n44328;
  assign n43047 = ~n44329;
  assign n44307 = ~n44330;
  assign n44337 = ~n44363;
  assign n44311 = n44369 & n44370;
  assign n44339 = n282 ^ n44373;
  assign n44394 = n44410 & n44411;
  assign n44342 = n44412 ^ n44413;
  assign n44430 = n44446 & n44447;
  assign n44193 = n44240 ^ n44241;
  assign n44242 = ~n44241;
  assign n44268 = n44246 & n425;
  assign n44265 = ~n44281;
  assign n44267 = ~n44246;
  assign n44247 = n44307 & n44308;
  assign n44300 = ~n44309;
  assign n44310 = n44337 & n44313;
  assign n44286 = n44338 ^ n44339;
  assign n44336 = ~n44311;
  assign n44340 = ~n44339;
  assign n44377 = n44342 & n281;
  assign n44374 = ~n44394;
  assign n44376 = ~n44342;
  assign n44414 = ~n44430;
  assign n42962 = ~n44193;
  assign n44197 = n44242 & n44243;
  assign n44245 = n44265 & n44266;
  assign n44256 = n44267 & n6844;
  assign n44219 = ~n44268;
  assign n44269 = n44300 & n44301;
  assign n44283 = n44247 & n44302;
  assign n44282 = ~n44247;
  assign n40399 = n44310 ^ n44311;
  assign n44315 = n44286 & n41666;
  assign n44314 = ~n44286;
  assign n44331 = n44336 & n44337;
  assign n44289 = n44340 & n44338;
  assign n44341 = n44374 & n44375;
  assign n44364 = n44376 & n9894;
  assign n44318 = ~n44377;
  assign n44378 = n44414 & n44415;
  assign n44215 = n44245 ^ n44246;
  assign n44249 = ~n44245;
  assign n44250 = ~n44256;
  assign n44248 = n44269 ^ n44270;
  assign n44272 = ~n44269;
  assign n44276 = n44282 & n44270;
  assign n44271 = ~n44283;
  assign n44280 = n40399 & n44293;
  assign n44284 = n40399 & n41674;
  assign n40454 = ~n40399;
  assign n44305 = n44314 & n41654;
  assign n44288 = ~n44315;
  assign n44312 = ~n44331;
  assign n44303 = ~n44289;
  assign n44316 = n44341 ^ n44342;
  assign n44343 = ~n44341;
  assign n44344 = ~n44364;
  assign n44345 = n280 ^ n44378;
  assign n44198 = n425 ^ n44215;
  assign n44204 = n44247 ^ n44248;
  assign n44233 = n44249 & n44250;
  assign n44257 = n44271 & n44272;
  assign n44252 = ~n44276;
  assign n44275 = n40454 & n44279;
  assign n43071 = ~n44280;
  assign n44277 = n40454 & n42959;
  assign n43027 = ~n44284;
  assign n44263 = ~n44305;
  assign n44285 = n44312 & n44313;
  assign n44290 = n281 ^ n44316;
  assign n44332 = n44343 & n44344;
  assign n44255 = n44345 ^ n44346;
  assign n44152 = n44197 ^ n44198;
  assign n44156 = n44198 & n44197;
  assign n44217 = n44204 & n424;
  assign n44216 = ~n44204;
  assign n44218 = ~n44233;
  assign n44251 = ~n44257;
  assign n43045 = ~n44275;
  assign n44259 = ~n44277;
  assign n44258 = n44285 ^ n44286;
  assign n44211 = n44289 ^ n44290;
  assign n44274 = n44290 & n44303;
  assign n44287 = ~n44285;
  assign n44317 = ~n44332;
  assign n42919 = ~n44152;
  assign n44209 = n44216 & n6815;
  assign n44177 = ~n44217;
  assign n44203 = n44218 & n44219;
  assign n44220 = n44251 & n44252;
  assign n43068 = n43071 & n43045;
  assign n40410 = n44258 ^ n41654;
  assign n44221 = n44259 & n44260;
  assign n44261 = n44258 & n41666;
  assign n44278 = n44287 & n44288;
  assign n44273 = n44317 & n44318;
  assign n44178 = n44203 ^ n44204;
  assign n44200 = ~n44209;
  assign n44199 = ~n44203;
  assign n44201 = n44220 ^ n44221;
  assign n44222 = ~n44220;
  assign n44232 = n40410 & n44244;
  assign n44234 = n40410 & n42883;
  assign n44236 = n44221 & n44253;
  assign n40376 = ~n40410;
  assign n44235 = ~n44221;
  assign n42968 = ~n44261;
  assign n44254 = n44273 ^ n44274;
  assign n44262 = ~n44278;
  assign n44157 = n424 ^ n44178;
  assign n44194 = n44199 & n44200;
  assign n44142 = n44201 ^ n44202;
  assign n43004 = ~n44232;
  assign n44229 = n40376 & n43020;
  assign n44224 = ~n44234;
  assign n44230 = n44235 & n44202;
  assign n44223 = ~n44236;
  assign n44167 = n44254 ^ n44255;
  assign n44237 = n44262 & n44263;
  assign n44085 = n44156 ^ n44157;
  assign n44120 = n44157 & n44156;
  assign n44180 = n44142 & n439;
  assign n44176 = ~n44194;
  assign n44179 = ~n44142;
  assign n44210 = n44222 & n44223;
  assign n44181 = n44224 & n44225;
  assign n43022 = ~n44229;
  assign n44226 = n44167 & n41605;
  assign n44206 = ~n44230;
  assign n44227 = ~n44167;
  assign n44212 = n44237 ^ n41602;
  assign n44239 = n44237 & n41602;
  assign n44238 = ~n44237;
  assign n42879 = ~n44085;
  assign n44158 = n44176 & n44177;
  assign n44173 = n44179 & n6709;
  assign n44144 = ~n44180;
  assign n44205 = ~n44210;
  assign n44171 = ~n44181;
  assign n40330 = n44211 ^ n44212;
  assign n44189 = ~n44226;
  assign n44213 = n44227 & n41563;
  assign n44231 = n44238 & n41643;
  assign n44228 = ~n44239;
  assign n44141 = n439 ^ n44158;
  assign n44160 = ~n44158;
  assign n44159 = ~n44173;
  assign n44192 = n40330 & n42962;
  assign n44182 = n44205 & n44206;
  assign n44195 = n40330 & n42867;
  assign n44196 = n40330 & n41602;
  assign n40345 = ~n40330;
  assign n44169 = ~n44213;
  assign n44214 = n44228 & n44211;
  assign n44208 = ~n44231;
  assign n44121 = n44141 ^ n44142;
  assign n44154 = n44159 & n44160;
  assign n44161 = n44181 ^ n44182;
  assign n44186 = n44182 & n44191;
  assign n42964 = ~n44192;
  assign n44190 = n40345 & n44193;
  assign n44185 = ~n44182;
  assign n44183 = ~n44195;
  assign n42926 = ~n44196;
  assign n44207 = ~n44214;
  assign n42838 = n44120 ^ n44121;
  assign n44088 = n44121 & n44120;
  assign n44143 = ~n44154;
  assign n44123 = n44161 ^ n44162;
  assign n44111 = n44183 & n44184;
  assign n44174 = n44185 & n44162;
  assign n44170 = ~n44186;
  assign n42988 = ~n44190;
  assign n44187 = n44207 & n44208;
  assign n44058 = ~n42838;
  assign n44122 = n44143 & n44144;
  assign n44146 = n44123 & n438;
  assign n44145 = ~n44123;
  assign n44163 = n44170 & n44171;
  assign n44165 = n44111 & n44172;
  assign n44164 = ~n44111;
  assign n44151 = ~n44174;
  assign n44166 = n44187 ^ n41605;
  assign n44188 = ~n44187;
  assign n44106 = n44122 ^ n44123;
  assign n44125 = ~n44122;
  assign n44136 = n44145 & n6678;
  assign n44108 = ~n44146;
  assign n44150 = ~n44163;
  assign n44155 = n44164 & n44132;
  assign n44134 = ~n44165;
  assign n40250 = n44166 ^ n44167;
  assign n44175 = n44188 & n44189;
  assign n44089 = n438 ^ n44106;
  assign n44124 = ~n44136;
  assign n44131 = n44150 & n44151;
  assign n44147 = n40250 & n44152;
  assign n44114 = ~n44155;
  assign n40315 = ~n40250;
  assign n44168 = ~n44175;
  assign n42801 = n44088 ^ n44089;
  assign n44043 = n44089 & n44088;
  assign n44118 = n44124 & n44125;
  assign n44112 = n44131 ^ n44132;
  assign n42946 = ~n44147;
  assign n44137 = n40315 & n42919;
  assign n44133 = ~n44131;
  assign n44138 = n40315 & n42827;
  assign n44139 = n40315 & n41605;
  assign n44153 = n44168 & n44169;
  assign n44025 = ~n42801;
  assign n44047 = ~n44043;
  assign n44083 = n44111 ^ n44112;
  assign n44107 = ~n44118;
  assign n44128 = n44133 & n44134;
  assign n42922 = ~n44137;
  assign n44126 = ~n44138;
  assign n42887 = ~n44139;
  assign n44149 = n44153 & n41566;
  assign n44148 = ~n44153;
  assign n44094 = n44083 & n437;
  assign n44102 = n44107 & n44108;
  assign n44093 = ~n44083;
  assign n44074 = n44126 & n44127;
  assign n44113 = ~n44128;
  assign n44140 = n44148 & n41524;
  assign n44130 = ~n44149;
  assign n44090 = n44093 & n6625;
  assign n44056 = ~n44094;
  assign n44073 = ~n44102;
  assign n44095 = n44113 & n44114;
  assign n44110 = n44074 & n44115;
  assign n44109 = ~n44074;
  assign n44129 = n44130 & n44135;
  assign n44117 = ~n44140;
  assign n44068 = n44073 ^ n44083;
  assign n44072 = ~n44090;
  assign n44075 = n44095 ^ n44096;
  assign n44097 = ~n44095;
  assign n44103 = n44109 & n44096;
  assign n44098 = ~n44110;
  assign n44116 = ~n44129;
  assign n44119 = n44117 & n44130;
  assign n44044 = n437 ^ n44068;
  assign n44069 = n44072 & n44073;
  assign n44031 = n44074 ^ n44075;
  assign n44091 = n44097 & n44098;
  assign n44077 = ~n44103;
  assign n44099 = n44116 & n44117;
  assign n44104 = ~n44119;
  assign n42758 = n44043 ^ n44044;
  assign n43990 = n44044 & n44047;
  assign n44057 = n44031 & n436;
  assign n44055 = ~n44069;
  assign n44054 = ~n44031;
  assign n44076 = ~n44091;
  assign n44079 = n44099 ^ n41515;
  assign n40187 = n44104 ^ n44105;
  assign n44100 = ~n44099;
  assign n43976 = ~n42758;
  assign n44048 = n44054 & n6577;
  assign n44030 = n44055 & n44056;
  assign n44014 = ~n44057;
  assign n44060 = n44076 & n44077;
  assign n40109 = n44079 ^ n44080;
  assign n44084 = n40187 & n42879;
  assign n44086 = n40187 & n42788;
  assign n44087 = n40187 & n41566;
  assign n44092 = n44100 & n44101;
  assign n40261 = ~n40187;
  assign n44012 = n44030 ^ n44031;
  assign n44033 = ~n44030;
  assign n44032 = ~n44048;
  assign n44035 = n44060 ^ n44061;
  assign n44059 = n40109 & n42838;
  assign n44064 = n44060 & n44061;
  assign n44062 = ~n44060;
  assign n40169 = ~n40109;
  assign n42881 = ~n44084;
  assign n44078 = n40261 & n44085;
  assign n44070 = ~n44086;
  assign n42847 = ~n44087;
  assign n44081 = ~n44092;
  assign n43991 = n436 ^ n44012;
  assign n44029 = n44032 & n44033;
  assign n44049 = n40169 & n44058;
  assign n42863 = ~n44059;
  assign n44050 = n44062 & n44063;
  assign n44051 = n40169 & n42777;
  assign n44045 = ~n44064;
  assign n44052 = n40169 & n41483;
  assign n44034 = n44070 & n44071;
  assign n42906 = ~n44078;
  assign n44065 = n44081 & n44082;
  assign n42738 = n43990 ^ n43991;
  assign n43992 = ~n43991;
  assign n44013 = ~n44029;
  assign n43994 = n44034 ^ n44035;
  assign n42841 = ~n44049;
  assign n44027 = ~n44050;
  assign n44036 = ~n44051;
  assign n42800 = ~n44052;
  assign n44039 = n44065 ^ n41486;
  assign n44046 = ~n44034;
  assign n44066 = ~n44065;
  assign n43960 = ~n42738;
  assign n43949 = n43992 & n43990;
  assign n43993 = n44013 & n44014;
  assign n44015 = n43994 & n6508;
  assign n44016 = ~n43994;
  assign n43982 = n44036 & n44037;
  assign n40044 = n44039 ^ n44040;
  assign n44038 = n44045 & n44046;
  assign n44053 = n44066 & n44067;
  assign n43972 = n43993 ^ n43994;
  assign n43996 = ~n43993;
  assign n43995 = ~n44015;
  assign n44008 = n44016 & n435;
  assign n44017 = n40044 & n44025;
  assign n44019 = n43982 & n44028;
  assign n44020 = n40044 & n42748;
  assign n44021 = n40044 & n41486;
  assign n44018 = ~n43982;
  assign n40122 = ~n40044;
  assign n44026 = ~n44038;
  assign n44041 = ~n44053;
  assign n43950 = n435 ^ n43972;
  assign n43988 = n43995 & n43996;
  assign n43974 = ~n44008;
  assign n42804 = ~n44017;
  assign n44009 = n40122 & n42801;
  assign n44010 = n44018 & n44003;
  assign n44007 = ~n44019;
  assign n44004 = ~n44020;
  assign n42767 = ~n44021;
  assign n44002 = n44026 & n44027;
  assign n44022 = n44041 & n44042;
  assign n42677 = n43949 ^ n43950;
  assign n43906 = n43950 & n43949;
  assign n43973 = ~n43988;
  assign n43983 = n44002 ^ n44003;
  assign n43940 = n44004 & n44005;
  assign n42823 = ~n44009;
  assign n43985 = ~n44010;
  assign n44006 = ~n44002;
  assign n43999 = n44022 ^ n41443;
  assign n44023 = ~n44022;
  assign n43892 = ~n42677;
  assign n43909 = ~n43906;
  assign n43967 = n43973 & n43974;
  assign n43948 = n43982 ^ n43983;
  assign n43987 = n43940 & n43989;
  assign n43986 = ~n43940;
  assign n39963 = n43998 ^ n43999;
  assign n43997 = n44006 & n44007;
  assign n44011 = n44023 & n44024;
  assign n43939 = ~n43967;
  assign n43962 = n43948 & n434;
  assign n43961 = ~n43948;
  assign n43975 = n39963 & n42758;
  assign n43977 = n43986 & n43964;
  assign n43966 = ~n43987;
  assign n39967 = ~n39963;
  assign n43984 = ~n43997;
  assign n44000 = ~n44011;
  assign n43927 = n43939 ^ n43948;
  assign n43952 = n43961 & n6432;
  assign n43918 = ~n43962;
  assign n42784 = ~n43975;
  assign n43968 = n39967 & n43976;
  assign n43943 = ~n43977;
  assign n43969 = n39967 & n42695;
  assign n43970 = n39967 & n41443;
  assign n43963 = n43984 & n43985;
  assign n43978 = n44000 & n44001;
  assign n43907 = n434 ^ n43927;
  assign n43938 = ~n43952;
  assign n43941 = n43963 ^ n43964;
  assign n42761 = ~n43968;
  assign n43953 = ~n43969;
  assign n42717 = ~n43970;
  assign n43965 = ~n43963;
  assign n39965 = n43978 ^ n43979;
  assign n43980 = ~n43978;
  assign n43855 = n43906 ^ n43907;
  assign n43908 = ~n43907;
  assign n43931 = n43938 & n43939;
  assign n43901 = n43940 ^ n43941;
  assign n43904 = n43953 & n43954;
  assign n43951 = n39965 & n43960;
  assign n43955 = n43965 & n43966;
  assign n43956 = n39965 & n42595;
  assign n43957 = n39965 & n41290;
  assign n39821 = ~n39965;
  assign n43971 = n43980 & n43981;
  assign n42634 = ~n43855;
  assign n43862 = n43908 & n43909;
  assign n43920 = n43901 & n433;
  assign n43917 = ~n43931;
  assign n43919 = ~n43901;
  assign n43933 = n43904 & n43944;
  assign n43932 = ~n43904;
  assign n42721 = ~n43951;
  assign n43947 = n39821 & n42738;
  assign n43942 = ~n43955;
  assign n43945 = ~n43956;
  assign n42685 = ~n43957;
  assign n43958 = ~n43971;
  assign n43900 = n43917 & n43918;
  assign n43910 = n43919 & n6316;
  assign n43880 = ~n43920;
  assign n43928 = n43932 & n43922;
  assign n43924 = ~n43933;
  assign n43921 = n43942 & n43943;
  assign n43884 = n43945 & n43946;
  assign n42740 = ~n43947;
  assign n43934 = n43958 & n43959;
  assign n43878 = n43900 ^ n43901;
  assign n43903 = ~n43900;
  assign n43902 = ~n43910;
  assign n43905 = n43921 ^ n43922;
  assign n43899 = ~n43928;
  assign n43926 = n43884 & n43929;
  assign n43923 = ~n43921;
  assign n43925 = ~n43884;
  assign n43912 = n43934 ^ n43935;
  assign n43936 = ~n43934;
  assign n43863 = n433 ^ n43878;
  assign n43893 = n43902 & n43903;
  assign n43865 = n43904 ^ n43905;
  assign n39781 = n43912 ^ n41327;
  assign n43911 = n43923 & n43924;
  assign n43913 = n43925 & n43869;
  assign n43886 = ~n43926;
  assign n43914 = n43912 & n41264;
  assign n43930 = n43936 & n43937;
  assign n42591 = n43862 ^ n43863;
  assign n43820 = n43863 & n43862;
  assign n43882 = n43865 & n432;
  assign n43879 = ~n43893;
  assign n43881 = ~n43865;
  assign n43891 = n39781 & n42677;
  assign n43894 = n39781 & n42622;
  assign n39791 = ~n39781;
  assign n43898 = ~n43911;
  assign n43871 = ~n43913;
  assign n42642 = ~n43914;
  assign n43915 = ~n43930;
  assign n43824 = ~n42591;
  assign n43864 = n43879 & n43880;
  assign n43872 = n43881 & n6292;
  assign n43842 = ~n43882;
  assign n42679 = ~n43891;
  assign n43889 = n39791 & n43892;
  assign n43887 = ~n43894;
  assign n43883 = n43898 & n43899;
  assign n43895 = n43915 & n43916;
  assign n43840 = n43864 ^ n43865;
  assign n43867 = ~n43864;
  assign n43866 = ~n43872;
  assign n43868 = n43883 ^ n43884;
  assign n43826 = n43887 & n43888;
  assign n42702 = ~n43889;
  assign n43885 = ~n43883;
  assign n43874 = n43895 ^ n41269;
  assign n43896 = ~n43895;
  assign n43821 = n432 ^ n43840;
  assign n43856 = n43866 & n43867;
  assign n43801 = n43868 ^ n43869;
  assign n43833 = ~n43826;
  assign n39673 = n43874 ^ n43875;
  assign n43873 = n43885 & n43886;
  assign n43890 = n43896 & n43897;
  assign n43770 = n43820 ^ n43821;
  assign n43780 = n43821 & n43820;
  assign n43844 = n43801 & n447;
  assign n43841 = ~n43856;
  assign n43843 = ~n43801;
  assign n43854 = n39673 & n42634;
  assign n43857 = n39673 & n42582;
  assign n43858 = n39673 & n41269;
  assign n39824 = ~n39673;
  assign n43870 = ~n43873;
  assign n43876 = ~n43890;
  assign n43782 = ~n43770;
  assign n43825 = n43841 & n43842;
  assign n43834 = n43843 & n6169;
  assign n43803 = ~n43844;
  assign n42636 = ~n43854;
  assign n43851 = n39824 & n43855;
  assign n43847 = ~n43857;
  assign n42599 = ~n43858;
  assign n43845 = n43870 & n43871;
  assign n43859 = n43876 & n43877;
  assign n43800 = n447 ^ n43825;
  assign n43822 = ~n43825;
  assign n43823 = ~n43834;
  assign n43827 = n43845 ^ n43846;
  assign n43765 = n43847 & n43848;
  assign n42656 = ~n43851;
  assign n43850 = n43845 & n43852;
  assign n43849 = ~n43845;
  assign n43837 = n43859 ^ n41110;
  assign n43860 = ~n43859;
  assign n43781 = n43800 ^ n43801;
  assign n43813 = n43822 & n43823;
  assign n43784 = n43826 ^ n43827;
  assign n43831 = n43765 & n43792;
  assign n43829 = ~n43765;
  assign n39600 = n43836 ^ n43837;
  assign n43835 = n43849 & n43846;
  assign n43832 = ~n43850;
  assign n43853 = n43860 & n43861;
  assign n42503 = n43780 ^ n43781;
  assign n43738 = n43781 & n43780;
  assign n43805 = n43784 & n446;
  assign n43802 = ~n43813;
  assign n43804 = ~n43784;
  assign n43812 = n39600 & n43824;
  assign n43814 = n43829 & n43830;
  assign n43815 = n39600 & n42489;
  assign n43794 = ~n43831;
  assign n43816 = n39600 & n41198;
  assign n43828 = n43832 & n43833;
  assign n39734 = ~n39600;
  assign n43810 = ~n43835;
  assign n43838 = ~n43853;
  assign n43730 = ~n42503;
  assign n43741 = ~n43738;
  assign n43783 = n43802 & n43803;
  assign n43795 = n43804 & n6144;
  assign n43760 = ~n43805;
  assign n43808 = n39734 & n42591;
  assign n42593 = ~n43812;
  assign n43768 = ~n43814;
  assign n43806 = ~n43815;
  assign n42548 = ~n43816;
  assign n43809 = ~n43828;
  assign n43817 = n43838 & n43839;
  assign n43761 = n43783 ^ n43784;
  assign n43786 = ~n43783;
  assign n43785 = ~n43795;
  assign n43723 = n43806 & n43807;
  assign n42614 = ~n43808;
  assign n43791 = n43809 & n43810;
  assign n43797 = n43817 ^ n41029;
  assign n43818 = ~n43817;
  assign n43739 = n446 ^ n43761;
  assign n43772 = n43785 & n43786;
  assign n43766 = n43791 ^ n43792;
  assign n43790 = n43723 & n43750;
  assign n43788 = ~n43723;
  assign n39530 = n43796 ^ n43797;
  assign n43793 = ~n43791;
  assign n43811 = n43818 & n43819;
  assign n42456 = n43738 ^ n43739;
  assign n43740 = ~n43739;
  assign n43733 = n43765 ^ n43766;
  assign n43759 = ~n43772;
  assign n43771 = n39530 & n43782;
  assign n43773 = n43788 & n43789;
  assign n43774 = n39530 & n42513;
  assign n43752 = ~n43790;
  assign n43775 = n39530 & n41029;
  assign n43787 = n43793 & n43794;
  assign n39660 = ~n39530;
  assign n43798 = ~n43811;
  assign n43691 = ~n42456;
  assign n43689 = n43740 & n43741;
  assign n43747 = n43733 & n6018;
  assign n43754 = n43759 & n43760;
  assign n43748 = ~n43733;
  assign n43764 = n39660 & n43770;
  assign n42553 = ~n43771;
  assign n43726 = ~n43773;
  assign n43762 = ~n43774;
  assign n42538 = ~n43775;
  assign n43767 = ~n43787;
  assign n43776 = n43798 & n43799;
  assign n43731 = ~n43747;
  assign n43742 = n43748 & n445;
  assign n43732 = ~n43754;
  assign n43683 = n43762 & n43763;
  assign n42574 = ~n43764;
  assign n43749 = n43767 & n43768;
  assign n43755 = n43776 ^ n43777;
  assign n43778 = ~n43776;
  assign n43722 = n43731 & n43732;
  assign n43712 = n43732 ^ n43733;
  assign n43714 = ~n43742;
  assign n43724 = n43749 ^ n43750;
  assign n43745 = n43683 & n43753;
  assign n43746 = n42574 & n42553;
  assign n43744 = ~n43683;
  assign n39464 = n40957 ^ n43755;
  assign n43751 = ~n43749;
  assign n43756 = n43755 & n40957;
  assign n43769 = n43778 & n43779;
  assign n43690 = n445 ^ n43712;
  assign n43713 = ~n43722;
  assign n43694 = n43723 ^ n43724;
  assign n43729 = n39464 & n42503;
  assign n43734 = n43744 & n43709;
  assign n43711 = ~n43745;
  assign n42572 = ~n43746;
  assign n43743 = n43751 & n43752;
  assign n39576 = ~n39464;
  assign n42454 = ~n43756;
  assign n43757 = ~n43769;
  assign n42407 = n43689 ^ n43690;
  assign n43688 = ~n43690;
  assign n43693 = n43713 & n43714;
  assign n43706 = n43694 & n5930;
  assign n43707 = ~n43694;
  assign n42528 = ~n43729;
  assign n43721 = n39576 & n43730;
  assign n43686 = ~n43734;
  assign n43727 = n39576 & n42386;
  assign n43725 = ~n43743;
  assign n43735 = n43757 & n43758;
  assign n43658 = n43688 & n43689;
  assign n43675 = n43693 ^ n43694;
  assign n43696 = ~n43693;
  assign n43695 = ~n43706;
  assign n43704 = n43707 & n444;
  assign n42507 = ~n43721;
  assign n43708 = n43725 & n43726;
  assign n43715 = ~n43727;
  assign n43718 = n43735 ^ n40961;
  assign n43736 = ~n43735;
  assign n43659 = n444 ^ n43675;
  assign n43661 = ~n43658;
  assign n43682 = n43695 & n43696;
  assign n43677 = ~n43704;
  assign n43684 = n43708 ^ n43709;
  assign n43654 = n43715 & n43716;
  assign n39399 = n43717 ^ n43718;
  assign n43710 = ~n43708;
  assign n43728 = n43736 & n43737;
  assign n43645 = n43658 ^ n43659;
  assign n43660 = ~n43659;
  assign n43676 = ~n43682;
  assign n43663 = n43683 ^ n43684;
  assign n43692 = n39399 & n42456;
  assign n43699 = n39399 & n42333;
  assign n43700 = n43654 & n43672;
  assign n43701 = n39399 & n40884;
  assign n43705 = n43710 & n43711;
  assign n43697 = ~n43654;
  assign n39417 = ~n39399;
  assign n43719 = ~n43728;
  assign n40478 = n43645 ^ n41413;
  assign n43646 = ~n43645;
  assign n43626 = n43660 & n43661;
  assign n43662 = n43676 & n43677;
  assign n43670 = n43663 & n443;
  assign n43669 = ~n43663;
  assign n43681 = n39417 & n43691;
  assign n42458 = ~n43692;
  assign n43687 = n43697 & n43698;
  assign n43679 = ~n43699;
  assign n43674 = ~n43700;
  assign n42414 = ~n43701;
  assign n43685 = ~n43705;
  assign n43702 = n43719 & n43720;
  assign n43625 = n40478 & n42460;
  assign n42529 = ~n40478;
  assign n43581 = n43646 & n41415;
  assign n43636 = n43646 & n41413;
  assign n43629 = ~n43626;
  assign n43647 = n43662 ^ n43663;
  assign n43653 = ~n43662;
  assign n43666 = n43669 & n5860;
  assign n43638 = ~n43670;
  assign n43622 = n43679 & n43680;
  assign n42482 = ~n43681;
  assign n43671 = n43685 & n43686;
  assign n43657 = ~n43687;
  assign n43678 = n43702 ^ n43703;
  assign n43614 = ~n43625;
  assign n42484 = ~n43636;
  assign n43627 = n443 ^ n43647;
  assign n43652 = ~n43666;
  assign n43655 = n43671 ^ n43672;
  assign n43631 = ~n43622;
  assign n39470 = n43668 ^ n43678;
  assign n43673 = ~n43671;
  assign n43599 = n43614 & n43615;
  assign n43616 = n43626 ^ n43627;
  assign n43628 = ~n43627;
  assign n43649 = n43652 & n43653;
  assign n43619 = n43654 ^ n43655;
  assign n43664 = n39470 & n42337;
  assign n43665 = n39470 & n43668;
  assign n43667 = n43673 & n43674;
  assign n41008 = ~n39470;
  assign n43586 = n43599 ^ n43600;
  assign n43601 = ~n43599;
  assign n43610 = n43616 & n41299;
  assign n43611 = ~n43616;
  assign n43589 = n43628 & n43629;
  assign n43639 = n43619 & n5793;
  assign n43637 = ~n43649;
  assign n43640 = ~n43619;
  assign n43650 = ~n43664;
  assign n42362 = ~n43665;
  assign n43656 = ~n43667;
  assign n42050 = n71 ^ n43586;
  assign n43467 = n43586 & n71;
  assign n43524 = n43601 & n43602;
  assign n43583 = ~n43610;
  assign n43604 = n43611 & n41313;
  assign n43592 = ~n43589;
  assign n43618 = n43637 & n43638;
  assign n43621 = ~n43639;
  assign n43632 = n43640 & n442;
  assign n43633 = n43650 & n43651;
  assign n43641 = n43656 & n43657;
  assign n43305 = ~n42050;
  assign n43597 = ~n43604;
  assign n43605 = n43618 ^ n43619;
  assign n43620 = ~n43618;
  assign n43607 = ~n43632;
  assign n43585 = n43633 ^ n43634;
  assign n43623 = n43641 ^ n43642;
  assign n43644 = n43641 & n43648;
  assign n43643 = ~n43641;
  assign n43588 = n43597 & n43581;
  assign n43580 = n43597 & n43583;
  assign n43590 = n442 ^ n43605;
  assign n43617 = n43620 & n43621;
  assign n43594 = n43622 ^ n43623;
  assign n43635 = n43643 & n43642;
  assign n43630 = ~n43644;
  assign n40290 = n43580 ^ n43581;
  assign n43582 = ~n43588;
  assign n43556 = n43589 ^ n43590;
  assign n43591 = ~n43590;
  assign n43609 = n43594 & n441;
  assign n43606 = ~n43617;
  assign n43608 = ~n43594;
  assign n43624 = n43630 & n43631;
  assign n43613 = ~n43635;
  assign n43569 = n40290 & n42355;
  assign n43570 = n40290 & n41313;
  assign n40457 = ~n40290;
  assign n43571 = n43582 & n43583;
  assign n43575 = n43556 & n41204;
  assign n43576 = ~n43556;
  assign n43563 = n43591 & n43592;
  assign n43593 = n43606 & n43607;
  assign n43603 = n43608 & n5708;
  assign n43579 = ~n43609;
  assign n43612 = ~n43624;
  assign n43560 = ~n43569;
  assign n42382 = ~n43570;
  assign n43557 = n43571 ^ n41250;
  assign n43573 = ~n43571;
  assign n43572 = ~n43575;
  assign n43574 = n43576 & n41250;
  assign n43566 = ~n43563;
  assign n43577 = n43593 ^ n43594;
  assign n43595 = ~n43593;
  assign n43596 = ~n43603;
  assign n43598 = n43612 & n43613;
  assign n40264 = n43556 ^ n43557;
  assign n43550 = n43560 & n43561;
  assign n43562 = n43572 & n43573;
  assign n43559 = ~n43574;
  assign n43564 = n441 ^ n43577;
  assign n43587 = n43595 & n43596;
  assign n43584 = n440 ^ n43598;
  assign n43542 = n40264 & n42287;
  assign n43543 = n40264 & n41204;
  assign n43548 = n43550 & n43551;
  assign n40258 = ~n40264;
  assign n43546 = ~n43550;
  assign n43558 = ~n43562;
  assign n43530 = n43563 ^ n43564;
  assign n43565 = ~n43564;
  assign n43568 = n43584 ^ n43585;
  assign n43578 = ~n43587;
  assign n43532 = ~n43542;
  assign n42318 = ~n43543;
  assign n43544 = n43546 & n43547;
  assign n43535 = ~n43548;
  assign n43545 = n43558 & n43559;
  assign n43552 = n43530 & n41141;
  assign n43553 = ~n43530;
  assign n43554 = n43565 & n43566;
  assign n43567 = n43578 & n43579;
  assign n43494 = n43532 & n43533;
  assign n43534 = n43535 & n43524;
  assign n43527 = ~n43544;
  assign n43531 = n43545 ^ n41141;
  assign n43538 = ~n43545;
  assign n43529 = ~n43552;
  assign n43549 = n43553 & n41159;
  assign n43555 = n43567 ^ n43568;
  assign n43522 = n43494 & n43510;
  assign n43520 = ~n43494;
  assign n40151 = n43530 ^ n43531;
  assign n43526 = ~n43534;
  assign n43523 = n43527 & n43535;
  assign n43539 = ~n43549;
  assign n43500 = n43554 ^ n43555;
  assign n43519 = n43520 & n43521;
  assign n43512 = ~n43522;
  assign n43513 = n43523 ^ n43524;
  assign n43525 = n43526 & n43527;
  assign n40267 = ~n40151;
  assign n43536 = n43538 & n43539;
  assign n43541 = n43500 & n41041;
  assign n43540 = ~n43500;
  assign n43508 = n43513 & n70;
  assign n43498 = ~n43519;
  assign n43514 = n40267 & n42228;
  assign n43515 = n40267 & n41159;
  assign n43507 = ~n43513;
  assign n43509 = ~n43525;
  assign n43528 = ~n43536;
  assign n43537 = n43540 & n41084;
  assign n43502 = ~n43541;
  assign n43505 = n43507 & n3685;
  assign n43478 = ~n43508;
  assign n43495 = n43509 ^ n43510;
  assign n43506 = n43512 & n43509;
  assign n43503 = ~n43514;
  assign n42267 = ~n43515;
  assign n43516 = n43528 & n43529;
  assign n43518 = ~n43537;
  assign n43451 = n43494 ^ n43495;
  assign n43460 = n43503 & n43504;
  assign n43496 = ~n43505;
  assign n43497 = ~n43506;
  assign n43499 = n43516 ^ n41084;
  assign n43517 = ~n43516;
  assign n43474 = n43451 & n69;
  assign n43473 = ~n43451;
  assign n43492 = n43460 & n43493;
  assign n43490 = n43496 & n43467;
  assign n43491 = n43496 & n43478;
  assign n43480 = n43497 & n43498;
  assign n43489 = ~n43460;
  assign n40065 = n43499 ^ n43500;
  assign n43511 = n43517 & n43518;
  assign n43466 = n43473 & n3604;
  assign n43436 = ~n43474;
  assign n43461 = n43480 ^ n43481;
  assign n43482 = n43489 & n43481;
  assign n43477 = ~n43490;
  assign n43468 = ~n43491;
  assign n43483 = n40065 & n42189;
  assign n43475 = ~n43492;
  assign n43484 = n40065 & n41084;
  assign n43476 = ~n43480;
  assign n40128 = ~n40065;
  assign n43501 = ~n43511;
  assign n43418 = n43460 ^ n43461;
  assign n43457 = ~n43466;
  assign n42012 = n43467 ^ n43468;
  assign n43469 = n43475 & n43476;
  assign n43472 = n43477 & n43478;
  assign n43459 = ~n43482;
  assign n43470 = ~n43483;
  assign n42232 = ~n43484;
  assign n43485 = n43501 & n43502;
  assign n43444 = n43418 & n68;
  assign n43443 = ~n43418;
  assign n43263 = ~n42012;
  assign n43458 = ~n43469;
  assign n43420 = n43470 & n43471;
  assign n43450 = ~n43472;
  assign n40034 = n43485 ^ n43486;
  assign n43487 = ~n43485;
  assign n43434 = n43443 & n3531;
  assign n43403 = ~n43444;
  assign n43429 = n43450 ^ n43451;
  assign n43449 = n43457 & n43450;
  assign n43437 = n43458 & n43459;
  assign n43454 = n43420 & n43438;
  assign n43452 = ~n43420;
  assign n43462 = n40034 & n42142;
  assign n43463 = n40034 & n41011;
  assign n40006 = ~n40034;
  assign n43479 = n43487 & n43488;
  assign n41973 = n69 ^ n43429;
  assign n43419 = ~n43434;
  assign n43421 = n43437 ^ n43438;
  assign n43435 = ~n43449;
  assign n43439 = ~n43437;
  assign n43445 = n43452 & n43453;
  assign n43440 = ~n43454;
  assign n43455 = ~n43462;
  assign n42177 = ~n43463;
  assign n43464 = ~n43479;
  assign n43386 = n43420 ^ n43421;
  assign n43235 = ~n41973;
  assign n43430 = n43435 & n43436;
  assign n43431 = n43439 & n43440;
  assign n43423 = ~n43445;
  assign n43389 = n43455 & n43456;
  assign n43446 = n43464 & n43465;
  assign n43404 = n43386 & n3431;
  assign n43405 = ~n43386;
  assign n43417 = ~n43430;
  assign n43422 = ~n43431;
  assign n43433 = n43389 & n43441;
  assign n43432 = ~n43389;
  assign n43424 = n43446 ^ n40892;
  assign n43447 = ~n43446;
  assign n43387 = ~n43404;
  assign n43398 = n43405 & n67;
  assign n43397 = n43417 ^ n43418;
  assign n43416 = n43419 & n43417;
  assign n43406 = n43422 & n43423;
  assign n39930 = n43424 ^ n43425;
  assign n43426 = n43432 & n43407;
  assign n43409 = ~n43433;
  assign n43442 = n43447 & n43448;
  assign n41914 = n68 ^ n43397;
  assign n43370 = ~n43398;
  assign n43390 = n43406 ^ n43407;
  assign n43402 = ~n43416;
  assign n43408 = ~n43406;
  assign n43411 = n39930 & n40892;
  assign n43412 = n39930 & n42097;
  assign n39955 = ~n39930;
  assign n43392 = ~n43426;
  assign n43427 = ~n43442;
  assign n43352 = n43389 ^ n43390;
  assign n41946 = ~n41914;
  assign n43385 = n43402 & n43403;
  assign n43401 = n43408 & n43409;
  assign n42132 = ~n43411;
  assign n43399 = ~n43412;
  assign n43413 = n43427 & n43428;
  assign n43372 = n43352 & n66;
  assign n43371 = ~n43352;
  assign n43368 = n43385 ^ n43386;
  assign n43388 = ~n43385;
  assign n43355 = n43399 & n43400;
  assign n43391 = ~n43401;
  assign n43394 = n43413 ^ n40831;
  assign n43414 = ~n43413;
  assign n43349 = n67 ^ n43368;
  assign n43366 = n43371 & n3384;
  assign n43332 = ~n43372;
  assign n43384 = n43387 & n43388;
  assign n43373 = n43391 & n43392;
  assign n43359 = ~n43355;
  assign n39836 = n43393 ^ n43394;
  assign n43410 = n43414 & n43415;
  assign n43152 = n43349 ^ n41914;
  assign n43350 = ~n43349;
  assign n43353 = ~n43366;
  assign n43356 = n43373 ^ n43374;
  assign n43376 = n43373 & n43380;
  assign n43369 = ~n43384;
  assign n43375 = ~n43373;
  assign n39892 = ~n39836;
  assign n43395 = ~n43410;
  assign n41890 = ~n43152;
  assign n43313 = n43350 & n41946;
  assign n43316 = n43355 ^ n43356;
  assign n43351 = n43369 & n43370;
  assign n43367 = n43375 & n43374;
  assign n43358 = ~n43376;
  assign n43377 = n39892 & n42062;
  assign n43378 = n39892 & n40831;
  assign n43381 = n43395 & n43396;
  assign n43335 = n43316 & n65;
  assign n43334 = ~n43316;
  assign n43333 = n43351 ^ n43352;
  assign n43357 = n43358 & n43359;
  assign n43354 = ~n43351;
  assign n43341 = ~n43367;
  assign n43360 = ~n43377;
  assign n42088 = ~n43378;
  assign n43363 = n43381 ^ n40780;
  assign n43382 = ~n43381;
  assign n43314 = n66 ^ n43333;
  assign n43330 = n43334 & n3342;
  assign n43293 = ~n43335;
  assign n43348 = n43353 & n43354;
  assign n43340 = ~n43357;
  assign n43299 = n43360 & n43361;
  assign n39766 = n43362 ^ n43363;
  assign n43379 = n43382 & n43383;
  assign n43115 = n43313 ^ n43314;
  assign n43272 = n43314 & n43313;
  assign n43318 = ~n43330;
  assign n43320 = n43340 & n43341;
  assign n43331 = ~n43348;
  assign n43344 = n43299 & n43321;
  assign n43342 = ~n43299;
  assign n39788 = ~n39766;
  assign n43364 = ~n43379;
  assign n41850 = ~n43115;
  assign n43300 = n43320 ^ n43321;
  assign n43315 = n43331 & n43332;
  assign n43322 = ~n43320;
  assign n43336 = n43342 & n43343;
  assign n43323 = ~n43344;
  assign n43337 = n39788 & n42018;
  assign n43338 = n39788 & n40761;
  assign n43345 = n43364 & n43365;
  assign n43269 = n43299 ^ n43300;
  assign n43291 = n43315 ^ n43316;
  assign n43319 = n43322 & n43323;
  assign n43317 = ~n43315;
  assign n43298 = ~n43336;
  assign n43324 = ~n43337;
  assign n42056 = ~n43338;
  assign n43326 = n43345 ^ n40738;
  assign n43346 = ~n43345;
  assign n43278 = n43269 & n3315;
  assign n43273 = n65 ^ n43291;
  assign n43279 = ~n43269;
  assign n43311 = n43317 & n43318;
  assign n43297 = ~n43319;
  assign n43257 = n43324 & n43325;
  assign n39682 = n43326 ^ n43327;
  assign n43339 = n43346 & n43347;
  assign n43067 = n43272 ^ n43273;
  assign n43230 = n43273 & n43272;
  assign n43267 = ~n43278;
  assign n43274 = n43279 & n64;
  assign n43280 = n43297 & n43298;
  assign n43292 = ~n43311;
  assign n43302 = n39682 & n41991;
  assign n43303 = n43257 & n43312;
  assign n43304 = n39682 & n42050;
  assign n43306 = n39682 & n40738;
  assign n43301 = ~n43257;
  assign n39707 = ~n39682;
  assign n43328 = ~n43339;
  assign n41813 = ~n43067;
  assign n43252 = ~n43274;
  assign n43258 = n43280 ^ n43281;
  assign n43288 = n43292 & n43293;
  assign n43282 = ~n43280;
  assign n43294 = n43301 & n43281;
  assign n43289 = ~n43302;
  assign n43283 = ~n43303;
  assign n42053 = ~n43304;
  assign n43295 = n39707 & n43305;
  assign n42011 = ~n43306;
  assign n43307 = n43328 & n43329;
  assign n43233 = n43257 ^ n43258;
  assign n43275 = n43282 & n43283;
  assign n43268 = ~n43288;
  assign n43219 = n43289 & n43290;
  assign n43260 = ~n43294;
  assign n42074 = ~n43295;
  assign n43284 = n43307 ^ n43308;
  assign n43309 = ~n43307;
  assign n43239 = n43233 & n79;
  assign n43238 = ~n43233;
  assign n43256 = n43267 & n43268;
  assign n43250 = n43268 ^ n43269;
  assign n43259 = ~n43275;
  assign n43271 = n43219 & n43276;
  assign n43270 = ~n43219;
  assign n39582 = n40685 ^ n43284;
  assign n43285 = ~n43284;
  assign n43296 = n43309 & n43310;
  assign n43236 = n43238 & n3280;
  assign n43197 = ~n43239;
  assign n43231 = n64 ^ n43250;
  assign n43251 = ~n43256;
  assign n43240 = n43259 & n43260;
  assign n43261 = n43270 & n43241;
  assign n43243 = ~n43271;
  assign n43262 = n39582 & n42012;
  assign n39630 = ~n39582;
  assign n43277 = n43285 & n40672;
  assign n43286 = ~n43296;
  assign n41777 = n43230 ^ n43231;
  assign n43192 = n43231 & n43230;
  assign n43217 = ~n43236;
  assign n43220 = n43240 ^ n43241;
  assign n43232 = n43251 & n43252;
  assign n43242 = ~n43240;
  assign n43222 = ~n43261;
  assign n43253 = n39630 & n41952;
  assign n42032 = ~n43262;
  assign n43254 = n39630 & n43263;
  assign n41971 = ~n43277;
  assign n43264 = n43286 & n43287;
  assign n43042 = ~n41777;
  assign n43179 = n43219 ^ n43220;
  assign n43210 = n43232 ^ n43233;
  assign n43218 = ~n43232;
  assign n43237 = n43242 & n43243;
  assign n43244 = ~n43253;
  assign n42015 = ~n43254;
  assign n43246 = n43264 ^ n40661;
  assign n43265 = ~n43264;
  assign n43193 = n79 ^ n43210;
  assign n43199 = n43179 & n78;
  assign n43198 = ~n43179;
  assign n43211 = n43217 & n43218;
  assign n43221 = ~n43237;
  assign n43182 = n43244 & n43245;
  assign n39516 = n43246 ^ n43247;
  assign n43255 = n43265 & n43266;
  assign n41761 = n43192 ^ n43193;
  assign n43137 = n43193 & n43192;
  assign n43194 = n43198 & n3229;
  assign n43161 = ~n43199;
  assign n43196 = ~n43211;
  assign n43200 = n43221 & n43222;
  assign n43224 = n43182 & n43234;
  assign n43225 = n39516 & n43235;
  assign n43223 = ~n43182;
  assign n39518 = ~n39516;
  assign n43248 = ~n43255;
  assign n42989 = ~n41761;
  assign n43181 = ~n43194;
  assign n43178 = n43196 & n43197;
  assign n43183 = n43200 ^ n43201;
  assign n43202 = ~n43200;
  assign n43212 = n43223 & n43201;
  assign n43213 = n39518 & n40661;
  assign n43214 = n39518 & n41905;
  assign n43203 = ~n43224;
  assign n43215 = n39518 & n41973;
  assign n41995 = ~n43225;
  assign n43226 = n43248 & n43249;
  assign n43162 = n43178 ^ n43179;
  assign n43140 = n43182 ^ n43183;
  assign n43180 = ~n43178;
  assign n43195 = n43202 & n43203;
  assign n43185 = ~n43212;
  assign n41943 = ~n43213;
  assign n43204 = ~n43214;
  assign n41976 = ~n43215;
  assign n43206 = n43226 ^ n43227;
  assign n43228 = ~n43226;
  assign n43138 = n78 ^ n43162;
  assign n43163 = n43140 & n77;
  assign n43159 = ~n43140;
  assign n43174 = n43180 & n43181;
  assign n43184 = ~n43195;
  assign n43143 = n43204 & n43205;
  assign n39433 = n43206 ^ n40607;
  assign n43207 = n43206 & n40607;
  assign n43216 = n43228 & n43229;
  assign n41695 = n43137 ^ n43138;
  assign n43095 = n43138 & n43137;
  assign n43157 = n43159 & n3182;
  assign n43120 = ~n43163;
  assign n43160 = ~n43174;
  assign n43164 = n43184 & n43185;
  assign n43188 = n43143 & n43165;
  assign n43186 = ~n43143;
  assign n39435 = ~n39433;
  assign n41877 = ~n43207;
  assign n43208 = ~n43216;
  assign n42948 = ~n41695;
  assign n43098 = ~n43095;
  assign n43141 = ~n43157;
  assign n43139 = n43160 & n43161;
  assign n43144 = n43164 ^ n43165;
  assign n43166 = ~n43164;
  assign n43175 = n43186 & n43187;
  assign n43176 = n39435 & n41862;
  assign n43167 = ~n43188;
  assign n43189 = n43208 & n43209;
  assign n43118 = n43139 ^ n43140;
  assign n43100 = n43143 ^ n43144;
  assign n43142 = ~n43139;
  assign n43158 = n43166 & n43167;
  assign n43146 = ~n43175;
  assign n43168 = ~n43176;
  assign n43171 = n43189 ^ n40552;
  assign n43190 = ~n43189;
  assign n43096 = n77 ^ n43118;
  assign n43121 = n43100 & n3147;
  assign n43122 = ~n43100;
  assign n43133 = n43141 & n43142;
  assign n43145 = ~n43158;
  assign n43103 = n43168 & n43169;
  assign n39405 = n43170 ^ n43171;
  assign n43177 = n43190 & n43191;
  assign n41657 = n43095 ^ n43096;
  assign n43097 = ~n43096;
  assign n43102 = ~n43121;
  assign n43116 = n43122 & n76;
  assign n43119 = ~n43133;
  assign n43123 = n43145 & n43146;
  assign n43148 = n39405 & n40573;
  assign n43149 = n39405 & n41829;
  assign n43150 = n43103 & n43156;
  assign n43151 = n39405 & n41890;
  assign n43147 = ~n43103;
  assign n39356 = ~n39405;
  assign n43172 = ~n43177;
  assign n42903 = ~n41657;
  assign n43052 = n43097 & n43098;
  assign n43077 = ~n43116;
  assign n43099 = n43119 & n43120;
  assign n43104 = n43123 ^ n43124;
  assign n43125 = ~n43123;
  assign n43134 = n43147 & n43124;
  assign n41849 = ~n43148;
  assign n43131 = ~n43149;
  assign n43126 = ~n43150;
  assign n41893 = ~n43151;
  assign n43135 = n39356 & n43152;
  assign n43153 = n43172 & n43173;
  assign n43075 = n43099 ^ n43100;
  assign n43055 = n43103 ^ n43104;
  assign n43101 = ~n43099;
  assign n43117 = n43125 & n43126;
  assign n43058 = n43131 & n43132;
  assign n43106 = ~n43134;
  assign n41910 = ~n43135;
  assign n43128 = n43153 ^ n40523;
  assign n43154 = ~n43153;
  assign n43053 = n76 ^ n43075;
  assign n43079 = n43055 & n75;
  assign n43078 = ~n43055;
  assign n43090 = n43101 & n43102;
  assign n43114 = n43058 & n43081;
  assign n43105 = ~n43117;
  assign n43112 = ~n43058;
  assign n39299 = n43127 ^ n43128;
  assign n43136 = n43154 & n43155;
  assign n41616 = n43052 ^ n43053;
  assign n43009 = n43053 & n43052;
  assign n43073 = n43078 & n3117;
  assign n43034 = ~n43079;
  assign n43076 = ~n43090;
  assign n43080 = n43105 & n43106;
  assign n43107 = n43112 & n43113;
  assign n43083 = ~n43114;
  assign n43108 = n39299 & n43115;
  assign n39343 = ~n39299;
  assign n43129 = ~n43136;
  assign n42859 = ~n41616;
  assign n43057 = ~n43073;
  assign n43054 = n43076 & n43077;
  assign n43059 = n43080 ^ n43081;
  assign n43082 = ~n43080;
  assign n43061 = ~n43107;
  assign n43091 = n39343 & n40520;
  assign n43092 = n39343 & n41772;
  assign n43093 = n39343 & n41850;
  assign n41874 = ~n43108;
  assign n43109 = n43129 & n43130;
  assign n43032 = n43054 ^ n43055;
  assign n43013 = n43058 ^ n43059;
  assign n43056 = ~n43054;
  assign n43074 = n43082 & n43083;
  assign n41818 = ~n43091;
  assign n43084 = ~n43092;
  assign n41855 = ~n43093;
  assign n43087 = n43109 ^ n40467;
  assign n43110 = ~n43109;
  assign n43010 = n75 ^ n43032;
  assign n43035 = n43013 & n3056;
  assign n43036 = ~n43013;
  assign n43048 = n43056 & n43057;
  assign n43060 = ~n43074;
  assign n43014 = n43084 & n43085;
  assign n39336 = n43086 ^ n43087;
  assign n43094 = n43110 & n43111;
  assign n41572 = n43009 ^ n43010;
  assign n43011 = ~n43010;
  assign n43008 = ~n43035;
  assign n43028 = n43036 & n74;
  assign n43033 = ~n43048;
  assign n43037 = n43060 & n43061;
  assign n43063 = n39336 & n40467;
  assign n43064 = n39336 & n41756;
  assign n43065 = n43014 & n43072;
  assign n43066 = n39336 & n41813;
  assign n43062 = ~n43014;
  assign n39260 = ~n39336;
  assign n43088 = ~n43094;
  assign n42820 = ~n41572;
  assign n42974 = n43011 & n43009;
  assign n42994 = ~n43028;
  assign n43012 = n43033 & n43034;
  assign n43015 = n43037 ^ n43038;
  assign n43039 = ~n43037;
  assign n43049 = n43062 & n43038;
  assign n41774 = ~n43063;
  assign n43046 = ~n43064;
  assign n43040 = ~n43065;
  assign n41816 = ~n43066;
  assign n43050 = n39260 & n43067;
  assign n43069 = n43088 & n43089;
  assign n42977 = ~n42974;
  assign n42992 = n43012 ^ n43013;
  assign n42979 = n43014 ^ n43015;
  assign n43007 = ~n43012;
  assign n43029 = n43039 & n43040;
  assign n42972 = n43046 & n43047;
  assign n43017 = ~n43049;
  assign n41837 = ~n43050;
  assign n39197 = n43068 ^ n43069;
  assign n43070 = ~n43069;
  assign n42975 = n74 ^ n42992;
  assign n42996 = n42979 & n73;
  assign n42995 = ~n42979;
  assign n43005 = n43007 & n43008;
  assign n43016 = ~n43029;
  assign n43025 = n42972 & n42998;
  assign n43023 = ~n42972;
  assign n43041 = n39197 & n41713;
  assign n43043 = n39197 & n41777;
  assign n39241 = ~n39197;
  assign n43051 = n43070 & n43071;
  assign n41534 = n42974 ^ n42975;
  assign n42976 = ~n42975;
  assign n42990 = n42995 & n3021;
  assign n42955 = ~n42996;
  assign n42993 = ~n43005;
  assign n42997 = n43016 & n43017;
  assign n43018 = n43023 & n43024;
  assign n43000 = ~n43025;
  assign n43030 = n39241 & n40399;
  assign n43026 = ~n43041;
  assign n43031 = n39241 & n43042;
  assign n41796 = ~n43043;
  assign n43044 = ~n43051;
  assign n42791 = ~n41534;
  assign n42932 = n42976 & n42977;
  assign n42981 = ~n42990;
  assign n42978 = n42993 & n42994;
  assign n42973 = n42997 ^ n42998;
  assign n42999 = ~n42997;
  assign n42983 = ~n43018;
  assign n42918 = n43026 & n43027;
  assign n41734 = ~n43030;
  assign n41780 = ~n43031;
  assign n43019 = n43044 & n43045;
  assign n42931 = ~n42932;
  assign n42935 = n42972 ^ n42973;
  assign n42953 = n42978 ^ n42979;
  assign n42980 = ~n42978;
  assign n42991 = n42999 & n43000;
  assign n43001 = n43019 ^ n43020;
  assign n43021 = ~n43019;
  assign n42933 = n73 ^ n42953;
  assign n42956 = n42935 & n2975;
  assign n42957 = ~n42935;
  assign n42969 = n42980 & n42981;
  assign n42982 = ~n42991;
  assign n39227 = n43001 ^ n40410;
  assign n43002 = n43001 & n40376;
  assign n43006 = n43021 & n43022;
  assign n41492 = n42932 ^ n42933;
  assign n42930 = ~n42933;
  assign n42937 = ~n42956;
  assign n42950 = n42957 & n72;
  assign n42954 = ~n42969;
  assign n42965 = n42982 & n42983;
  assign n42984 = n39227 & n41654;
  assign n42985 = n39227 & n42989;
  assign n39159 = ~n39227;
  assign n41703 = ~n43002;
  assign n43003 = ~n43006;
  assign n42749 = ~n41492;
  assign n42891 = n42930 & n42931;
  assign n42916 = ~n42950;
  assign n42934 = n42954 & n42955;
  assign n42960 = n42965 & n42966;
  assign n42958 = ~n42965;
  assign n42970 = n39159 & n41761;
  assign n42967 = ~n42984;
  assign n41740 = ~n42985;
  assign n42986 = n43003 & n43004;
  assign n42894 = ~n42891;
  assign n42914 = n42934 ^ n42935;
  assign n42936 = ~n42934;
  assign n42951 = n42958 & n42959;
  assign n42939 = ~n42960;
  assign n42908 = n42967 & n42968;
  assign n41763 = ~n42970;
  assign n42961 = n42986 ^ n40345;
  assign n42987 = ~n42986;
  assign n42892 = n72 ^ n42914;
  assign n42927 = n42936 & n42937;
  assign n42938 = n42939 & n42918;
  assign n42924 = ~n42951;
  assign n42949 = n42908 & n42952;
  assign n42947 = ~n42908;
  assign n39192 = n42961 ^ n42962;
  assign n42971 = n42987 & n42988;
  assign n42696 = n42891 ^ n42892;
  assign n42893 = ~n42892;
  assign n42915 = ~n42927;
  assign n42923 = ~n42938;
  assign n42917 = n42924 & n42939;
  assign n42940 = n42947 & n42883;
  assign n42941 = n39192 & n40345;
  assign n42942 = n39192 & n42948;
  assign n42943 = n39192 & n41643;
  assign n42910 = ~n42949;
  assign n39125 = ~n39192;
  assign n42963 = ~n42971;
  assign n41449 = ~n42696;
  assign n42850 = n42893 & n42894;
  assign n42895 = n42915 & n42916;
  assign n42875 = n42917 ^ n42918;
  assign n42907 = n42923 & n42924;
  assign n42885 = ~n42940;
  assign n41665 = ~n42941;
  assign n41698 = ~n42942;
  assign n42925 = ~n42943;
  assign n42928 = n39125 & n41695;
  assign n42944 = n42963 & n42964;
  assign n42874 = n87 ^ n42895;
  assign n42897 = n42875 & n87;
  assign n42882 = n42907 ^ n42908;
  assign n42877 = ~n42895;
  assign n42896 = ~n42875;
  assign n42909 = ~n42907;
  assign n42842 = n42925 & n42926;
  assign n41719 = ~n42928;
  assign n42920 = n42944 ^ n40250;
  assign n42945 = ~n42944;
  assign n42851 = n42874 ^ n42875;
  assign n42837 = n42882 ^ n42883;
  assign n42888 = n42896 & n2910;
  assign n42854 = ~n42897;
  assign n42898 = n42909 & n42910;
  assign n42912 = n42842 & n42913;
  assign n42911 = ~n42842;
  assign n39105 = n42919 ^ n42920;
  assign n42929 = n42945 & n42946;
  assign n41423 = n42850 ^ n42851;
  assign n42793 = n42851 & n42850;
  assign n42865 = n42837 & n86;
  assign n42864 = ~n42837;
  assign n42876 = ~n42888;
  assign n42884 = ~n42898;
  assign n42899 = n42911 & n42867;
  assign n42900 = n39105 & n40250;
  assign n42901 = n39105 & n41657;
  assign n42869 = ~n42912;
  assign n42902 = n39105 & n41563;
  assign n39117 = ~n39105;
  assign n42921 = ~n42929;
  assign n42665 = ~n41423;
  assign n42852 = n42864 & n2896;
  assign n42815 = ~n42865;
  assign n42872 = n42876 & n42877;
  assign n42866 = n42884 & n42885;
  assign n42845 = ~n42899;
  assign n41615 = ~n42900;
  assign n41660 = ~n42901;
  assign n42886 = ~n42902;
  assign n42889 = n39117 & n42903;
  assign n42904 = n42921 & n42922;
  assign n42834 = ~n42852;
  assign n42843 = n42866 ^ n42867;
  assign n42853 = ~n42872;
  assign n42868 = ~n42866;
  assign n42805 = n42886 & n42887;
  assign n41682 = ~n42889;
  assign n42878 = n42904 ^ n40261;
  assign n42905 = ~n42904;
  assign n42796 = n42842 ^ n42843;
  assign n42836 = n42853 & n42854;
  assign n42855 = n42868 & n42869;
  assign n42871 = n42805 & n42873;
  assign n42870 = ~n42805;
  assign n39128 = n42878 ^ n42879;
  assign n42890 = n42905 & n42906;
  assign n42825 = n42796 & n85;
  assign n42813 = n42836 ^ n42837;
  assign n42824 = ~n42796;
  assign n42835 = ~n42836;
  assign n42844 = ~n42855;
  assign n42856 = n42870 & n42827;
  assign n42857 = n39128 & n41616;
  assign n42858 = n39128 & n41524;
  assign n42829 = ~n42871;
  assign n42860 = n39128 & n40261;
  assign n39062 = ~n39128;
  assign n42880 = ~n42890;
  assign n42794 = n86 ^ n42813;
  assign n42816 = n42824 & n2826;
  assign n42773 = ~n42825;
  assign n42833 = n42834 & n42835;
  assign n42826 = n42844 & n42845;
  assign n42808 = ~n42856;
  assign n41619 = ~n42857;
  assign n42846 = ~n42858;
  assign n42848 = n39062 & n42859;
  assign n41571 = ~n42860;
  assign n42861 = n42880 & n42881;
  assign n42610 = n42793 ^ n42794;
  assign n42752 = n42794 & n42793;
  assign n42797 = ~n42816;
  assign n42806 = n42826 ^ n42827;
  assign n42814 = ~n42833;
  assign n42828 = ~n42826;
  assign n42762 = n42846 & n42847;
  assign n41639 = ~n42848;
  assign n42839 = n42861 ^ n40109;
  assign n42862 = ~n42861;
  assign n41339 = ~n42610;
  assign n42755 = n42805 ^ n42806;
  assign n42795 = n42814 & n42815;
  assign n42817 = n42828 & n42829;
  assign n42831 = n42762 & n42832;
  assign n42830 = ~n42762;
  assign n39028 = n42838 ^ n42839;
  assign n42849 = n42862 & n42863;
  assign n42786 = n42755 & n84;
  assign n42771 = n42795 ^ n42796;
  assign n42785 = ~n42755;
  assign n42798 = ~n42795;
  assign n42807 = ~n42817;
  assign n42818 = n42830 & n42788;
  assign n42819 = n39028 & n41572;
  assign n42790 = ~n42831;
  assign n39032 = ~n39028;
  assign n42840 = ~n42849;
  assign n42753 = n85 ^ n42771;
  assign n42774 = n42785 & n2783;
  assign n42732 = ~n42786;
  assign n42792 = n42797 & n42798;
  assign n42787 = n42807 & n42808;
  assign n42765 = ~n42818;
  assign n42809 = n39032 & n40109;
  assign n42810 = n39032 & n41515;
  assign n41600 = ~n42819;
  assign n42811 = n39032 & n42820;
  assign n42821 = n42840 & n42841;
  assign n41274 = n42752 ^ n42753;
  assign n42710 = n42753 & n42752;
  assign n42757 = ~n42774;
  assign n42763 = n42787 ^ n42788;
  assign n42772 = ~n42792;
  assign n42789 = ~n42787;
  assign n41532 = ~n42809;
  assign n42799 = ~n42810;
  assign n41575 = ~n42811;
  assign n42802 = n42821 ^ n40044;
  assign n42822 = ~n42821;
  assign n42570 = ~n41274;
  assign n42713 = n42762 ^ n42763;
  assign n42754 = n42772 & n42773;
  assign n42775 = n42789 & n42790;
  assign n42722 = n42799 & n42800;
  assign n38964 = n42801 ^ n42802;
  assign n42812 = n42822 & n42823;
  assign n42742 = n42713 & n83;
  assign n42730 = n42754 ^ n42755;
  assign n42741 = ~n42713;
  assign n42756 = ~n42754;
  assign n42764 = ~n42775;
  assign n42778 = n38964 & n40122;
  assign n42779 = n38964 & n41433;
  assign n42780 = n42722 & n42744;
  assign n42781 = n38964 & n42791;
  assign n42776 = ~n42722;
  assign n38996 = ~n38964;
  assign n42803 = ~n42812;
  assign n42711 = n84 ^ n42730;
  assign n42733 = n42741 & n2766;
  assign n42691 = ~n42742;
  assign n42751 = n42756 & n42757;
  assign n42743 = n42764 & n42765;
  assign n42768 = n42776 & n42777;
  assign n41491 = ~n42778;
  assign n42766 = ~n42779;
  assign n42746 = ~n42780;
  assign n42769 = n38996 & n41534;
  assign n41536 = ~n42781;
  assign n42782 = n42803 & n42804;
  assign n41210 = n42710 ^ n42711;
  assign n42668 = n42711 & n42710;
  assign n42714 = ~n42733;
  assign n42723 = n42743 ^ n42744;
  assign n42731 = ~n42751;
  assign n42745 = ~n42743;
  assign n42680 = n42766 & n42767;
  assign n42725 = ~n42768;
  assign n41559 = ~n42769;
  assign n42759 = n42782 ^ n39963;
  assign n42783 = ~n42782;
  assign n42558 = ~n41210;
  assign n42671 = ~n42668;
  assign n42673 = n42722 ^ n42723;
  assign n42712 = n42731 & n42732;
  assign n42734 = n42745 & n42746;
  assign n42750 = n42680 & n42706;
  assign n42747 = ~n42680;
  assign n38937 = n42758 ^ n42759;
  assign n42770 = n42783 & n42784;
  assign n42703 = n42673 & n2673;
  assign n42689 = n42712 ^ n42713;
  assign n42704 = ~n42673;
  assign n42715 = ~n42712;
  assign n42724 = ~n42734;
  assign n42735 = n42747 & n42748;
  assign n42736 = n38937 & n42749;
  assign n42708 = ~n42750;
  assign n38975 = ~n38937;
  assign n42760 = ~n42770;
  assign n42669 = n83 ^ n42689;
  assign n42675 = ~n42703;
  assign n42692 = n42704 & n82;
  assign n42709 = n42714 & n42715;
  assign n42705 = n42724 & n42725;
  assign n42683 = ~n42735;
  assign n42726 = n38975 & n39963;
  assign n41520 = ~n42736;
  assign n42727 = n38975 & n41492;
  assign n42728 = n38975 & n41437;
  assign n42737 = n42760 & n42761;
  assign n41132 = n42668 ^ n42669;
  assign n42670 = ~n42669;
  assign n42647 = ~n42692;
  assign n42681 = n42705 ^ n42706;
  assign n42690 = ~n42709;
  assign n42707 = ~n42705;
  assign n41459 = ~n42726;
  assign n41495 = ~n42727;
  assign n42716 = ~n42728;
  assign n42718 = n42737 ^ n42738;
  assign n42739 = ~n42737;
  assign n42492 = ~n41132;
  assign n42625 = n42670 & n42671;
  assign n42630 = n42680 ^ n42681;
  assign n42672 = n42690 & n42691;
  assign n42693 = n42707 & n42708;
  assign n42637 = n42716 & n42717;
  assign n38884 = n39965 ^ n42718;
  assign n42719 = n42718 & n39821;
  assign n42729 = n42739 & n42740;
  assign n42628 = ~n42625;
  assign n42657 = n42630 & n2621;
  assign n42645 = n42672 ^ n42673;
  assign n42658 = ~n42630;
  assign n42674 = ~n42672;
  assign n42682 = ~n42693;
  assign n42697 = n38884 & n41379;
  assign n42698 = n42637 & n42660;
  assign n42699 = n38884 & n41449;
  assign n42694 = ~n42637;
  assign n38955 = ~n38884;
  assign n41405 = ~n42719;
  assign n42720 = ~n42729;
  assign n42626 = n82 ^ n42645;
  assign n42632 = ~n42657;
  assign n42648 = n42658 & n81;
  assign n42666 = n42674 & n42675;
  assign n42659 = n42682 & n42683;
  assign n42686 = n42694 & n42695;
  assign n42687 = n38955 & n42696;
  assign n42684 = ~n42697;
  assign n42662 = ~n42698;
  assign n41451 = ~n42699;
  assign n42700 = n42720 & n42721;
  assign n41051 = n42625 ^ n42626;
  assign n42627 = ~n42626;
  assign n42603 = ~n42648;
  assign n42638 = n42659 ^ n42660;
  assign n42646 = ~n42666;
  assign n42661 = ~n42659;
  assign n42618 = n42684 & n42685;
  assign n42640 = ~n42686;
  assign n41477 = ~n42687;
  assign n42676 = n42700 ^ n39791;
  assign n42701 = ~n42700;
  assign n42442 = ~n41051;
  assign n42352 = n42627 & n42628;
  assign n42587 = n42637 ^ n42638;
  assign n42629 = n42646 & n42647;
  assign n42649 = n42661 & n42662;
  assign n42664 = n42618 & n42667;
  assign n42663 = ~n42618;
  assign n38853 = n42676 ^ n42677;
  assign n42688 = n42701 & n42702;
  assign n42615 = n42587 & n2593;
  assign n42604 = n42629 ^ n42630;
  assign n42616 = ~n42587;
  assign n42631 = ~n42629;
  assign n42639 = ~n42649;
  assign n42650 = n42663 & n42595;
  assign n42651 = n38853 & n39791;
  assign n42652 = n38853 & n41327;
  assign n42620 = ~n42664;
  assign n42653 = n38853 & n42665;
  assign n38940 = ~n38853;
  assign n42678 = ~n42688;
  assign n42377 = n81 ^ n42604;
  assign n42589 = ~n42615;
  assign n42605 = n42616 & n80;
  assign n42624 = n42631 & n42632;
  assign n42617 = n42639 & n42640;
  assign n42597 = ~n42650;
  assign n41353 = ~n42651;
  assign n42643 = n38940 & n41423;
  assign n42641 = ~n42652;
  assign n41393 = ~n42653;
  assign n42654 = n42678 & n42679;
  assign n42585 = ~n42377;
  assign n42565 = ~n42605;
  assign n42594 = n42617 ^ n42618;
  assign n42602 = ~n42624;
  assign n42619 = ~n42617;
  assign n42578 = n42641 & n42642;
  assign n41425 = ~n42643;
  assign n42633 = n42654 ^ n39824;
  assign n42655 = ~n42654;
  assign n42541 = n42585 & n42352;
  assign n42519 = n42594 ^ n42595;
  assign n42586 = n42602 & n42603;
  assign n42606 = n42619 & n42620;
  assign n42623 = n42578 & n42555;
  assign n42621 = ~n42578;
  assign n38816 = n42633 ^ n42634;
  assign n42644 = n42655 & n42656;
  assign n42576 = n42519 & n95;
  assign n42563 = n42586 ^ n42587;
  assign n42575 = ~n42519;
  assign n42588 = ~n42586;
  assign n42596 = ~n42606;
  assign n42607 = n42621 & n42622;
  assign n42608 = n38816 & n39824;
  assign n42609 = n38816 & n41339;
  assign n42611 = n38816 & n41195;
  assign n42580 = ~n42623;
  assign n38906 = ~n38816;
  assign n42635 = ~n42644;
  assign n42542 = n80 ^ n42563;
  assign n42566 = n42575 & n2483;
  assign n42521 = ~n42576;
  assign n42584 = n42588 & n42589;
  assign n42577 = n42596 & n42597;
  assign n42557 = ~n42607;
  assign n41292 = ~n42608;
  assign n41341 = ~n42609;
  assign n42600 = n38906 & n42610;
  assign n42598 = ~n42611;
  assign n42612 = n42635 & n42636;
  assign n40496 = n42541 ^ n42542;
  assign n42543 = ~n42542;
  assign n42546 = ~n42566;
  assign n42554 = n42577 ^ n42578;
  assign n42564 = ~n42584;
  assign n42579 = ~n42577;
  assign n42533 = n42598 & n42599;
  assign n41368 = ~n42600;
  assign n42590 = n42612 ^ n39734;
  assign n42613 = ~n42612;
  assign n38663 = n40496 ^ n40478;
  assign n42517 = n40496 & n42529;
  assign n42421 = n40496 & n40478;
  assign n42495 = n42543 & n42541;
  assign n42500 = n42554 ^ n42555;
  assign n42544 = n42564 & n42565;
  assign n42567 = n42579 & n42580;
  assign n42583 = n42533 & n42509;
  assign n42581 = ~n42533;
  assign n38800 = n42590 ^ n42591;
  assign n42601 = n42613 & n42614;
  assign n42494 = n38663 & n41415;
  assign n41445 = ~n42517;
  assign n42498 = ~n42495;
  assign n42530 = n42500 & n2398;
  assign n42518 = n95 ^ n42544;
  assign n42531 = ~n42500;
  assign n42545 = ~n42544;
  assign n42556 = ~n42567;
  assign n42568 = n42581 & n42582;
  assign n42569 = n38800 & n41274;
  assign n42535 = ~n42583;
  assign n38837 = ~n38800;
  assign n42592 = ~n42601;
  assign n42483 = ~n42494;
  assign n42496 = n42518 ^ n42519;
  assign n42502 = ~n42530;
  assign n42522 = n42531 & n94;
  assign n42539 = n42545 & n42546;
  assign n42532 = n42556 & n42557;
  assign n42511 = ~n42568;
  assign n41311 = ~n42569;
  assign n42559 = n38837 & n39734;
  assign n42560 = n38837 & n42570;
  assign n42561 = n38837 & n41110;
  assign n42571 = n42592 & n42593;
  assign n42461 = n42483 & n42484;
  assign n42485 = n42495 ^ n42496;
  assign n42497 = ~n42496;
  assign n42476 = ~n42522;
  assign n42508 = n42532 ^ n42533;
  assign n42520 = ~n42539;
  assign n42534 = ~n42532;
  assign n41209 = ~n42559;
  assign n41277 = ~n42560;
  assign n42547 = ~n42561;
  assign n38792 = n42571 ^ n42572;
  assign n42573 = ~n42571;
  assign n42435 = n42461 ^ n42462;
  assign n42459 = ~n42461;
  assign n42472 = n42485 & n40290;
  assign n42473 = ~n42485;
  assign n42447 = n42497 & n42498;
  assign n42450 = n42508 ^ n42509;
  assign n42499 = n42520 & n42521;
  assign n42523 = n42534 & n42535;
  assign n42463 = n42547 & n42548;
  assign n42549 = n38792 & n42558;
  assign n42550 = n38792 & n39660;
  assign n42551 = n38792 & n41114;
  assign n38763 = ~n38792;
  assign n42562 = n42573 & n42574;
  assign n40571 = n231 ^ n42435;
  assign n42230 = n42435 & n231;
  assign n42307 = n42459 & n42460;
  assign n42423 = ~n42472;
  assign n42467 = n42473 & n40457;
  assign n42486 = n42450 & n2323;
  assign n42474 = n42499 ^ n42500;
  assign n42487 = ~n42450;
  assign n42501 = ~n42499;
  assign n42510 = ~n42523;
  assign n42525 = n42463 & n42536;
  assign n42524 = ~n42463;
  assign n41213 = ~n42549;
  assign n41155 = ~n42550;
  assign n42540 = n38763 & n41210;
  assign n42537 = ~n42551;
  assign n42552 = ~n42562;
  assign n40595 = ~n40571;
  assign n42446 = ~n42467;
  assign n42448 = n94 ^ n42474;
  assign n42452 = ~n42486;
  assign n42477 = n42487 & n93;
  assign n42493 = n42501 & n42502;
  assign n42488 = n42510 & n42511;
  assign n42515 = n42524 & n42489;
  assign n42491 = ~n42525;
  assign n42409 = n42537 & n42538;
  assign n41246 = ~n42540;
  assign n42526 = n42552 & n42553;
  assign n42444 = n42446 & n42421;
  assign n42420 = n42446 & n42423;
  assign n42366 = n42447 ^ n42448;
  assign n42399 = n42448 & n42447;
  assign n42419 = ~n42477;
  assign n42464 = n42488 ^ n42489;
  assign n42475 = ~n42493;
  assign n42490 = ~n42488;
  assign n42466 = ~n42515;
  assign n42514 = n42409 & n42439;
  assign n42512 = ~n42409;
  assign n42504 = n42526 ^ n39464;
  assign n42527 = ~n42526;
  assign n38626 = n42420 ^ n42421;
  assign n42424 = n42366 & n40264;
  assign n42422 = ~n42444;
  assign n42425 = ~n42366;
  assign n42402 = ~n42399;
  assign n42404 = n42463 ^ n42464;
  assign n42449 = n42475 & n42476;
  assign n42478 = n42490 & n42491;
  assign n38731 = n42503 ^ n42504;
  assign n42505 = n42512 & n42513;
  assign n42441 = ~n42514;
  assign n42516 = n42527 & n42528;
  assign n42396 = n38626 & n40457;
  assign n42397 = n38626 & n41299;
  assign n38621 = ~n38626;
  assign n42398 = n42422 & n42423;
  assign n42369 = ~n42424;
  assign n42415 = n42425 & n40258;
  assign n42437 = n42404 & n92;
  assign n42426 = n42449 ^ n42450;
  assign n42436 = ~n42404;
  assign n42451 = ~n42449;
  assign n42465 = ~n42478;
  assign n42479 = n38731 & n42492;
  assign n38757 = ~n38731;
  assign n42412 = ~n42505;
  assign n42506 = ~n42516;
  assign n41333 = ~n42396;
  assign n42381 = ~n42397;
  assign n42367 = n42398 ^ n40264;
  assign n42395 = ~n42398;
  assign n42394 = ~n42415;
  assign n42400 = n93 ^ n42426;
  assign n42427 = n42436 & n2217;
  assign n42374 = ~n42437;
  assign n42445 = n42451 & n42452;
  assign n42438 = n42465 & n42466;
  assign n41177 = ~n42479;
  assign n42468 = n38757 & n39464;
  assign n42469 = n38757 & n41132;
  assign n42470 = n38757 & n41033;
  assign n42480 = n42506 & n42507;
  assign n38611 = n42366 ^ n42367;
  assign n42363 = n42381 & n42382;
  assign n42391 = n42394 & n42395;
  assign n42315 = n42399 ^ n42400;
  assign n42401 = ~n42400;
  assign n42406 = ~n42427;
  assign n42410 = n42438 ^ n42439;
  assign n42418 = ~n42445;
  assign n42440 = ~n42438;
  assign n41070 = ~n42468;
  assign n41135 = ~n42469;
  assign n42453 = ~n42470;
  assign n42455 = n42480 ^ n39417;
  assign n42481 = ~n42480;
  assign n42356 = n42363 & n42364;
  assign n38589 = ~n38611;
  assign n42354 = ~n42363;
  assign n42370 = n42315 & n40151;
  assign n42368 = ~n42391;
  assign n42371 = ~n42315;
  assign n42346 = n42401 & n42402;
  assign n42349 = n42409 ^ n42410;
  assign n42403 = n42418 & n42419;
  assign n42428 = n42440 & n42441;
  assign n42357 = n42453 & n42454;
  assign n38724 = n42455 ^ n42456;
  assign n42471 = n42481 & n42482;
  assign n42338 = n38589 & n40258;
  assign n42339 = n38589 & n41250;
  assign n42342 = n42354 & n42355;
  assign n42328 = ~n42356;
  assign n42343 = n42368 & n42369;
  assign n42344 = ~n42370;
  assign n42365 = n42371 & n40267;
  assign n42383 = n42349 & n2139;
  assign n42372 = n42403 ^ n42404;
  assign n42384 = ~n42349;
  assign n42405 = ~n42403;
  assign n42411 = ~n42428;
  assign n42430 = n38724 & n39417;
  assign n42431 = n38724 & n42442;
  assign n42432 = n38724 & n40961;
  assign n42433 = n42357 & n42443;
  assign n42429 = ~n42357;
  assign n38701 = ~n38724;
  assign n42457 = ~n42471;
  assign n42327 = n42328 & n42307;
  assign n41279 = ~n42338;
  assign n42317 = ~n42339;
  assign n42313 = ~n42342;
  assign n42316 = n42343 ^ n40151;
  assign n42345 = ~n42343;
  assign n42320 = ~n42365;
  assign n42347 = n92 ^ n42372;
  assign n42351 = ~n42383;
  assign n42375 = n42384 & n91;
  assign n42392 = n42405 & n42406;
  assign n42385 = n42411 & n42412;
  assign n42416 = n42429 & n42386;
  assign n40993 = ~n42430;
  assign n41116 = ~n42431;
  assign n42417 = n38701 & n41051;
  assign n42413 = ~n42432;
  assign n42388 = ~n42433;
  assign n42434 = n42457 & n42458;
  assign n38563 = n42315 ^ n42316;
  assign n42264 = n42317 & n42318;
  assign n42312 = ~n42327;
  assign n42306 = n42313 & n42328;
  assign n42340 = n42344 & n42345;
  assign n42329 = n42346 ^ n42347;
  assign n42298 = n42347 & n42346;
  assign n42324 = ~n42375;
  assign n42358 = n42385 ^ n42386;
  assign n42373 = ~n42392;
  assign n42387 = ~n42385;
  assign n42308 = n42413 & n42414;
  assign n42360 = ~n42416;
  assign n41074 = ~n42417;
  assign n42408 = n42434 ^ n39470;
  assign n42294 = n42264 & n42305;
  assign n42285 = n42306 ^ n42307;
  assign n42293 = ~n42264;
  assign n42286 = n42312 & n42313;
  assign n38585 = ~n38563;
  assign n42321 = n42329 & n40128;
  assign n42319 = ~n42340;
  assign n42271 = ~n42329;
  assign n42302 = n42357 ^ n42358;
  assign n42348 = n42373 & n42374;
  assign n42376 = n42387 & n42388;
  assign n42390 = n42308 & n42393;
  assign n42389 = ~n42308;
  assign n38713 = n42407 ^ n42408;
  assign n42281 = n42285 & n230;
  assign n42265 = n42286 ^ n42287;
  assign n42288 = n42293 & n42287;
  assign n42289 = n38585 & n40151;
  assign n42290 = n38585 & n41141;
  assign n42279 = ~n42294;
  assign n42278 = ~n42285;
  assign n42280 = ~n42286;
  assign n42295 = n42319 & n42320;
  assign n42314 = n42271 & n40065;
  assign n42296 = ~n42321;
  assign n42331 = n42302 & n90;
  assign n42322 = n42348 ^ n42349;
  assign n42330 = ~n42302;
  assign n42350 = ~n42348;
  assign n42359 = ~n42376;
  assign n42353 = n42377 ^ n38713;
  assign n42378 = n42389 & n42333;
  assign n42379 = n38713 & n39470;
  assign n42380 = n38713 & n40933;
  assign n42335 = ~n42390;
  assign n39539 = ~n38713;
  assign n42209 = n42264 ^ n42265;
  assign n42269 = n42278 & n19809;
  assign n42268 = n42279 & n42280;
  assign n42236 = ~n42281;
  assign n42259 = ~n42288;
  assign n41179 = ~n42289;
  assign n42266 = ~n42290;
  assign n42270 = n42295 ^ n40128;
  assign n42297 = ~n42295;
  assign n42273 = ~n42314;
  assign n42299 = n91 ^ n42322;
  assign n42325 = n42330 & n2082;
  assign n42276 = ~n42331;
  assign n42341 = n42350 & n42351;
  assign n41037 = n42352 ^ n42353;
  assign n42332 = n42359 & n42360;
  assign n42311 = ~n42378;
  assign n40972 = ~n42379;
  assign n42361 = ~n42380;
  assign n42240 = n42209 & n229;
  assign n42239 = ~n42209;
  assign n42203 = n42266 & n42267;
  assign n42258 = ~n42268;
  assign n42260 = ~n42269;
  assign n38552 = n42270 ^ n42271;
  assign n42291 = n42296 & n42297;
  assign n42219 = n42298 ^ n42299;
  assign n42300 = ~n42299;
  assign n42303 = ~n42325;
  assign n42309 = n42332 ^ n42333;
  assign n42323 = ~n42341;
  assign n42334 = ~n42332;
  assign n42336 = n42361 & n42362;
  assign n42226 = n42239 & n19742;
  assign n42187 = ~n42240;
  assign n42227 = n42258 & n42259;
  assign n42245 = n42260 & n42230;
  assign n42229 = n42260 & n42236;
  assign n42246 = n38552 & n40128;
  assign n42247 = n42203 & n42261;
  assign n42248 = n38552 & n41041;
  assign n42244 = ~n42203;
  assign n38532 = ~n38552;
  assign n42272 = ~n42291;
  assign n42252 = n42300 & n42298;
  assign n42255 = n42308 ^ n42309;
  assign n42301 = n42323 & n42324;
  assign n42326 = n42334 & n42335;
  assign n42263 = n42336 ^ n42337;
  assign n42206 = ~n42226;
  assign n42204 = n42227 ^ n42228;
  assign n42205 = n42229 ^ n42230;
  assign n42234 = ~n42227;
  assign n42241 = n42244 & n42228;
  assign n42235 = ~n42245;
  assign n41119 = ~n42246;
  assign n42233 = ~n42247;
  assign n42231 = ~n42248;
  assign n42249 = n42272 & n42273;
  assign n42283 = n42255 & n89;
  assign n42274 = n42301 ^ n42302;
  assign n42282 = ~n42255;
  assign n42304 = ~n42301;
  assign n42310 = ~n42326;
  assign n42154 = n42203 ^ n42204;
  assign n40542 = n42205 ^ n40571;
  assign n42161 = n42205 & n40571;
  assign n42159 = n42231 & n42232;
  assign n42218 = n42233 & n42234;
  assign n42208 = n42235 & n42236;
  assign n42211 = ~n42241;
  assign n42220 = n42249 ^ n40034;
  assign n42251 = n42249 & n40006;
  assign n42250 = ~n42249;
  assign n42253 = n90 ^ n42274;
  assign n42277 = n42282 & n2029;
  assign n42225 = ~n42283;
  assign n42292 = n42303 & n42304;
  assign n42284 = n42310 & n42311;
  assign n42185 = n42154 & n228;
  assign n41799 = ~n40542;
  assign n42184 = ~n42154;
  assign n42183 = n42208 ^ n42209;
  assign n42213 = n42159 & n42216;
  assign n42212 = ~n42159;
  assign n42210 = ~n42218;
  assign n42207 = ~n42208;
  assign n38493 = n42219 ^ n42220;
  assign n42242 = n42250 & n40034;
  assign n42237 = ~n42251;
  assign n42238 = n42252 ^ n42253;
  assign n42199 = n42253 & n42252;
  assign n42257 = ~n42277;
  assign n42262 = n88 ^ n42284;
  assign n42275 = ~n42292;
  assign n42162 = n229 ^ n42183;
  assign n42173 = n42184 & n19716;
  assign n42138 = ~n42185;
  assign n42197 = n42206 & n42207;
  assign n42188 = n42210 & n42211;
  assign n42198 = n42212 & n42189;
  assign n42190 = ~n42213;
  assign n38500 = ~n38493;
  assign n42221 = n42237 & n42219;
  assign n42222 = n42238 & n39955;
  assign n42215 = ~n42242;
  assign n42169 = ~n42238;
  assign n42202 = n42262 ^ n42263;
  assign n42254 = n42275 & n42276;
  assign n40528 = n42161 ^ n42162;
  assign n42163 = ~n42173;
  assign n42164 = ~n42162;
  assign n42160 = n42188 ^ n42189;
  assign n42186 = ~n42197;
  assign n42191 = ~n42188;
  assign n42166 = ~n42198;
  assign n42195 = n38500 & n40006;
  assign n42196 = n38500 & n40967;
  assign n42214 = ~n42221;
  assign n42217 = n42169 & n39930;
  assign n42194 = ~n42222;
  assign n42223 = n42254 ^ n42255;
  assign n42256 = ~n42254;
  assign n41758 = ~n40528;
  assign n42120 = n42159 ^ n42160;
  assign n42112 = n42164 & n42161;
  assign n42174 = n42186 & n42187;
  assign n42175 = n42190 & n42191;
  assign n41043 = ~n42195;
  assign n42176 = ~n42196;
  assign n42192 = n42214 & n42215;
  assign n42171 = ~n42217;
  assign n42200 = n89 ^ n42223;
  assign n42243 = n42256 & n42257;
  assign n42140 = n42120 & n227;
  assign n42115 = ~n42112;
  assign n42139 = ~n42120;
  assign n42153 = ~n42174;
  assign n42165 = ~n42175;
  assign n42123 = n42176 & n42177;
  assign n42168 = n42192 ^ n39955;
  assign n42193 = ~n42192;
  assign n42127 = n42199 ^ n42200;
  assign n42181 = n42200 & n42199;
  assign n42224 = ~n42243;
  assign n42134 = n42139 & n19695;
  assign n42103 = ~n42140;
  assign n42133 = n42153 ^ n42154;
  assign n42152 = n42163 & n42153;
  assign n42141 = n42165 & n42166;
  assign n42156 = n42123 & n42167;
  assign n38435 = n42168 ^ n42169;
  assign n42155 = ~n42123;
  assign n42178 = n42193 & n42194;
  assign n42179 = n42127 & n39836;
  assign n42180 = ~n42127;
  assign n42201 = n42224 & n42225;
  assign n42113 = n228 ^ n42133;
  assign n42121 = ~n42134;
  assign n42124 = n42141 ^ n42142;
  assign n42145 = n38435 & n40905;
  assign n42146 = n38435 & n39955;
  assign n42137 = ~n42152;
  assign n42144 = ~n42141;
  assign n42150 = n42155 & n42142;
  assign n42143 = ~n42156;
  assign n38465 = ~n38435;
  assign n42170 = ~n42178;
  assign n42149 = ~n42179;
  assign n42172 = n42180 & n39892;
  assign n42182 = n42201 ^ n42202;
  assign n40493 = n42112 ^ n42113;
  assign n42086 = n42123 ^ n42124;
  assign n42114 = ~n42113;
  assign n42119 = n42137 & n42138;
  assign n42135 = n42143 & n42144;
  assign n42131 = ~n42145;
  assign n40942 = ~n42146;
  assign n42126 = ~n42150;
  assign n42147 = n42170 & n42171;
  assign n42130 = ~n42172;
  assign n42089 = n42181 ^ n42182;
  assign n41721 = ~n40493;
  assign n42105 = n42086 & n226;
  assign n42083 = n42114 & n42115;
  assign n42104 = ~n42086;
  assign n42101 = n42119 ^ n42120;
  assign n42077 = n42131 & n42132;
  assign n42122 = ~n42119;
  assign n42125 = ~n42135;
  assign n42128 = n42147 ^ n39836;
  assign n42148 = ~n42147;
  assign n42157 = n42089 & n39788;
  assign n42158 = ~n42089;
  assign n42084 = n227 ^ n42101;
  assign n42094 = n42104 & n19641;
  assign n42067 = ~n42105;
  assign n42111 = n42077 & n42117;
  assign n42116 = n42121 & n42122;
  assign n42110 = ~n42077;
  assign n42118 = n42125 & n42126;
  assign n38412 = n42127 ^ n42128;
  assign n42136 = n42148 & n42149;
  assign n42092 = ~n42157;
  assign n42151 = n42158 & n39766;
  assign n40428 = n42083 ^ n42084;
  assign n42041 = n42084 & n42083;
  assign n42081 = ~n42094;
  assign n42106 = n42110 & n42097;
  assign n42095 = ~n42111;
  assign n42102 = ~n42116;
  assign n42096 = ~n42118;
  assign n38439 = ~n38412;
  assign n42129 = ~n42136;
  assign n42109 = ~n42151;
  assign n41684 = ~n40428;
  assign n42044 = ~n42041;
  assign n42093 = n42095 & n42096;
  assign n42078 = n42096 ^ n42097;
  assign n42085 = n42102 & n42103;
  assign n42080 = ~n42106;
  assign n42098 = n38439 & n39836;
  assign n42099 = n38439 & n40860;
  assign n42107 = n42129 & n42130;
  assign n42046 = n42077 ^ n42078;
  assign n42065 = n42085 ^ n42086;
  assign n42079 = ~n42093;
  assign n42082 = ~n42085;
  assign n40899 = ~n42098;
  assign n42087 = ~n42099;
  assign n42090 = n42107 ^ n39766;
  assign n42108 = ~n42107;
  assign n42042 = n226 ^ n42065;
  assign n42059 = n42046 & n19596;
  assign n42060 = ~n42046;
  assign n42061 = n42079 & n42080;
  assign n42076 = n42081 & n42082;
  assign n42037 = n42087 & n42088;
  assign n38381 = n42089 ^ n42090;
  assign n42100 = n42108 & n42109;
  assign n40379 = n42041 ^ n42042;
  assign n42043 = ~n42042;
  assign n42047 = ~n42059;
  assign n42054 = n42060 & n225;
  assign n42038 = n42061 ^ n42062;
  assign n42058 = ~n42061;
  assign n42069 = n38381 & n39766;
  assign n42070 = n42037 & n42075;
  assign n42071 = n38381 & n40780;
  assign n42066 = ~n42076;
  assign n42068 = ~n42037;
  assign n38403 = ~n38381;
  assign n42091 = ~n42100;
  assign n41645 = ~n40379;
  assign n42008 = n42037 ^ n42038;
  assign n42003 = n42043 & n42044;
  assign n42028 = ~n42054;
  assign n42045 = n42066 & n42067;
  assign n42063 = n42068 & n42062;
  assign n40811 = ~n42069;
  assign n42057 = ~n42070;
  assign n42055 = ~n42071;
  assign n42072 = n42091 & n42092;
  assign n42022 = n42008 & n224;
  assign n42021 = ~n42008;
  assign n42006 = ~n42003;
  assign n42026 = n42045 ^ n42046;
  assign n41997 = n42055 & n42056;
  assign n42049 = n42057 & n42058;
  assign n42048 = ~n42045;
  assign n42034 = ~n42063;
  assign n42051 = n42072 ^ n39682;
  assign n42073 = ~n42072;
  assign n42016 = n42021 & n19565;
  assign n41984 = ~n42022;
  assign n42004 = n225 ^ n42026;
  assign n42036 = n41997 & n42040;
  assign n42039 = n42047 & n42048;
  assign n42035 = ~n41997;
  assign n42033 = ~n42049;
  assign n38346 = n42050 ^ n42051;
  assign n42064 = n42073 & n42074;
  assign n41606 = n42003 ^ n42004;
  assign n42001 = ~n42016;
  assign n42005 = ~n42004;
  assign n42017 = n42033 & n42034;
  assign n42029 = n42035 & n42018;
  assign n42019 = ~n42036;
  assign n42027 = ~n42039;
  assign n38371 = ~n38346;
  assign n42052 = ~n42064;
  assign n40333 = ~n41606;
  assign n41967 = n42005 & n42006;
  assign n41998 = n42017 ^ n42018;
  assign n42007 = n42027 & n42028;
  assign n42020 = ~n42017;
  assign n42000 = ~n42029;
  assign n42023 = n38371 & n39707;
  assign n42024 = n38371 & n40715;
  assign n42030 = n42052 & n42053;
  assign n41966 = n41997 ^ n41998;
  assign n41989 = n42007 ^ n42008;
  assign n42009 = n42019 & n42020;
  assign n42002 = ~n42007;
  assign n40756 = ~n42023;
  assign n42010 = ~n42024;
  assign n42013 = n42030 ^ n39582;
  assign n42031 = ~n42030;
  assign n41978 = n41966 & n239;
  assign n41968 = n224 ^ n41989;
  assign n41977 = ~n41966;
  assign n41996 = n42001 & n42002;
  assign n41999 = ~n42009;
  assign n41960 = n42010 & n42011;
  assign n38309 = n42012 ^ n42013;
  assign n42025 = n42031 & n42032;
  assign n40272 = n41967 ^ n41968;
  assign n41927 = n41968 & n41967;
  assign n41969 = n41977 & n19533;
  assign n41937 = ~n41978;
  assign n41983 = ~n41996;
  assign n41979 = n41999 & n42000;
  assign n41992 = n41960 & n41980;
  assign n41990 = ~n41960;
  assign n38344 = ~n38309;
  assign n42014 = ~n42025;
  assign n41556 = ~n40272;
  assign n41930 = ~n41927;
  assign n41959 = ~n41969;
  assign n41961 = n41979 ^ n41980;
  assign n41965 = n41983 & n41984;
  assign n41982 = ~n41979;
  assign n41985 = n41990 & n41991;
  assign n41986 = n38344 & n39582;
  assign n41987 = n38344 & n40685;
  assign n41981 = ~n41992;
  assign n41993 = n42014 & n42015;
  assign n41916 = n41960 ^ n41961;
  assign n41947 = n41965 ^ n41966;
  assign n41958 = ~n41965;
  assign n41972 = n41981 & n41982;
  assign n41963 = ~n41985;
  assign n40707 = ~n41986;
  assign n41970 = ~n41987;
  assign n41974 = n41993 ^ n39516;
  assign n41994 = ~n41993;
  assign n41928 = n239 ^ n41947;
  assign n41938 = n41916 & n19483;
  assign n41939 = ~n41916;
  assign n41950 = n41958 & n41959;
  assign n41941 = n41970 & n41971;
  assign n41962 = ~n41972;
  assign n38270 = n41973 ^ n41974;
  assign n41988 = n41994 & n41995;
  assign n40205 = n41927 ^ n41928;
  assign n41929 = ~n41928;
  assign n41918 = ~n41938;
  assign n41932 = n41939 & n238;
  assign n41936 = ~n41950;
  assign n41940 = n41962 & n41963;
  assign n41953 = n38270 & n39516;
  assign n41954 = n38270 & n40636;
  assign n41955 = n41941 & n41920;
  assign n41951 = ~n41941;
  assign n38299 = ~n38270;
  assign n41975 = ~n41988;
  assign n41527 = ~n40205;
  assign n41880 = n41929 & n41930;
  assign n41901 = ~n41932;
  assign n41915 = n41936 & n41937;
  assign n41919 = n41940 ^ n41941;
  assign n41945 = ~n41940;
  assign n41948 = n41951 & n41952;
  assign n40676 = ~n41953;
  assign n41942 = ~n41954;
  assign n41944 = ~n41955;
  assign n41964 = n41975 & n41976;
  assign n41879 = ~n41880;
  assign n41899 = n41915 ^ n41916;
  assign n41883 = n41919 ^ n41920;
  assign n41917 = ~n41915;
  assign n41886 = n41942 & n41943;
  assign n41933 = n41944 & n41945;
  assign n41922 = ~n41948;
  assign n41957 = n41964 & n39433;
  assign n41956 = ~n41964;
  assign n41881 = n238 ^ n41899;
  assign n41902 = n41883 & n19432;
  assign n41903 = ~n41883;
  assign n41911 = n41917 & n41918;
  assign n41924 = n41886 & n41931;
  assign n41923 = ~n41886;
  assign n41921 = ~n41933;
  assign n41949 = n41956 & n39435;
  assign n41935 = ~n41957;
  assign n40131 = n41880 ^ n41881;
  assign n41878 = ~n41881;
  assign n41885 = ~n41902;
  assign n41896 = n41903 & n237;
  assign n41900 = ~n41911;
  assign n41904 = n41921 & n41922;
  assign n41912 = n41923 & n41905;
  assign n41907 = ~n41924;
  assign n41934 = n41935 & n41946;
  assign n41926 = ~n41949;
  assign n41487 = ~n40131;
  assign n41840 = n41878 & n41879;
  assign n41867 = ~n41896;
  assign n41882 = n41900 & n41901;
  assign n41887 = n41904 ^ n41905;
  assign n41906 = ~n41904;
  assign n41889 = ~n41912;
  assign n41925 = ~n41934;
  assign n41913 = n41926 & n41935;
  assign n41856 = ~n41840;
  assign n41865 = n41882 ^ n41883;
  assign n41843 = n41886 ^ n41887;
  assign n41884 = ~n41882;
  assign n41897 = n41906 & n41907;
  assign n38230 = n41913 ^ n41914;
  assign n41908 = n41925 & n41926;
  assign n41841 = n237 ^ n41865;
  assign n41869 = n41843 & n236;
  assign n41868 = ~n41843;
  assign n41875 = n41884 & n41885;
  assign n41888 = ~n41897;
  assign n41891 = n41908 ^ n39405;
  assign n38261 = ~n38230;
  assign n41909 = ~n41908;
  assign n40099 = n41840 ^ n41841;
  assign n41805 = n41841 & n41856;
  assign n41858 = n41868 & n19414;
  assign n41825 = ~n41869;
  assign n41866 = ~n41875;
  assign n41870 = n41888 & n41889;
  assign n38192 = n41890 ^ n41891;
  assign n41894 = n38261 & n40602;
  assign n41895 = n38261 & n39433;
  assign n41898 = n41909 & n41910;
  assign n41439 = ~n40099;
  assign n41845 = ~n41858;
  assign n41842 = n41866 & n41867;
  assign n41847 = n41870 ^ n41871;
  assign n41853 = ~n41870;
  assign n38228 = ~n38192;
  assign n41876 = ~n41894;
  assign n40630 = ~n41895;
  assign n41892 = ~n41898;
  assign n41823 = n41842 ^ n41843;
  assign n41844 = ~n41842;
  assign n41859 = n38228 & n40552;
  assign n41860 = n38228 & n39356;
  assign n41846 = n41876 & n41877;
  assign n41872 = n41892 & n41893;
  assign n41806 = n236 ^ n41823;
  assign n41838 = n41844 & n41845;
  assign n41809 = n41846 ^ n41847;
  assign n41848 = ~n41859;
  assign n40590 = ~n41860;
  assign n41863 = n41846 & n41871;
  assign n41851 = n41872 ^ n39299;
  assign n41861 = ~n41846;
  assign n41873 = ~n41872;
  assign n40026 = n41805 ^ n41806;
  assign n41807 = ~n41806;
  assign n41826 = n41809 & n19360;
  assign n41824 = ~n41838;
  assign n41827 = ~n41809;
  assign n41781 = n41848 & n41849;
  assign n38190 = n41850 ^ n41851;
  assign n41857 = n41861 & n41862;
  assign n41852 = ~n41863;
  assign n41864 = n41873 & n41874;
  assign n41381 = ~n40026;
  assign n41768 = n41807 & n41805;
  assign n41808 = n41824 & n41825;
  assign n41811 = ~n41826;
  assign n41819 = n41827 & n235;
  assign n41830 = n41781 & n41804;
  assign n41831 = n38190 & n40523;
  assign n41832 = n38190 & n39299;
  assign n41828 = ~n41781;
  assign n38153 = ~n38190;
  assign n41839 = n41852 & n41853;
  assign n41834 = ~n41857;
  assign n41854 = ~n41864;
  assign n41787 = n41808 ^ n41809;
  assign n41810 = ~n41808;
  assign n41789 = ~n41819;
  assign n41820 = n41828 & n41829;
  assign n41812 = ~n41830;
  assign n41817 = ~n41831;
  assign n40539 = ~n41832;
  assign n41833 = ~n41839;
  assign n41835 = n41854 & n41855;
  assign n41769 = n235 ^ n41787;
  assign n41800 = n41810 & n41811;
  assign n41749 = n41817 & n41818;
  assign n41791 = ~n41820;
  assign n41821 = n41833 & n41834;
  assign n41814 = n41835 ^ n39336;
  assign n41836 = ~n41835;
  assign n39905 = n41768 ^ n41769;
  assign n41726 = n41769 & n41768;
  assign n41788 = ~n41800;
  assign n41798 = n41749 & n41801;
  assign n41797 = ~n41749;
  assign n38112 = n41813 ^ n41814;
  assign n41803 = ~n41821;
  assign n41822 = n41836 & n41837;
  assign n41308 = ~n39905;
  assign n41770 = n41788 & n41789;
  assign n41792 = n41797 & n41772;
  assign n41775 = ~n41798;
  assign n41793 = n38112 & n41799;
  assign n38151 = ~n38112;
  assign n41782 = n41803 ^ n41804;
  assign n41802 = n41812 & n41803;
  assign n41815 = ~n41822;
  assign n41751 = n234 ^ n41770;
  assign n41743 = ~n41770;
  assign n41752 = n41781 ^ n41782;
  assign n41754 = ~n41792;
  assign n41783 = n38151 & n40489;
  assign n40559 = ~n41793;
  assign n41784 = n38151 & n40542;
  assign n41785 = n38151 & n39260;
  assign n41790 = ~n41802;
  assign n41794 = n41815 & n41816;
  assign n41727 = n41751 ^ n41752;
  assign n41766 = n41752 & n234;
  assign n41765 = ~n41752;
  assign n41773 = ~n41783;
  assign n40544 = ~n41784;
  assign n40505 = ~n41785;
  assign n41771 = n41790 & n41791;
  assign n41778 = n41794 ^ n39197;
  assign n41795 = ~n41794;
  assign n39827 = n41726 ^ n41727;
  assign n41728 = ~n41727;
  assign n41764 = n41765 & n19316;
  assign n41724 = ~n41766;
  assign n41750 = n41771 ^ n41772;
  assign n41708 = n41773 & n41774;
  assign n38073 = n41777 ^ n41778;
  assign n41776 = ~n41771;
  assign n41786 = n41795 & n41796;
  assign n41242 = ~n39827;
  assign n41661 = n41728 & n41726;
  assign n41701 = n41749 ^ n41750;
  assign n41742 = ~n41764;
  assign n41757 = n41708 & n41732;
  assign n41759 = n38073 & n40528;
  assign n41755 = ~n41708;
  assign n38110 = ~n38073;
  assign n41767 = n41775 & n41776;
  assign n41779 = ~n41786;
  assign n41730 = n41701 & n233;
  assign n41729 = ~n41701;
  assign n41741 = n41742 & n41743;
  assign n41744 = n41755 & n41756;
  assign n41735 = ~n41757;
  assign n41745 = n38110 & n39197;
  assign n41746 = n38110 & n40454;
  assign n41747 = n38110 & n41758;
  assign n40530 = ~n41759;
  assign n41753 = ~n41767;
  assign n41760 = n41779 & n41780;
  assign n41722 = n41729 & n19279;
  assign n41686 = ~n41730;
  assign n41723 = ~n41741;
  assign n41711 = ~n41744;
  assign n40476 = ~n41745;
  assign n41733 = ~n41746;
  assign n40510 = ~n41747;
  assign n41731 = n41753 & n41754;
  assign n41737 = n41760 ^ n41761;
  assign n41762 = ~n41760;
  assign n41704 = ~n41722;
  assign n41720 = n41723 & n41724;
  assign n41709 = n41731 ^ n41732;
  assign n41692 = n41733 & n41734;
  assign n38015 = n39227 ^ n41737;
  assign n41738 = n41737 & n39159;
  assign n41736 = ~n41731;
  assign n41748 = n41762 & n41763;
  assign n41668 = n41708 ^ n41709;
  assign n41700 = ~n41720;
  assign n41714 = n38015 & n40410;
  assign n41715 = n41692 & n41674;
  assign n41716 = n38015 & n41721;
  assign n41712 = ~n41692;
  assign n38071 = ~n38015;
  assign n41725 = n41735 & n41736;
  assign n40433 = ~n41738;
  assign n41739 = ~n41748;
  assign n41689 = n41668 & n19255;
  assign n41683 = n41700 ^ n41701;
  assign n41699 = n41704 & n41700;
  assign n41690 = ~n41668;
  assign n41705 = n41712 & n41713;
  assign n41702 = ~n41714;
  assign n41693 = ~n41715;
  assign n40472 = ~n41716;
  assign n41706 = n38071 & n40493;
  assign n41710 = ~n41725;
  assign n41717 = n41739 & n41740;
  assign n41662 = n233 ^ n41683;
  assign n41670 = ~n41689;
  assign n41687 = n41690 & n232;
  assign n41685 = ~n41699;
  assign n41632 = n41702 & n41703;
  assign n41676 = ~n41705;
  assign n40495 = ~n41706;
  assign n41691 = n41710 & n41711;
  assign n41696 = n41717 ^ n39192;
  assign n41718 = ~n41717;
  assign n39754 = n41661 ^ n41662;
  assign n41623 = n41662 & n41661;
  assign n41667 = n41685 & n41686;
  assign n41647 = ~n41687;
  assign n41673 = n41691 ^ n41692;
  assign n41641 = ~n41632;
  assign n37978 = n41695 ^ n41696;
  assign n41694 = ~n41691;
  assign n41707 = n41718 & n41719;
  assign n41173 = ~n39754;
  assign n41648 = n41667 ^ n41668;
  assign n41608 = n41673 ^ n41674;
  assign n41669 = ~n41667;
  assign n41677 = n37978 & n40330;
  assign n41678 = n37978 & n41684;
  assign n41679 = n37978 & n39125;
  assign n38026 = ~n37978;
  assign n41688 = n41693 & n41694;
  assign n41697 = ~n41707;
  assign n41624 = n232 ^ n41648;
  assign n41651 = n41608 & n19197;
  assign n41663 = n41669 & n41670;
  assign n41652 = ~n41608;
  assign n41671 = n38026 & n40428;
  assign n41664 = ~n41677;
  assign n40431 = ~n41678;
  assign n40387 = ~n41679;
  assign n41675 = ~n41688;
  assign n41680 = n41697 & n41698;
  assign n39679 = n41623 ^ n41624;
  assign n41581 = n41624 & n41623;
  assign n41627 = ~n41651;
  assign n41649 = n41652 & n247;
  assign n41646 = ~n41663;
  assign n41576 = n41664 & n41665;
  assign n40449 = ~n41671;
  assign n41653 = n41675 & n41676;
  assign n41658 = n41680 ^ n39105;
  assign n41681 = ~n41680;
  assign n41091 = ~n39679;
  assign n41584 = ~n41581;
  assign n41625 = n41646 & n41647;
  assign n41610 = ~n41649;
  assign n41644 = n41576 & n41602;
  assign n41633 = n41653 ^ n41654;
  assign n41642 = ~n41576;
  assign n37959 = n41657 ^ n41658;
  assign n41656 = n41653 & n41666;
  assign n41655 = ~n41653;
  assign n41672 = n41681 & n41682;
  assign n41607 = n247 ^ n41625;
  assign n41586 = n41632 ^ n41633;
  assign n41626 = ~n41625;
  assign n41635 = n41642 & n41643;
  assign n41604 = ~n41644;
  assign n41636 = n37959 & n41645;
  assign n37989 = ~n37959;
  assign n41650 = n41655 & n41654;
  assign n41640 = ~n41656;
  assign n41659 = ~n41672;
  assign n41582 = n41607 ^ n41608;
  assign n41613 = n41586 & n246;
  assign n41620 = n41626 & n41627;
  assign n41612 = ~n41586;
  assign n41580 = ~n41635;
  assign n41628 = n37989 & n40315;
  assign n41629 = n37989 & n40379;
  assign n40406 = ~n41636;
  assign n41630 = n37989 & n39117;
  assign n41634 = n41640 & n41641;
  assign n41622 = ~n41650;
  assign n41637 = n41659 & n41660;
  assign n39603 = n41581 ^ n41582;
  assign n41583 = ~n41582;
  assign n41611 = n41612 & n19179;
  assign n41569 = ~n41613;
  assign n41609 = ~n41620;
  assign n41614 = ~n41628;
  assign n40382 = ~n41629;
  assign n40344 = ~n41630;
  assign n41621 = ~n41634;
  assign n41617 = n41637 ^ n39128;
  assign n41638 = ~n41637;
  assign n41035 = ~n39603;
  assign n40994 = n41583 & n41584;
  assign n41585 = n41609 & n41610;
  assign n41588 = ~n41611;
  assign n41538 = n41614 & n41615;
  assign n37918 = n41616 ^ n41617;
  assign n41601 = n41621 & n41622;
  assign n41631 = n41638 & n41639;
  assign n41567 = n41585 ^ n41586;
  assign n41587 = ~n41585;
  assign n41577 = n41601 ^ n41602;
  assign n41596 = n41538 & n41605;
  assign n41597 = n37918 & n41606;
  assign n41595 = ~n41538;
  assign n37949 = ~n37918;
  assign n41603 = ~n41601;
  assign n41618 = ~n41631;
  assign n40955 = n246 ^ n41567;
  assign n41545 = n41576 ^ n41577;
  assign n41578 = n41587 & n41588;
  assign n41589 = n41595 & n41563;
  assign n41590 = n37949 & n40187;
  assign n41565 = ~n41596;
  assign n41591 = n37949 & n39062;
  assign n40361 = ~n41597;
  assign n41592 = n37949 & n40333;
  assign n41594 = n41603 & n41604;
  assign n41598 = n41618 & n41619;
  assign n41502 = n40955 & n40994;
  assign n41560 = n41545 & n19125;
  assign n41561 = ~n41545;
  assign n41568 = ~n41578;
  assign n41541 = ~n41589;
  assign n41570 = ~n41590;
  assign n40286 = ~n41591;
  assign n40336 = ~n41592;
  assign n41579 = ~n41594;
  assign n41573 = n41598 ^ n39028;
  assign n41599 = ~n41598;
  assign n41542 = ~n41560;
  assign n41551 = n41561 & n245;
  assign n41544 = n41568 & n41569;
  assign n41498 = n41570 & n41571;
  assign n37881 = n41572 ^ n41573;
  assign n41562 = n41579 & n41580;
  assign n41593 = n41599 & n41600;
  assign n41528 = n41544 ^ n41545;
  assign n41530 = ~n41551;
  assign n41543 = ~n41544;
  assign n41539 = n41562 ^ n41563;
  assign n41554 = n41498 & n41566;
  assign n41555 = n37881 & n40272;
  assign n41553 = ~n41498;
  assign n37909 = ~n37881;
  assign n41564 = ~n41562;
  assign n41574 = ~n41593;
  assign n41503 = n245 ^ n41528;
  assign n41506 = n41538 ^ n41539;
  assign n41537 = n41542 & n41543;
  assign n41546 = n41553 & n41524;
  assign n41547 = n37909 & n40169;
  assign n41526 = ~n41554;
  assign n40303 = ~n41555;
  assign n41548 = n37909 & n39028;
  assign n41549 = n37909 & n41556;
  assign n41552 = n41564 & n41565;
  assign n41557 = n41574 & n41575;
  assign n38672 = n41502 ^ n41503;
  assign n41504 = ~n41503;
  assign n41522 = n41506 & n244;
  assign n41521 = ~n41506;
  assign n41529 = ~n41537;
  assign n41501 = ~n41546;
  assign n41531 = ~n41547;
  assign n40204 = ~n41548;
  assign n40275 = ~n41549;
  assign n41540 = ~n41552;
  assign n41533 = n41557 ^ n38996;
  assign n41558 = ~n41557;
  assign n37741 = n38672 ^ n38663;
  assign n41383 = n38672 & n38663;
  assign n41463 = n41504 & n41502;
  assign n41512 = n41521 & n19082;
  assign n41479 = ~n41522;
  assign n41505 = n41529 & n41530;
  assign n41456 = n41531 & n41532;
  assign n37843 = n41533 ^ n41534;
  assign n41523 = n41540 & n41541;
  assign n41550 = n41558 & n41559;
  assign n41462 = n37741 & n40478;
  assign n41488 = n41505 ^ n41506;
  assign n41497 = ~n41512;
  assign n41496 = ~n41505;
  assign n41499 = n41523 ^ n41524;
  assign n41516 = n41456 & n41483;
  assign n41517 = n37843 & n41527;
  assign n41514 = ~n41456;
  assign n37879 = ~n37843;
  assign n41525 = ~n41523;
  assign n41535 = ~n41550;
  assign n41444 = ~n41462;
  assign n41464 = n244 ^ n41488;
  assign n41489 = n41496 & n41497;
  assign n41455 = n41498 ^ n41499;
  assign n41507 = n41514 & n41515;
  assign n41485 = ~n41516;
  assign n41508 = n37879 & n40044;
  assign n40237 = ~n41517;
  assign n41509 = n37879 & n38996;
  assign n41510 = n37879 & n40205;
  assign n41513 = n41525 & n41526;
  assign n41518 = n41535 & n41536;
  assign n41412 = n41444 & n41445;
  assign n41446 = n41463 ^ n41464;
  assign n41396 = n41464 & n41463;
  assign n41481 = n41455 & n243;
  assign n41478 = ~n41489;
  assign n41480 = ~n41455;
  assign n41461 = ~n41507;
  assign n41490 = ~n41508;
  assign n40148 = ~n41509;
  assign n40208 = ~n41510;
  assign n41500 = ~n41513;
  assign n41493 = n41518 ^ n38937;
  assign n41519 = ~n41518;
  assign n41385 = n41412 ^ n41413;
  assign n41414 = ~n41412;
  assign n41441 = n41446 & n38621;
  assign n41440 = ~n41446;
  assign n41399 = ~n41396;
  assign n41454 = n41478 & n41479;
  assign n41468 = n41480 & n19042;
  assign n41429 = ~n41481;
  assign n41394 = n41490 & n41491;
  assign n37841 = n41492 ^ n41493;
  assign n41482 = n41500 & n41501;
  assign n41511 = n41519 & n41520;
  assign n39154 = n391 ^ n41385;
  assign n41126 = n41385 & n391;
  assign n41236 = n41414 & n41415;
  assign n41426 = n41440 & n38626;
  assign n41409 = ~n41441;
  assign n41427 = n41454 ^ n41455;
  assign n41452 = ~n41454;
  assign n41453 = ~n41468;
  assign n41457 = n41482 ^ n41483;
  assign n41471 = n37841 & n39967;
  assign n41472 = n41394 & n41486;
  assign n41473 = n37841 & n41487;
  assign n41474 = n37841 & n38937;
  assign n41470 = ~n41394;
  assign n37802 = ~n37841;
  assign n41484 = ~n41482;
  assign n41494 = ~n41511;
  assign n40300 = ~n39154;
  assign n41408 = n41409 & n41383;
  assign n41387 = ~n41426;
  assign n41397 = n243 ^ n41427;
  assign n41447 = n41452 & n41453;
  assign n41401 = n41456 ^ n41457;
  assign n41465 = n41470 & n41433;
  assign n41458 = ~n41471;
  assign n41435 = ~n41472;
  assign n40134 = ~n41473;
  assign n41466 = n37802 & n40131;
  assign n40077 = ~n41474;
  assign n41469 = n41484 & n41485;
  assign n41475 = n41494 & n41495;
  assign n41330 = n41396 ^ n41397;
  assign n41386 = ~n41408;
  assign n41382 = n41387 & n41409;
  assign n41398 = ~n41397;
  assign n41430 = n41401 & n19000;
  assign n41428 = ~n41447;
  assign n41431 = ~n41401;
  assign n41442 = n41458 & n41459;
  assign n41407 = ~n41465;
  assign n40176 = ~n41466;
  assign n41460 = ~n41469;
  assign n41448 = n41475 ^ n38955;
  assign n41476 = ~n41475;
  assign n37542 = n41382 ^ n41383;
  assign n41369 = n41330 & n38589;
  assign n41357 = n41386 & n41387;
  assign n41370 = ~n41330;
  assign n41344 = n41398 & n41399;
  assign n41400 = n41428 & n41429;
  assign n41403 = ~n41430;
  assign n41416 = n41431 & n242;
  assign n41438 = n41442 & n41443;
  assign n41436 = ~n41442;
  assign n37763 = n41448 ^ n41449;
  assign n41432 = n41460 & n41461;
  assign n41467 = n41476 & n41477;
  assign n41354 = n37542 & n40290;
  assign n41331 = n41357 ^ n38611;
  assign n37714 = ~n37542;
  assign n41315 = ~n41369;
  assign n41358 = n41370 & n38611;
  assign n41342 = ~n41357;
  assign n41347 = ~n41344;
  assign n41371 = n41400 ^ n41401;
  assign n41402 = ~n41400;
  assign n41373 = ~n41416;
  assign n41395 = n41432 ^ n41433;
  assign n41418 = n41436 & n41437;
  assign n41377 = ~n41438;
  assign n41419 = n37763 & n39965;
  assign n41420 = n37763 & n38955;
  assign n41421 = n37763 & n41439;
  assign n37792 = ~n37763;
  assign n41434 = ~n41432;
  assign n41450 = ~n41467;
  assign n37532 = n41330 ^ n41331;
  assign n41332 = ~n41354;
  assign n41343 = ~n41358;
  assign n41345 = n242 ^ n41371;
  assign n41384 = n41394 ^ n41395;
  assign n41388 = n41402 & n41403;
  assign n41351 = ~n41418;
  assign n41404 = ~n41419;
  assign n40002 = ~n41420;
  assign n40061 = ~n41421;
  assign n41410 = n37792 & n40099;
  assign n41417 = n41434 & n41435;
  assign n41422 = n41450 & n41451;
  assign n41300 = n37532 & n40264;
  assign n37530 = ~n37532;
  assign n41312 = n41332 & n41333;
  assign n41334 = n41342 & n41343;
  assign n41254 = n41344 ^ n41345;
  assign n41346 = ~n41345;
  assign n41375 = n41384 & n241;
  assign n41372 = ~n41388;
  assign n41374 = ~n41384;
  assign n41323 = n41404 & n41405;
  assign n41389 = n41351 & n41377;
  assign n40101 = ~n41410;
  assign n41406 = ~n41417;
  assign n41390 = n41422 ^ n41423;
  assign n41424 = ~n41422;
  assign n41278 = ~n41300;
  assign n41301 = n41312 & n41313;
  assign n41298 = ~n41312;
  assign n41316 = n41254 & n38563;
  assign n41314 = ~n41334;
  assign n41317 = ~n41254;
  assign n41283 = n41346 & n41347;
  assign n41319 = n41372 & n41373;
  assign n41359 = n41374 & n18956;
  assign n41321 = ~n41375;
  assign n41380 = n41323 & n41290;
  assign n41378 = ~n41323;
  assign n41361 = ~n41389;
  assign n37690 = n38853 ^ n41390;
  assign n41360 = n41406 & n41407;
  assign n41391 = n41390 & n38940;
  assign n41411 = n41424 & n41425;
  assign n41163 = n41278 & n41279;
  assign n41295 = n41298 & n41299;
  assign n41271 = ~n41301;
  assign n41280 = n41314 & n41315;
  assign n41282 = ~n41316;
  assign n41302 = n41317 & n38585;
  assign n41348 = ~n41319;
  assign n41349 = ~n41359;
  assign n41286 = n41360 ^ n41361;
  assign n41363 = n41378 & n41379;
  assign n41325 = ~n41380;
  assign n41364 = n37690 & n39781;
  assign n41365 = n37690 & n41381;
  assign n37761 = ~n37690;
  assign n41376 = ~n41360;
  assign n39926 = ~n41391;
  assign n41392 = ~n41411;
  assign n41251 = n41163 & n41204;
  assign n41249 = ~n41163;
  assign n41270 = n41271 & n41236;
  assign n41255 = n41280 ^ n38563;
  assign n41253 = ~n41295;
  assign n41281 = ~n41280;
  assign n41248 = ~n41302;
  assign n41335 = n41348 & n41349;
  assign n41318 = n41349 & n41321;
  assign n41337 = n41286 & n240;
  assign n41336 = ~n41286;
  assign n41294 = ~n41363;
  assign n41352 = ~n41364;
  assign n41355 = n37761 & n40026;
  assign n39985 = ~n41365;
  assign n41362 = n41376 & n41377;
  assign n41366 = n41392 & n41393;
  assign n41234 = n41249 & n41250;
  assign n41216 = ~n41251;
  assign n37437 = n41254 ^ n41255;
  assign n41252 = ~n41270;
  assign n41235 = n41253 & n41271;
  assign n41272 = n41281 & n41282;
  assign n41284 = n41318 ^ n41319;
  assign n41320 = ~n41335;
  assign n41329 = n41336 & n18899;
  assign n41260 = ~n41337;
  assign n41226 = n41352 & n41353;
  assign n40028 = ~n41355;
  assign n41350 = ~n41362;
  assign n41338 = n41366 ^ n38906;
  assign n41367 = ~n41366;
  assign n41181 = ~n41234;
  assign n41217 = n41235 ^ n41236;
  assign n37455 = ~n37437;
  assign n41237 = n41252 & n41253;
  assign n41247 = ~n41272;
  assign n41182 = n41283 ^ n41284;
  assign n41219 = n41284 & n41283;
  assign n41285 = n41320 & n41321;
  assign n41288 = ~n41329;
  assign n41328 = n41226 & n41264;
  assign n41326 = ~n41226;
  assign n37642 = n41338 ^ n41339;
  assign n41322 = n41350 & n41351;
  assign n41356 = n41367 & n41368;
  assign n41202 = n41217 & n390;
  assign n41205 = n37455 & n40267;
  assign n41201 = ~n41217;
  assign n41203 = ~n41237;
  assign n41218 = n41247 & n41248;
  assign n41257 = n41182 & n38532;
  assign n41256 = ~n41182;
  assign n41222 = ~n41219;
  assign n41258 = n41285 ^ n41286;
  assign n41287 = ~n41285;
  assign n41289 = n41322 ^ n41323;
  assign n41304 = n41326 & n41327;
  assign n41305 = n37642 & n39673;
  assign n41265 = ~n41328;
  assign n41306 = n37642 & n39905;
  assign n41307 = n37642 & n38906;
  assign n37720 = ~n37642;
  assign n41324 = ~n41322;
  assign n41340 = ~n41356;
  assign n41199 = n41201 & n16646;
  assign n41128 = ~n41202;
  assign n41164 = n41203 ^ n41204;
  assign n41178 = ~n41205;
  assign n41200 = n41216 & n41203;
  assign n41183 = n41218 ^ n38552;
  assign n41214 = ~n41218;
  assign n41238 = n41256 & n38552;
  assign n41215 = ~n41257;
  assign n41220 = n240 ^ n41258;
  assign n41273 = n41287 & n41288;
  assign n41189 = n41289 ^ n41290;
  assign n41229 = ~n41304;
  assign n41291 = ~n41305;
  assign n39907 = ~n41306;
  assign n39849 = ~n41307;
  assign n41296 = n37720 & n41308;
  assign n41303 = n41324 & n41325;
  assign n41309 = n41340 & n41341;
  assign n41077 = n41163 ^ n41164;
  assign n41097 = n41178 & n41179;
  assign n37379 = n41182 ^ n41183;
  assign n41165 = ~n41199;
  assign n41180 = ~n41200;
  assign n41206 = n41214 & n41215;
  assign n41100 = n41219 ^ n41220;
  assign n41185 = ~n41238;
  assign n41221 = ~n41220;
  assign n41261 = n41189 & n18888;
  assign n41259 = ~n41273;
  assign n41262 = ~n41189;
  assign n41152 = n41291 & n41292;
  assign n39948 = ~n41296;
  assign n41293 = ~n41303;
  assign n41275 = n41309 ^ n38800;
  assign n41310 = ~n41309;
  assign n41124 = n41077 & n389;
  assign n41123 = ~n41077;
  assign n41143 = n37379 & n40065;
  assign n41144 = n41097 & n41159;
  assign n41158 = n41165 & n41126;
  assign n41125 = n41165 & n41128;
  assign n41142 = ~n41097;
  assign n37394 = ~n37379;
  assign n41140 = n41180 & n41181;
  assign n41186 = n41100 & n38500;
  assign n41184 = ~n41206;
  assign n41187 = ~n41100;
  assign n41146 = n41221 & n41222;
  assign n41223 = n41259 & n41260;
  assign n41225 = ~n41261;
  assign n41239 = n41262 & n255;
  assign n41268 = n41152 & n41269;
  assign n41267 = ~n41152;
  assign n37617 = n41274 ^ n41275;
  assign n41263 = n41293 & n41294;
  assign n41297 = n41310 & n41311;
  assign n41117 = n41123 & n16551;
  assign n41048 = ~n41124;
  assign n39080 = n41125 ^ n41126;
  assign n41098 = n41140 ^ n41141;
  assign n41129 = n41142 & n41141;
  assign n41118 = ~n41143;
  assign n41121 = ~n41144;
  assign n41127 = ~n41158;
  assign n41120 = ~n41140;
  assign n41145 = n41184 & n41185;
  assign n41096 = ~n41186;
  assign n41166 = n41187 & n38493;
  assign n41149 = ~n41146;
  assign n41188 = n255 ^ n41223;
  assign n41224 = ~n41223;
  assign n41191 = ~n41239;
  assign n41227 = n41263 ^ n41264;
  assign n41241 = n41267 & n41195;
  assign n41197 = ~n41268;
  assign n41243 = n37617 & n39827;
  assign n37657 = ~n37617;
  assign n41266 = ~n41263;
  assign n41276 = ~n41297;
  assign n41003 = n41097 ^ n41098;
  assign n41083 = ~n41117;
  assign n39106 = ~n39080;
  assign n41000 = n41118 & n41119;
  assign n41099 = n41120 & n41121;
  assign n41122 = n41127 & n41128;
  assign n41079 = ~n41129;
  assign n41101 = n41145 ^ n38493;
  assign n41138 = ~n41145;
  assign n41139 = ~n41166;
  assign n41147 = n41188 ^ n41189;
  assign n41207 = n41224 & n41225;
  assign n41151 = n41226 ^ n41227;
  assign n41157 = ~n41241;
  assign n41230 = n37657 & n39600;
  assign n41231 = n37657 & n41242;
  assign n39874 = ~n41243;
  assign n41232 = n37657 & n38800;
  assign n41240 = n41265 & n41266;
  assign n41244 = n41276 & n41277;
  assign n41054 = n41003 & n388;
  assign n41053 = ~n41003;
  assign n41081 = n41000 & n41084;
  assign n41080 = ~n41000;
  assign n41078 = ~n41099;
  assign n37354 = n41100 ^ n41101;
  assign n41076 = ~n41122;
  assign n41130 = n41138 & n41139;
  assign n41020 = n41146 ^ n41147;
  assign n41148 = ~n41147;
  assign n41192 = n41151 & n18839;
  assign n41190 = ~n41207;
  assign n41193 = ~n41151;
  assign n41208 = ~n41230;
  assign n39830 = ~n41231;
  assign n39753 = ~n41232;
  assign n41228 = ~n41240;
  assign n41211 = n41244 ^ n38792;
  assign n41245 = ~n41244;
  assign n41046 = n41053 & n16413;
  assign n40974 = ~n41054;
  assign n41038 = n41076 ^ n41077;
  assign n41040 = n41078 & n41079;
  assign n41055 = n41080 & n41041;
  assign n41045 = ~n41081;
  assign n41056 = n37354 & n40034;
  assign n41075 = n41083 & n41076;
  assign n37323 = ~n37354;
  assign n41102 = n41020 & n38465;
  assign n41095 = ~n41130;
  assign n41103 = ~n41020;
  assign n41060 = n41148 & n41149;
  assign n41150 = n41190 & n41191;
  assign n41137 = ~n41192;
  assign n41167 = n41193 & n254;
  assign n41067 = n41208 & n41209;
  assign n37567 = n41210 ^ n41211;
  assign n41194 = n41228 & n41229;
  assign n41233 = n41245 & n41246;
  assign n40998 = n389 ^ n41038;
  assign n41001 = n41040 ^ n41041;
  assign n41010 = ~n41046;
  assign n41044 = ~n41040;
  assign n41005 = ~n41055;
  assign n41042 = ~n41056;
  assign n41047 = ~n41075;
  assign n41057 = n41095 & n41096;
  assign n41059 = ~n41102;
  assign n41085 = n41103 & n38435;
  assign n41104 = n41150 ^ n41151;
  assign n41136 = ~n41150;
  assign n41106 = ~n41167;
  assign n41153 = n41194 ^ n41195;
  assign n41170 = n41067 & n41198;
  assign n41171 = n37567 & n39530;
  assign n41172 = n37567 & n38763;
  assign n41174 = n37567 & n39754;
  assign n41169 = ~n41067;
  assign n37605 = ~n37567;
  assign n41196 = ~n41194;
  assign n41212 = ~n41233;
  assign n39052 = n40998 ^ n39080;
  assign n40935 = n41000 ^ n41001;
  assign n40920 = n40998 & n39080;
  assign n40926 = n41042 & n41043;
  assign n41018 = n41044 & n41045;
  assign n41039 = n41047 & n41048;
  assign n41019 = n41057 ^ n38465;
  assign n41058 = ~n41057;
  assign n41022 = ~n41085;
  assign n41061 = n254 ^ n41104;
  assign n41131 = n41136 & n41137;
  assign n41064 = n41152 ^ n41153;
  assign n41160 = n41169 & n41110;
  assign n41112 = ~n41170;
  assign n41154 = ~n41171;
  assign n39677 = ~n41172;
  assign n41161 = n37605 & n41173;
  assign n39757 = ~n41174;
  assign n41168 = n41196 & n41197;
  assign n41175 = n41212 & n41213;
  assign n40965 = n40935 & n387;
  assign n40172 = ~n39052;
  assign n40964 = ~n40935;
  assign n40923 = ~n40920;
  assign n41007 = n40926 & n41011;
  assign n41006 = ~n40926;
  assign n41004 = ~n41018;
  assign n37285 = n41019 ^ n41020;
  assign n41002 = ~n41039;
  assign n41049 = n41058 & n41059;
  assign n40944 = n41060 ^ n41061;
  assign n41062 = ~n41061;
  assign n41108 = n41064 & n253;
  assign n41105 = ~n41131;
  assign n41107 = ~n41064;
  assign n40988 = n41154 & n41155;
  assign n41072 = ~n41160;
  assign n39797 = ~n41161;
  assign n41156 = ~n41168;
  assign n41133 = n41175 ^ n38731;
  assign n41176 = ~n41175;
  assign n40940 = n40964 & n16311;
  assign n40888 = ~n40965;
  assign n40963 = n41002 ^ n41003;
  assign n40966 = n41004 & n41005;
  assign n40978 = n41006 & n40967;
  assign n40969 = ~n41007;
  assign n40999 = n41010 & n41002;
  assign n37309 = ~n37285;
  assign n41021 = ~n41049;
  assign n40982 = n41062 & n41060;
  assign n41063 = n41105 & n41106;
  assign n41086 = n41107 & n18788;
  assign n41025 = ~n41108;
  assign n41115 = n40988 & n41029;
  assign n41113 = ~n40988;
  assign n37507 = n41132 ^ n41133;
  assign n41109 = n41156 & n41157;
  assign n41162 = n41176 & n41177;
  assign n40924 = ~n40940;
  assign n40921 = n388 ^ n40963;
  assign n40927 = n40966 ^ n40967;
  assign n40968 = ~n40966;
  assign n40929 = ~n40978;
  assign n40975 = n37309 & n39930;
  assign n40973 = ~n40999;
  assign n40979 = n41021 & n41022;
  assign n41023 = n41063 ^ n41064;
  assign n41065 = ~n41063;
  assign n41066 = ~n41086;
  assign n41068 = n41109 ^ n41110;
  assign n41088 = n41113 & n41114;
  assign n41089 = n37507 & n39576;
  assign n41031 = ~n41115;
  assign n41090 = n37507 & n38731;
  assign n41092 = n37507 & n39679;
  assign n37553 = ~n37507;
  assign n41111 = ~n41109;
  assign n41134 = ~n41162;
  assign n39016 = n40920 ^ n40921;
  assign n40852 = n40926 ^ n40927;
  assign n40922 = ~n40921;
  assign n40943 = n40968 & n40969;
  assign n40934 = n40973 & n40974;
  assign n40941 = ~n40975;
  assign n40945 = n40979 ^ n38412;
  assign n40981 = n40979 & n38412;
  assign n40980 = ~n40979;
  assign n40983 = n253 ^ n41023;
  assign n41050 = n41065 & n41066;
  assign n40985 = n41067 ^ n41068;
  assign n40991 = ~n41088;
  assign n41069 = ~n41089;
  assign n39615 = ~n41090;
  assign n41082 = n37553 & n41091;
  assign n39681 = ~n41092;
  assign n41087 = n41111 & n41112;
  assign n41093 = n41134 & n41135;
  assign n40890 = n40852 & n386;
  assign n40114 = ~n39016;
  assign n40889 = ~n40852;
  assign n40866 = n40922 & n40923;
  assign n40900 = n40934 ^ n40935;
  assign n40855 = n40941 & n40942;
  assign n40928 = ~n40943;
  assign n37247 = n40944 ^ n40945;
  assign n40925 = ~n40934;
  assign n40976 = n40980 & n38439;
  assign n40970 = ~n40981;
  assign n40862 = n40982 ^ n40983;
  assign n40908 = n40983 & n40982;
  assign n41027 = n40985 & n252;
  assign n41024 = ~n41050;
  assign n41026 = ~n40985;
  assign n40916 = n41069 & n41070;
  assign n39719 = ~n41082;
  assign n41071 = ~n41087;
  assign n41052 = n41093 ^ n38724;
  assign n41094 = n41093 & n41116;
  assign n40873 = n40889 & n16246;
  assign n40827 = ~n40890;
  assign n40867 = n387 ^ n40900;
  assign n40869 = ~n40866;
  assign n40903 = n40924 & n40925;
  assign n40891 = n40928 & n40929;
  assign n40906 = n37247 & n39892;
  assign n40907 = n40855 & n40892;
  assign n40904 = ~n40855;
  assign n37270 = ~n37247;
  assign n40946 = n40970 & n40944;
  assign n40948 = n40862 & n38403;
  assign n40931 = ~n40976;
  assign n40947 = ~n40862;
  assign n40911 = ~n40908;
  assign n40984 = n41024 & n41025;
  assign n41012 = n41026 & n18712;
  assign n40951 = ~n41027;
  assign n41034 = n40916 & n40957;
  assign n41032 = ~n40916;
  assign n37446 = n41051 ^ n41052;
  assign n41028 = n41071 & n41072;
  assign n41073 = ~n41094;
  assign n40047 = n40866 ^ n40867;
  assign n40853 = ~n40873;
  assign n40868 = ~n40867;
  assign n40856 = n40891 ^ n40892;
  assign n40887 = ~n40903;
  assign n40893 = ~n40891;
  assign n40901 = n40904 & n40905;
  assign n40898 = ~n40906;
  assign n40894 = ~n40907;
  assign n40930 = ~n40946;
  assign n40936 = n40947 & n38381;
  assign n40897 = ~n40948;
  assign n40949 = n40984 ^ n40985;
  assign n40986 = ~n40984;
  assign n40987 = ~n41012;
  assign n40989 = n41028 ^ n41029;
  assign n41014 = n41032 & n41033;
  assign n40959 = ~n41034;
  assign n41015 = n37446 & n39399;
  assign n41016 = n37446 & n38701;
  assign n41017 = n37446 & n41035;
  assign n37491 = ~n37446;
  assign n41030 = ~n41028;
  assign n41036 = n41073 & n41074;
  assign n40024 = ~n40047;
  assign n40799 = n40855 ^ n40856;
  assign n40795 = n40868 & n40869;
  assign n40851 = n40887 & n40888;
  assign n40874 = n40893 & n40894;
  assign n40802 = n40898 & n40899;
  assign n40858 = ~n40901;
  assign n40895 = n40930 & n40931;
  assign n40865 = ~n40936;
  assign n40909 = n252 ^ n40949;
  assign n40977 = n40986 & n40987;
  assign n40913 = n40988 ^ n40989;
  assign n40919 = ~n41014;
  assign n40992 = ~n41015;
  assign n41009 = n37491 & n39603;
  assign n39538 = ~n41016;
  assign n39606 = ~n41017;
  assign n41013 = n41030 & n41031;
  assign n40995 = n41036 ^ n41037;
  assign n40829 = n40799 & n16138;
  assign n40825 = ~n40799;
  assign n40828 = n40851 ^ n40852;
  assign n40861 = n40802 & n40831;
  assign n40854 = ~n40851;
  assign n40859 = ~n40802;
  assign n40857 = ~n40874;
  assign n40863 = n40895 ^ n38381;
  assign n40896 = ~n40895;
  assign n40806 = n40908 ^ n40909;
  assign n40910 = ~n40909;
  assign n40952 = n40913 & n18693;
  assign n40950 = ~n40977;
  assign n40953 = ~n40913;
  assign n40847 = n40992 & n40993;
  assign n40954 = n40994 ^ n40995;
  assign n40996 = n40995 & n41008;
  assign n39644 = ~n41009;
  assign n40997 = n40995 & n38713;
  assign n40990 = ~n41013;
  assign n38734 = ~n40995;
  assign n40814 = n40825 & n385;
  assign n40796 = n386 ^ n40828;
  assign n40800 = ~n40829;
  assign n40839 = n40853 & n40854;
  assign n40830 = n40857 & n40858;
  assign n40840 = n40859 & n40860;
  assign n40833 = ~n40861;
  assign n37213 = n40862 ^ n40863;
  assign n40875 = n40896 & n40897;
  assign n40876 = n40806 & n38371;
  assign n40877 = ~n40806;
  assign n40841 = n40910 & n40911;
  assign n40912 = n40950 & n40951;
  assign n40915 = ~n40952;
  assign n40937 = n40953 & n251;
  assign n39564 = n40954 ^ n40955;
  assign n40962 = n40847 & n40884;
  assign n40960 = ~n40847;
  assign n40956 = n40990 & n40991;
  assign n40971 = ~n40996;
  assign n39507 = ~n40997;
  assign n38966 = n40795 ^ n40796;
  assign n40797 = ~n40796;
  assign n40770 = ~n40814;
  assign n40803 = n40830 ^ n40831;
  assign n40834 = n37213 & n39788;
  assign n40826 = ~n40839;
  assign n40832 = ~n40830;
  assign n40805 = ~n40840;
  assign n37236 = ~n37213;
  assign n40864 = ~n40875;
  assign n40809 = ~n40876;
  assign n40870 = n40877 & n38346;
  assign n40878 = n40912 ^ n40913;
  assign n40914 = ~n40912;
  assign n40880 = ~n40937;
  assign n40917 = n40956 ^ n40957;
  assign n40939 = n40960 & n40961;
  assign n40886 = ~n40962;
  assign n40932 = n40971 & n40972;
  assign n40958 = ~n40956;
  assign n39970 = ~n38966;
  assign n40744 = n40797 & n40795;
  assign n40747 = n40802 ^ n40803;
  assign n40798 = n40826 & n40827;
  assign n40815 = n40832 & n40833;
  assign n40810 = ~n40834;
  assign n40835 = n40864 & n40865;
  assign n40837 = ~n40870;
  assign n40842 = n251 ^ n40878;
  assign n40902 = n40914 & n40915;
  assign n40844 = n40916 ^ n40917;
  assign n40794 = n40932 ^ n40933;
  assign n40850 = ~n40939;
  assign n40938 = n40958 & n40959;
  assign n40771 = n40747 & n16072;
  assign n40772 = ~n40747;
  assign n40768 = n40798 ^ n40799;
  assign n40734 = n40810 & n40811;
  assign n40801 = ~n40798;
  assign n40804 = ~n40815;
  assign n40807 = n40835 ^ n38346;
  assign n40836 = ~n40835;
  assign n40750 = n40841 ^ n40842;
  assign n40785 = n40842 & n40841;
  assign n40881 = n40844 & n18624;
  assign n40879 = ~n40902;
  assign n40882 = ~n40844;
  assign n40918 = ~n40938;
  assign n40745 = n385 ^ n40768;
  assign n40748 = ~n40771;
  assign n40758 = n40772 & n384;
  assign n40781 = n40734 & n40761;
  assign n40783 = n40800 & n40801;
  assign n40784 = n40804 & n40805;
  assign n40779 = ~n40734;
  assign n37203 = n40806 ^ n40807;
  assign n40816 = n40836 & n40837;
  assign n40817 = n40750 & n38344;
  assign n40818 = ~n40750;
  assign n40788 = ~n40785;
  assign n40843 = n40879 & n40880;
  assign n40846 = ~n40881;
  assign n40871 = n40882 & n250;
  assign n40883 = n40918 & n40919;
  assign n38931 = n40744 ^ n40745;
  assign n40697 = n40745 & n40744;
  assign n40725 = ~n40758;
  assign n40773 = n40779 & n40780;
  assign n40774 = n37203 & n39682;
  assign n40759 = ~n40781;
  assign n40769 = ~n40783;
  assign n40760 = ~n40784;
  assign n37177 = ~n37203;
  assign n40808 = ~n40816;
  assign n40753 = ~n40817;
  assign n40812 = n40818 & n38309;
  assign n40819 = n40843 ^ n40844;
  assign n40845 = ~n40843;
  assign n40821 = ~n40871;
  assign n40848 = n40883 ^ n40884;
  assign n40885 = ~n40883;
  assign n39871 = ~n38931;
  assign n40700 = ~n40697;
  assign n40754 = n40759 & n40760;
  assign n40735 = n40760 ^ n40761;
  assign n40746 = n40769 & n40770;
  assign n40737 = ~n40773;
  assign n40755 = ~n40774;
  assign n40775 = n40808 & n40809;
  assign n40777 = ~n40812;
  assign n40786 = n250 ^ n40819;
  assign n40838 = n40845 & n40846;
  assign n40790 = n40847 ^ n40848;
  assign n40872 = n40885 & n40886;
  assign n40702 = n40734 ^ n40735;
  assign n40723 = n40746 ^ n40747;
  assign n40736 = ~n40754;
  assign n40689 = n40755 & n40756;
  assign n40749 = ~n40746;
  assign n40751 = n40775 ^ n38309;
  assign n40776 = ~n40775;
  assign n40778 = n40785 ^ n40786;
  assign n40787 = ~n40786;
  assign n40822 = n40790 & n18560;
  assign n40820 = ~n40838;
  assign n40823 = ~n40790;
  assign n40849 = ~n40872;
  assign n40698 = n384 ^ n40723;
  assign n40713 = n40702 & n399;
  assign n40712 = ~n40702;
  assign n40714 = n40736 & n40737;
  assign n40731 = n40689 & n40738;
  assign n40733 = n40748 & n40749;
  assign n40730 = ~n40689;
  assign n37143 = n40750 ^ n40751;
  assign n40762 = n40776 & n40777;
  assign n40764 = n40778 & n38299;
  assign n40763 = ~n40778;
  assign n40739 = n40787 & n40788;
  assign n40789 = n40820 & n40821;
  assign n40792 = ~n40822;
  assign n40813 = n40823 & n249;
  assign n40824 = n40849 & n40850;
  assign n38878 = n40697 ^ n40698;
  assign n40699 = ~n40698;
  assign n40705 = n40712 & n15958;
  assign n40670 = ~n40713;
  assign n40690 = n40714 ^ n40715;
  assign n40717 = ~n40714;
  assign n40726 = n40730 & n40715;
  assign n40727 = n37143 & n39630;
  assign n40716 = ~n40731;
  assign n40724 = ~n40733;
  assign n37168 = ~n37143;
  assign n40752 = ~n40762;
  assign n40757 = n40763 & n38270;
  assign n40729 = ~n40764;
  assign n40765 = n40789 ^ n40790;
  assign n40791 = ~n40789;
  assign n40767 = ~n40813;
  assign n40793 = n248 ^ n40824;
  assign n39794 = ~n38878;
  assign n40646 = n40689 ^ n40690;
  assign n40655 = n40699 & n40700;
  assign n40692 = ~n40705;
  assign n40708 = n40716 & n40717;
  assign n40701 = n40724 & n40725;
  assign n40694 = ~n40726;
  assign n40706 = ~n40727;
  assign n40709 = n40752 & n40753;
  assign n40704 = ~n40757;
  assign n40740 = n249 ^ n40765;
  assign n40782 = n40791 & n40792;
  assign n40743 = n40793 ^ n40794;
  assign n40668 = n40646 & n398;
  assign n40667 = ~n40646;
  assign n40658 = ~n40655;
  assign n40678 = n40701 ^ n40702;
  assign n40649 = n40706 & n40707;
  assign n40693 = ~n40708;
  assign n40691 = ~n40701;
  assign n40728 = ~n40709;
  assign n40732 = n40729 & n40704;
  assign n40659 = n40739 ^ n40740;
  assign n40741 = ~n40740;
  assign n40766 = ~n40782;
  assign n40664 = n40667 & n15897;
  assign n40633 = ~n40668;
  assign n40656 = n399 ^ n40678;
  assign n40683 = n40691 & n40692;
  assign n40671 = n40693 & n40694;
  assign n40686 = n40649 & n40672;
  assign n40684 = ~n40649;
  assign n40718 = n40728 & n40729;
  assign n40720 = n40659 & n38261;
  assign n40710 = ~n40732;
  assign n40719 = ~n40659;
  assign n40721 = n40741 & n40739;
  assign n40742 = n40766 & n40767;
  assign n38848 = n40655 ^ n40656;
  assign n40648 = ~n40664;
  assign n40657 = ~n40656;
  assign n40650 = n40671 ^ n40672;
  assign n40669 = ~n40683;
  assign n40674 = ~n40671;
  assign n40679 = n40684 & n40685;
  assign n40673 = ~n40686;
  assign n37110 = n40709 ^ n40710;
  assign n40703 = ~n40718;
  assign n40711 = n40719 & n38230;
  assign n40663 = ~n40720;
  assign n40722 = n40742 ^ n40743;
  assign n39735 = ~n38848;
  assign n40615 = n40649 ^ n40650;
  assign n40610 = n40657 & n40658;
  assign n40665 = n40669 & n40670;
  assign n40666 = n40673 & n40674;
  assign n40652 = ~n40679;
  assign n40687 = n37110 & n39518;
  assign n40680 = n40703 & n40704;
  assign n37113 = ~n37110;
  assign n40682 = ~n40711;
  assign n40622 = n40721 ^ n40722;
  assign n40634 = n40615 & n15813;
  assign n40631 = ~n40615;
  assign n40645 = ~n40665;
  assign n40651 = ~n40666;
  assign n40660 = n40680 ^ n38230;
  assign n40675 = ~n40687;
  assign n40681 = ~n40680;
  assign n40695 = n40622 & n38192;
  assign n40696 = ~n40622;
  assign n40627 = n40631 & n397;
  assign n40616 = ~n40634;
  assign n40626 = n40645 ^ n40646;
  assign n40644 = n40648 & n40645;
  assign n40635 = n40651 & n40652;
  assign n37053 = n40659 ^ n40660;
  assign n40618 = n40675 & n40676;
  assign n40677 = n40681 & n40682;
  assign n40643 = ~n40695;
  assign n40688 = n40696 & n38228;
  assign n40611 = n398 ^ n40626;
  assign n40598 = ~n40627;
  assign n40619 = n40635 ^ n40636;
  assign n40632 = ~n40644;
  assign n40637 = ~n40635;
  assign n40640 = n37053 & n39435;
  assign n37083 = ~n37053;
  assign n40654 = n40618 & n40661;
  assign n40653 = ~n40618;
  assign n40662 = ~n40677;
  assign n40625 = ~n40688;
  assign n38811 = n40610 ^ n40611;
  assign n40576 = n40611 & n40610;
  assign n40581 = n40618 ^ n40619;
  assign n40614 = n40632 & n40633;
  assign n40629 = ~n40640;
  assign n40647 = n40653 & n40636;
  assign n40638 = ~n40654;
  assign n40641 = n40662 & n40663;
  assign n39641 = ~n38811;
  assign n40600 = n40581 & n396;
  assign n40579 = ~n40576;
  assign n40599 = ~n40581;
  assign n40596 = n40614 ^ n40615;
  assign n40617 = ~n40614;
  assign n40584 = n40629 & n40630;
  assign n40628 = n40637 & n40638;
  assign n40623 = n40641 ^ n38192;
  assign n40621 = ~n40647;
  assign n40642 = ~n40641;
  assign n40577 = n397 ^ n40596;
  assign n40593 = n40599 & n15732;
  assign n40562 = ~n40600;
  assign n40612 = n40616 & n40617;
  assign n40588 = ~n40584;
  assign n37029 = n40622 ^ n40623;
  assign n40620 = ~n40628;
  assign n40639 = n40642 & n40643;
  assign n38775 = n40576 ^ n40577;
  assign n40578 = ~n40577;
  assign n40583 = ~n40593;
  assign n40597 = ~n40612;
  assign n40601 = n40620 & n40621;
  assign n37050 = ~n37029;
  assign n40624 = ~n40639;
  assign n39578 = ~n38775;
  assign n39533 = n40578 & n40579;
  assign n40580 = n40597 & n40598;
  assign n40585 = n40601 ^ n40602;
  assign n40604 = n40601 & n40607;
  assign n40605 = n37050 & n39405;
  assign n40603 = ~n40601;
  assign n40613 = n40624 & n40625;
  assign n40560 = n40580 ^ n40581;
  assign n40546 = n40584 ^ n40585;
  assign n40582 = ~n40580;
  assign n40594 = n40603 & n40602;
  assign n40587 = ~n40604;
  assign n40589 = ~n40605;
  assign n40609 = n40613 & n38153;
  assign n40608 = ~n40613;
  assign n39489 = n396 ^ n40560;
  assign n40564 = n40546 & n395;
  assign n40563 = ~n40546;
  assign n40572 = n40582 & n40583;
  assign n40586 = n40587 & n40588;
  assign n40534 = n40589 & n40590;
  assign n40567 = ~n40594;
  assign n40606 = n40608 & n38190;
  assign n40592 = ~n40609;
  assign n40511 = n39489 & n39533;
  assign n40556 = n40563 & n15662;
  assign n40533 = ~n40564;
  assign n40561 = ~n40572;
  assign n40569 = n40534 & n40573;
  assign n40566 = ~n40586;
  assign n40568 = ~n40534;
  assign n40591 = n40592 & n40595;
  assign n40575 = ~n40606;
  assign n40514 = ~n40511;
  assign n40550 = ~n40556;
  assign n40545 = n40561 & n40562;
  assign n40551 = n40566 & n40567;
  assign n40565 = n40568 & n40552;
  assign n40554 = ~n40569;
  assign n40574 = ~n40591;
  assign n40570 = n40575 & n40592;
  assign n40531 = n40545 ^ n40546;
  assign n40535 = n40551 ^ n40552;
  assign n40549 = ~n40545;
  assign n40553 = ~n40551;
  assign n40537 = ~n40565;
  assign n37000 = n40570 ^ n40571;
  assign n40557 = n40574 & n40575;
  assign n40512 = n395 ^ n40531;
  assign n40503 = n40534 ^ n40535;
  assign n40540 = n40549 & n40550;
  assign n40547 = n40553 & n40554;
  assign n40541 = n40557 ^ n38151;
  assign n37061 = ~n37000;
  assign n40558 = ~n40557;
  assign n37747 = n40511 ^ n40512;
  assign n40513 = ~n40512;
  assign n40518 = n40503 & n394;
  assign n40517 = ~n40503;
  assign n40532 = ~n40540;
  assign n36960 = n40541 ^ n40542;
  assign n40536 = ~n40547;
  assign n40548 = n37061 & n39343;
  assign n40555 = n40558 & n40559;
  assign n40473 = n40496 ^ n37747;
  assign n40477 = n38663 ^ n37747;
  assign n36790 = n37741 ^ n37747;
  assign n40394 = n37747 & n37741;
  assign n40464 = n40513 & n40514;
  assign n40515 = n40517 & n15572;
  assign n40480 = ~n40518;
  assign n40526 = n40532 & n40533;
  assign n40519 = n40536 & n40537;
  assign n36991 = ~n36960;
  assign n40538 = ~n40548;
  assign n40543 = ~n40555;
  assign n38582 = n167 ^ n40473;
  assign n40322 = n40477 & n40478;
  assign n40194 = n40473 & n167;
  assign n40498 = ~n40515;
  assign n40501 = n40519 ^ n40520;
  assign n40499 = ~n40526;
  assign n40521 = n36991 & n39336;
  assign n40506 = ~n40519;
  assign n40500 = n40538 & n40539;
  assign n40527 = n40543 & n40544;
  assign n40458 = n40322 & n40290;
  assign n40199 = ~n38582;
  assign n40456 = ~n40322;
  assign n40497 = n40498 & n40499;
  assign n40460 = n40500 ^ n40501;
  assign n40485 = n40499 ^ n40503;
  assign n40504 = ~n40521;
  assign n40524 = n40500 & n40520;
  assign n40508 = n40527 ^ n40528;
  assign n40522 = ~n40500;
  assign n40529 = ~n40527;
  assign n40451 = n40456 & n40457;
  assign n40305 = ~n40458;
  assign n40465 = n394 ^ n40485;
  assign n40481 = n40460 & n15529;
  assign n40479 = ~n40497;
  assign n40482 = ~n40460;
  assign n40441 = n40504 & n40505;
  assign n36904 = n40508 ^ n38110;
  assign n40516 = n40522 & n40523;
  assign n40507 = ~n40524;
  assign n40525 = n40529 & n40530;
  assign n40337 = ~n40451;
  assign n40452 = n40464 ^ n40465;
  assign n40412 = n40465 & n40464;
  assign n40459 = n40479 & n40480;
  assign n40462 = ~n40481;
  assign n40474 = n40482 & n393;
  assign n40490 = n40441 & n40467;
  assign n40491 = n36904 & n39241;
  assign n40488 = ~n40441;
  assign n36978 = ~n36904;
  assign n40502 = n40506 & n40507;
  assign n40487 = ~n40516;
  assign n40509 = ~n40525;
  assign n40439 = n40452 & n37542;
  assign n40440 = ~n40452;
  assign n40435 = n40459 ^ n40460;
  assign n40415 = ~n40412;
  assign n40461 = ~n40459;
  assign n40437 = ~n40474;
  assign n40483 = n40488 & n40489;
  assign n40468 = ~n40490;
  assign n40475 = ~n40491;
  assign n40486 = ~n40502;
  assign n40492 = n40509 & n40510;
  assign n40413 = n393 ^ n40435;
  assign n40396 = ~n40439;
  assign n40434 = n40440 & n37714;
  assign n40450 = n40461 & n40462;
  assign n40425 = n40475 & n40476;
  assign n40444 = ~n40483;
  assign n40466 = n40486 & n40487;
  assign n40470 = n40492 ^ n40493;
  assign n40494 = ~n40492;
  assign n40346 = n40412 ^ n40413;
  assign n40414 = ~n40413;
  assign n40421 = ~n40434;
  assign n40436 = ~n40450;
  assign n40455 = n40425 & n40399;
  assign n40442 = n40466 ^ n40467;
  assign n40453 = ~n40425;
  assign n36865 = n40470 ^ n38015;
  assign n40469 = ~n40466;
  assign n40484 = n40494 & n40495;
  assign n40388 = n40346 & n37530;
  assign n40389 = ~n40346;
  assign n40365 = n40414 & n40415;
  assign n40416 = n40421 & n40394;
  assign n40393 = n40421 & n40396;
  assign n40417 = n40436 & n40437;
  assign n40418 = n40441 ^ n40442;
  assign n40445 = n40453 & n40454;
  assign n40446 = n36865 & n39227;
  assign n40426 = ~n40455;
  assign n36963 = ~n36865;
  assign n40463 = n40468 & n40469;
  assign n40471 = ~n40484;
  assign n40371 = ~n40388;
  assign n40383 = n40389 & n37532;
  assign n36621 = n40393 ^ n40394;
  assign n40372 = ~n40365;
  assign n40395 = ~n40416;
  assign n40391 = n40417 ^ n40418;
  assign n40407 = ~n40417;
  assign n40422 = n40418 & n15486;
  assign n40423 = ~n40418;
  assign n40401 = ~n40445;
  assign n40432 = ~n40446;
  assign n40443 = ~n40463;
  assign n40447 = n40471 & n40472;
  assign n38631 = n37542 ^ n36621;
  assign n40352 = ~n40383;
  assign n36764 = ~n36621;
  assign n40366 = n392 ^ n40391;
  assign n40390 = n40395 & n40396;
  assign n40408 = ~n40422;
  assign n40419 = n40423 & n392;
  assign n40354 = n40432 & n40433;
  assign n40424 = n40443 & n40444;
  assign n40429 = n40447 ^ n37978;
  assign n40448 = ~n40447;
  assign n40323 = n38631 ^ n38626;
  assign n40326 = n40365 ^ n40366;
  assign n40306 = n40366 & n40372;
  assign n40368 = ~n40390;
  assign n40397 = n40407 & n40408;
  assign n40385 = ~n40419;
  assign n40411 = n40354 & n40376;
  assign n40398 = n40424 ^ n40425;
  assign n40409 = ~n40354;
  assign n36831 = n40428 ^ n40429;
  assign n40427 = ~n40424;
  assign n40438 = n40448 & n40449;
  assign n40289 = n40322 ^ n40323;
  assign n40324 = n40323 & n40337;
  assign n40348 = n40326 & n37437;
  assign n40349 = ~n40326;
  assign n40347 = n40368 ^ n37532;
  assign n40367 = n40371 & n40368;
  assign n40384 = ~n40397;
  assign n40340 = n40398 ^ n40399;
  assign n40402 = n40409 & n40410;
  assign n40403 = n36831 & n39192;
  assign n40378 = ~n40411;
  assign n36877 = ~n36831;
  assign n40420 = n40426 & n40427;
  assign n40430 = ~n40438;
  assign n40276 = n40289 ^ n40290;
  assign n40304 = ~n40324;
  assign n36588 = n40346 ^ n40347;
  assign n40321 = ~n40348;
  assign n40338 = n40349 & n37455;
  assign n40351 = ~n40367;
  assign n40362 = n40384 & n40385;
  assign n40373 = n40340 & n15473;
  assign n40374 = ~n40340;
  assign n40357 = ~n40402;
  assign n40386 = ~n40403;
  assign n40400 = ~n40420;
  assign n40404 = n40430 & n40431;
  assign n40263 = n40276 & n166;
  assign n40262 = ~n40276;
  assign n40277 = n40304 & n40305;
  assign n38618 = n36588 ^ n37532;
  assign n36590 = ~n36588;
  assign n40292 = ~n40338;
  assign n40325 = n40351 & n40352;
  assign n40339 = n407 ^ n40362;
  assign n40364 = ~n40362;
  assign n40363 = ~n40373;
  assign n40369 = n40374 & n407;
  assign n40294 = n40386 & n40387;
  assign n40375 = n40400 & n40401;
  assign n40380 = n40404 ^ n37959;
  assign n40405 = ~n40404;
  assign n40255 = n40262 & n17578;
  assign n40196 = ~n40263;
  assign n40238 = n40277 ^ n40264;
  assign n40239 = n38618 ^ n38611;
  assign n40223 = ~n40277;
  assign n38594 = n40325 ^ n40326;
  assign n40307 = n40339 ^ n40340;
  assign n40320 = ~n40325;
  assign n40353 = n40363 & n40364;
  assign n40342 = ~n40369;
  assign n40355 = n40375 ^ n40376;
  assign n40313 = ~n40294;
  assign n36892 = n40379 ^ n40380;
  assign n40377 = ~n40375;
  assign n40392 = n40405 & n40406;
  assign n40160 = n40238 ^ n40239;
  assign n40227 = ~n40255;
  assign n40256 = n40239 & n40264;
  assign n40257 = ~n40239;
  assign n40116 = n38594 ^ n38563;
  assign n36491 = n38594 ^ n37437;
  assign n40229 = n40306 ^ n40307;
  assign n40243 = n40307 & n40306;
  assign n40317 = n40320 & n40321;
  assign n40341 = ~n40353;
  assign n40309 = n40354 ^ n40355;
  assign n40358 = n36892 & n39105;
  assign n36814 = ~n36892;
  assign n40370 = n40377 & n40378;
  assign n40381 = ~n40392;
  assign n40209 = n40160 & n17487;
  assign n40221 = n40227 & n40194;
  assign n40193 = n40227 & n40196;
  assign n40210 = ~n40160;
  assign n40191 = ~n40256;
  assign n40240 = n40257 & n40258;
  assign n40265 = n40116 & n40151;
  assign n40266 = ~n40116;
  assign n36526 = ~n36491;
  assign n40279 = n40229 & n37379;
  assign n40278 = ~n40229;
  assign n40246 = ~n40243;
  assign n40291 = ~n40317;
  assign n40308 = n40341 & n40342;
  assign n40327 = n40309 & n15399;
  assign n40328 = ~n40309;
  assign n40343 = ~n40358;
  assign n40356 = ~n40370;
  assign n40359 = n40381 & n40382;
  assign n38525 = n40193 ^ n40194;
  assign n40161 = ~n40209;
  assign n40197 = n40210 & n165;
  assign n40195 = ~n40221;
  assign n40222 = ~n40240;
  assign n40153 = ~n40265;
  assign n40259 = n40266 & n40267;
  assign n40269 = n40278 & n37394;
  assign n40213 = ~n40279;
  assign n40268 = n40291 & n40292;
  assign n40280 = n40308 ^ n40309;
  assign n40310 = ~n40308;
  assign n40311 = ~n40327;
  assign n40318 = n40328 & n406;
  assign n40217 = n40343 & n40344;
  assign n40329 = n40356 & n40357;
  assign n40334 = n40359 ^ n37918;
  assign n40360 = ~n40359;
  assign n38554 = ~n38525;
  assign n40159 = n40195 & n40196;
  assign n40125 = ~n40197;
  assign n40211 = n40222 & n40223;
  assign n40119 = ~n40259;
  assign n40228 = n40268 ^ n37394;
  assign n40242 = ~n40269;
  assign n40244 = n406 ^ n40280;
  assign n40241 = ~n40268;
  assign n40293 = n40310 & n40311;
  assign n40282 = ~n40318;
  assign n40316 = n40217 & n40250;
  assign n40295 = n40329 ^ n40330;
  assign n40314 = ~n40217;
  assign n36812 = n40333 ^ n40334;
  assign n40332 = n40329 & n40345;
  assign n40331 = ~n40329;
  assign n40350 = n40360 & n40361;
  assign n40123 = n40159 ^ n40160;
  assign n40162 = ~n40159;
  assign n40190 = ~n40211;
  assign n36474 = n40228 ^ n40229;
  assign n40230 = n40241 & n40242;
  assign n40136 = n40243 ^ n40244;
  assign n40245 = ~n40244;
  assign n40281 = ~n40293;
  assign n40248 = n40294 ^ n40295;
  assign n40297 = n40314 & n40315;
  assign n40298 = n36812 & n39128;
  assign n40252 = ~n40316;
  assign n40299 = n36812 & n39154;
  assign n36771 = ~n36812;
  assign n40319 = n40331 & n40330;
  assign n40312 = ~n40332;
  assign n40335 = ~n40350;
  assign n40087 = n165 ^ n40123;
  assign n40149 = n40161 & n40162;
  assign n40150 = n40190 & n40191;
  assign n38568 = n36474 ^ n37379;
  assign n40198 = n36474 & n38582;
  assign n36420 = ~n36474;
  assign n40215 = n40136 & n37323;
  assign n40212 = ~n40230;
  assign n40214 = ~n40136;
  assign n40180 = n40245 & n40246;
  assign n40247 = n40281 & n40282;
  assign n40271 = n40248 & n405;
  assign n40270 = ~n40248;
  assign n40220 = ~n40297;
  assign n40285 = ~n40298;
  assign n39139 = ~n40299;
  assign n40287 = n36771 & n40300;
  assign n40296 = n40312 & n40313;
  assign n40284 = ~n40319;
  assign n40301 = n40335 & n40336;
  assign n38502 = n40087 ^ n38525;
  assign n40003 = n40087 & n38525;
  assign n40124 = ~n40149;
  assign n40115 = n40150 ^ n40151;
  assign n40032 = n38568 ^ n38552;
  assign n40152 = ~n40150;
  assign n38584 = ~n40198;
  assign n40192 = n36420 & n40199;
  assign n40177 = n40212 & n40213;
  assign n40200 = n40214 & n37354;
  assign n40178 = ~n40215;
  assign n40183 = ~n40180;
  assign n40216 = n40247 ^ n40248;
  assign n40231 = ~n40247;
  assign n40260 = n40270 & n15354;
  assign n40202 = ~n40271;
  assign n40143 = n40285 & n40286;
  assign n39156 = ~n40287;
  assign n40283 = ~n40296;
  assign n40273 = n40301 ^ n37881;
  assign n40302 = ~n40301;
  assign n40030 = ~n38502;
  assign n40079 = n40115 ^ n40116;
  assign n40078 = n40124 & n40125;
  assign n40126 = n40032 & n40065;
  assign n40127 = ~n40032;
  assign n40135 = n40152 & n40153;
  assign n40137 = n40177 ^ n37354;
  assign n38597 = ~n40192;
  assign n40179 = ~n40177;
  assign n40139 = ~n40200;
  assign n40181 = n405 ^ n40216;
  assign n40232 = ~n40260;
  assign n40254 = n40143 & n40261;
  assign n40253 = ~n40143;
  assign n36723 = n40272 ^ n40273;
  assign n40249 = n40283 & n40284;
  assign n40288 = n40302 & n40303;
  assign n40048 = n40078 ^ n40079;
  assign n40080 = n40079 & n17421;
  assign n40081 = ~n40079;
  assign n40055 = ~n40078;
  assign n40051 = ~n40126;
  assign n40117 = n40127 & n40128;
  assign n40118 = ~n40135;
  assign n36402 = n40136 ^ n40137;
  assign n40163 = n40178 & n40179;
  assign n40066 = n40180 ^ n40181;
  assign n40182 = ~n40181;
  assign n40224 = n40231 & n40232;
  assign n40218 = n40249 ^ n40250;
  assign n40234 = n40253 & n40187;
  assign n40189 = ~n40254;
  assign n36769 = ~n36723;
  assign n40251 = ~n40249;
  assign n40274 = ~n40288;
  assign n40004 = n164 ^ n40048;
  assign n40054 = ~n40080;
  assign n40062 = n40081 & n164;
  assign n38509 = n36402 ^ n37354;
  assign n40082 = ~n40117;
  assign n40102 = n40118 & n40119;
  assign n36346 = ~n36402;
  assign n40140 = n40066 & n37309;
  assign n40138 = ~n40163;
  assign n40141 = ~n40066;
  assign n40089 = n40182 & n40183;
  assign n40165 = n40217 ^ n40218;
  assign n40201 = ~n40224;
  assign n40146 = ~n40234;
  assign n40225 = n36769 & n39032;
  assign n40233 = n40251 & n40252;
  assign n40235 = n40274 & n40275;
  assign n38468 = n40003 ^ n40004;
  assign n39897 = n40004 & n40003;
  assign n40049 = n40054 & n40055;
  assign n40017 = ~n40062;
  assign n39972 = n38509 ^ n38493;
  assign n40064 = ~n40102;
  assign n40103 = n40138 & n40139;
  assign n40069 = ~n40140;
  assign n40129 = n40141 & n37285;
  assign n40092 = ~n40089;
  assign n40184 = n40165 & n15327;
  assign n40164 = n40201 & n40202;
  assign n40185 = ~n40165;
  assign n40203 = ~n40225;
  assign n40219 = ~n40233;
  assign n40206 = n40235 ^ n37843;
  assign n40236 = ~n40235;
  assign n39949 = ~n38468;
  assign n40016 = ~n40049;
  assign n40035 = n39972 & n40006;
  assign n40033 = ~n39972;
  assign n40031 = n40064 ^ n40065;
  assign n40063 = n40082 & n40064;
  assign n40067 = n40103 ^ n37285;
  assign n40104 = ~n40103;
  assign n40105 = ~n40129;
  assign n40130 = n40164 ^ n40165;
  assign n40154 = ~n40184;
  assign n40166 = n40185 & n404;
  assign n40155 = ~n40164;
  assign n40072 = n40203 & n40204;
  assign n36672 = n40205 ^ n40206;
  assign n40186 = n40219 & n40220;
  assign n40226 = n40236 & n40237;
  assign n39978 = n40016 & n40017;
  assign n39979 = n40031 ^ n40032;
  assign n40018 = n40033 & n40034;
  assign n40008 = ~n40035;
  assign n40050 = ~n40063;
  assign n36273 = n40066 ^ n40067;
  assign n40088 = n40104 & n40105;
  assign n40090 = n404 ^ n40130;
  assign n40142 = n40154 & n40155;
  assign n40121 = ~n40166;
  assign n40144 = n40186 ^ n40187;
  assign n40170 = n40072 & n40109;
  assign n40171 = n36672 & n38964;
  assign n40173 = n36672 & n39052;
  assign n40168 = ~n40072;
  assign n36710 = ~n36672;
  assign n40188 = ~n40186;
  assign n40207 = ~n40226;
  assign n39938 = n39978 ^ n39979;
  assign n39952 = ~n39978;
  assign n39987 = n39979 & n163;
  assign n39986 = ~n39979;
  assign n39974 = ~n40018;
  assign n38485 = n37309 ^ n36273;
  assign n40029 = n36273 & n38502;
  assign n40005 = n40050 & n40051;
  assign n36309 = ~n36273;
  assign n40068 = ~n40088;
  assign n39989 = n40089 ^ n40090;
  assign n40091 = ~n40090;
  assign n40120 = ~n40142;
  assign n40084 = n40143 ^ n40144;
  assign n40156 = n40168 & n40169;
  assign n40111 = ~n40170;
  assign n40147 = ~n40171;
  assign n40157 = n36710 & n40172;
  assign n39054 = ~n40173;
  assign n40167 = n40188 & n40189;
  assign n40174 = n40207 & n40208;
  assign n39898 = n163 ^ n39938;
  assign n39980 = n39986 & n17333;
  assign n39910 = ~n39987;
  assign n39891 = n38485 ^ n38435;
  assign n39971 = n40005 ^ n40006;
  assign n38504 = ~n40029;
  assign n40015 = n36309 & n40030;
  assign n40007 = ~n40005;
  assign n40036 = n40068 & n40069;
  assign n40057 = n39989 & n37270;
  assign n40056 = ~n39989;
  assign n40009 = n40091 & n40092;
  assign n40083 = n40120 & n40121;
  assign n40107 = n40084 & n403;
  assign n40106 = ~n40084;
  assign n39997 = n40147 & n40148;
  assign n40075 = ~n40156;
  assign n39071 = ~n40157;
  assign n40145 = ~n40167;
  assign n40132 = n40174 ^ n37841;
  assign n40175 = ~n40174;
  assign n38452 = n39897 ^ n39898;
  assign n39899 = ~n39898;
  assign n39878 = n39971 ^ n39972;
  assign n39953 = n39891 & n39930;
  assign n39951 = ~n39980;
  assign n39954 = ~n39891;
  assign n39988 = n40007 & n40008;
  assign n38521 = ~n40015;
  assign n39990 = n40036 ^ n37247;
  assign n40038 = ~n40036;
  assign n40052 = n40056 & n37247;
  assign n40037 = ~n40057;
  assign n40012 = ~n40009;
  assign n40053 = n40083 ^ n40084;
  assign n40071 = ~n40083;
  assign n40093 = n40106 & n15296;
  assign n40040 = ~n40107;
  assign n40113 = n39997 & n40122;
  assign n40112 = ~n39997;
  assign n36613 = n40131 ^ n40132;
  assign n40108 = n40145 & n40146;
  assign n40158 = n40175 & n40176;
  assign n39864 = ~n38452;
  assign n39812 = n39899 & n39897;
  assign n39927 = n39878 & n17249;
  assign n39928 = ~n39878;
  assign n39939 = n39951 & n39952;
  assign n39880 = ~n39953;
  assign n39940 = n39954 & n39955;
  assign n39973 = ~n39988;
  assign n36254 = n39989 ^ n39990;
  assign n40019 = n40037 & n40038;
  assign n39992 = ~n40052;
  assign n40010 = n403 ^ n40053;
  assign n40070 = ~n40093;
  assign n40073 = n40108 ^ n40109;
  assign n40095 = n40112 & n40044;
  assign n40046 = ~n40113;
  assign n40096 = n36613 & n38975;
  assign n40097 = n36613 & n40114;
  assign n36660 = ~n36613;
  assign n40110 = ~n40108;
  assign n40133 = ~n40158;
  assign n39875 = ~n39927;
  assign n39908 = n39928 & n162;
  assign n39909 = ~n39939;
  assign n39911 = ~n39940;
  assign n38449 = n36254 ^ n37247;
  assign n39950 = n36254 & n38468;
  assign n39929 = n39973 & n39974;
  assign n36201 = ~n36254;
  assign n39901 = n40009 ^ n40010;
  assign n39991 = ~n40019;
  assign n40011 = ~n40010;
  assign n40058 = n40070 & n40071;
  assign n39994 = n40072 ^ n40073;
  assign n40000 = ~n40095;
  assign n40076 = ~n40096;
  assign n39019 = ~n40097;
  assign n40085 = n36660 & n39016;
  assign n40094 = n40110 & n40111;
  assign n40098 = n40133 & n40134;
  assign n39833 = ~n39908;
  assign n39877 = n39909 & n39910;
  assign n39800 = n38449 ^ n38439;
  assign n39890 = n39929 ^ n39930;
  assign n39937 = n36201 & n39949;
  assign n38471 = ~n39950;
  assign n39912 = ~n39929;
  assign n39975 = n39901 & n37213;
  assign n39981 = n39991 & n39992;
  assign n39976 = ~n39901;
  assign n39914 = n40011 & n40012;
  assign n40041 = n39994 & n15251;
  assign n40039 = ~n40058;
  assign n40042 = ~n39994;
  assign n39922 = n40076 & n40077;
  assign n39037 = ~n40085;
  assign n40074 = ~n40094;
  assign n40059 = n40098 ^ n40099;
  assign n40100 = ~n40098;
  assign n39831 = n39877 ^ n39878;
  assign n39815 = n39890 ^ n39891;
  assign n39881 = n39800 & n39892;
  assign n39876 = ~n39877;
  assign n39882 = ~n39800;
  assign n39900 = n39911 & n39912;
  assign n38489 = ~n39937;
  assign n39894 = ~n39975;
  assign n39956 = n39976 & n37236;
  assign n39931 = ~n39981;
  assign n39917 = ~n39914;
  assign n39993 = n40039 & n40040;
  assign n39996 = ~n40041;
  assign n40020 = n40042 & n402;
  assign n39934 = ~n39922;
  assign n36509 = n37763 ^ n40059;
  assign n40043 = n40074 & n40075;
  assign n40086 = n40100 & n40101;
  assign n39813 = n162 ^ n39831;
  assign n39853 = n39815 & n17182;
  assign n39865 = n39875 & n39876;
  assign n39854 = ~n39815;
  assign n39802 = ~n39881;
  assign n39866 = n39882 & n39836;
  assign n39879 = ~n39900;
  assign n39902 = n39931 ^ n37213;
  assign n39932 = ~n39956;
  assign n39957 = n39993 ^ n39994;
  assign n39995 = ~n39993;
  assign n39959 = ~n40020;
  assign n39998 = n40043 ^ n40044;
  assign n40022 = n36509 & n38884;
  assign n40023 = n36509 & n40047;
  assign n36643 = ~n36509;
  assign n40045 = ~n40043;
  assign n40060 = ~n40086;
  assign n38407 = n39812 ^ n39813;
  assign n39726 = n39813 & n39812;
  assign n39810 = ~n39853;
  assign n39834 = n39854 & n161;
  assign n39832 = ~n39865;
  assign n39838 = ~n39866;
  assign n39835 = n39879 & n39880;
  assign n36167 = n39901 ^ n39902;
  assign n39913 = n39931 & n39932;
  assign n39915 = n402 ^ n39957;
  assign n39982 = n39995 & n39996;
  assign n39919 = n39997 ^ n39998;
  assign n40001 = ~n40022;
  assign n38980 = ~n40023;
  assign n40013 = n36643 & n40024;
  assign n40021 = n40045 & n40046;
  assign n40025 = n40060 & n40061;
  assign n39763 = ~n38407;
  assign n39729 = ~n39726;
  assign n39814 = n39832 & n39833;
  assign n39761 = ~n39834;
  assign n39799 = n39835 ^ n39836;
  assign n39852 = n36167 & n39864;
  assign n39837 = ~n39835;
  assign n38418 = n36167 ^ n37213;
  assign n36133 = ~n36167;
  assign n39893 = ~n39913;
  assign n39816 = n39914 ^ n39915;
  assign n39916 = ~n39915;
  assign n39961 = n39919 & n401;
  assign n39958 = ~n39982;
  assign n39960 = ~n39919;
  assign n39859 = n40001 & n40002;
  assign n39001 = ~n40013;
  assign n39999 = ~n40021;
  assign n39983 = n40025 ^ n40026;
  assign n40027 = ~n40025;
  assign n39721 = n39799 ^ n39800;
  assign n39764 = n39814 ^ n39815;
  assign n39811 = ~n39814;
  assign n39736 = n38418 ^ n38403;
  assign n39825 = n39837 & n39838;
  assign n38437 = ~n39852;
  assign n39851 = n36133 & n38452;
  assign n39855 = n39893 & n39894;
  assign n39883 = n39816 & n37177;
  assign n39884 = ~n39816;
  assign n39840 = n39916 & n39917;
  assign n39918 = n39958 & n39959;
  assign n39941 = n39960 & n15210;
  assign n39887 = ~n39961;
  assign n39968 = n39859 & n39821;
  assign n39964 = ~n39859;
  assign n39977 = n39001 & n38980;
  assign n36439 = n39983 ^ n37690;
  assign n39962 = n39999 & n40000;
  assign n40014 = n40027 & n40028;
  assign n39727 = n161 ^ n39764;
  assign n39759 = n39721 & n160;
  assign n39758 = ~n39721;
  assign n39789 = n39736 & n39766;
  assign n39798 = n39810 & n39811;
  assign n39787 = ~n39736;
  assign n39801 = ~n39825;
  assign n38454 = ~n39851;
  assign n39817 = n39855 ^ n37203;
  assign n39857 = ~n39855;
  assign n39856 = ~n39883;
  assign n39867 = n39884 & n37203;
  assign n39843 = ~n39840;
  assign n39885 = n39918 ^ n39919;
  assign n39920 = ~n39918;
  assign n39921 = ~n39941;
  assign n39923 = n39962 ^ n39963;
  assign n39942 = n39964 & n39965;
  assign n39861 = ~n39968;
  assign n39944 = n36439 & n38853;
  assign n39945 = n36439 & n39970;
  assign n39969 = n39962 & n39963;
  assign n38999 = ~n39977;
  assign n36603 = ~n36439;
  assign n39966 = ~n39962;
  assign n39984 = ~n40014;
  assign n38374 = n39726 ^ n39727;
  assign n39728 = ~n39727;
  assign n39744 = n39758 & n17111;
  assign n39687 = ~n39759;
  assign n39776 = n39787 & n39788;
  assign n39767 = ~n39789;
  assign n39760 = ~n39798;
  assign n39765 = n39801 & n39802;
  assign n36105 = n39816 ^ n39817;
  assign n39839 = n39856 & n39857;
  assign n39819 = ~n39867;
  assign n39841 = n401 ^ n39885;
  assign n39903 = n39920 & n39921;
  assign n39845 = n39922 ^ n39923;
  assign n39823 = ~n39942;
  assign n39925 = ~n39944;
  assign n39935 = n36603 & n38966;
  assign n38948 = ~n39945;
  assign n39943 = n39966 & n39967;
  assign n39933 = ~n39969;
  assign n39946 = n39984 & n39985;
  assign n39683 = ~n38374;
  assign n39646 = n39728 & n39729;
  assign n39722 = ~n39744;
  assign n39720 = n39760 & n39761;
  assign n39737 = n39765 ^ n39766;
  assign n39762 = n36105 & n38407;
  assign n39725 = ~n39776;
  assign n38389 = n36105 ^ n37203;
  assign n39768 = ~n39765;
  assign n36071 = ~n36105;
  assign n39818 = ~n39839;
  assign n39739 = n39840 ^ n39841;
  assign n39842 = ~n39841;
  assign n39888 = n39845 & n15157;
  assign n39886 = ~n39903;
  assign n39889 = ~n39845;
  assign n39741 = n39925 & n39926;
  assign n39924 = n39933 & n39934;
  assign n38968 = ~n39935;
  assign n39896 = ~n39943;
  assign n39904 = n39946 ^ n37720;
  assign n39947 = ~n39946;
  assign n39649 = ~n39646;
  assign n39685 = n39720 ^ n39721;
  assign n39651 = n39736 ^ n39737;
  assign n39628 = n38389 ^ n38371;
  assign n39723 = ~n39720;
  assign n38410 = ~n39762;
  assign n39745 = n36071 & n39763;
  assign n39746 = n39767 & n39768;
  assign n39777 = n39818 & n39819;
  assign n39804 = n39739 & n37143;
  assign n39803 = ~n39739;
  assign n39771 = n39842 & n39843;
  assign n39844 = n39886 & n39887;
  assign n39847 = ~n39888;
  assign n39868 = n39889 & n400;
  assign n39751 = ~n39741;
  assign n36468 = n39904 ^ n39905;
  assign n39895 = ~n39924;
  assign n39936 = n39947 & n39948;
  assign n39647 = n160 ^ n39685;
  assign n39688 = n39651 & n17044;
  assign n39689 = ~n39651;
  assign n39705 = n39628 & n39682;
  assign n39708 = n39722 & n39723;
  assign n39706 = ~n39628;
  assign n38423 = ~n39745;
  assign n39724 = ~n39746;
  assign n39738 = n39777 ^ n37168;
  assign n39769 = ~n39777;
  assign n39790 = n39803 & n37168;
  assign n39731 = ~n39804;
  assign n39805 = n39844 ^ n39845;
  assign n39846 = ~n39844;
  assign n39807 = ~n39868;
  assign n39869 = n36468 & n38816;
  assign n39870 = n36468 & n38931;
  assign n39858 = n39895 & n39896;
  assign n36366 = ~n36468;
  assign n39906 = ~n39936;
  assign n38339 = n39646 ^ n39647;
  assign n39648 = ~n39647;
  assign n39653 = ~n39688;
  assign n39668 = n39689 & n175;
  assign n39617 = ~n39705;
  assign n39698 = n39706 & n39707;
  assign n39686 = ~n39708;
  assign n39709 = n39724 & n39725;
  assign n36047 = n39738 ^ n39739;
  assign n39770 = ~n39790;
  assign n39772 = n400 ^ n39805;
  assign n39826 = n39846 & n39847;
  assign n39820 = n39858 ^ n39859;
  assign n39848 = ~n39869;
  assign n38913 = ~n39870;
  assign n39862 = n36366 & n39871;
  assign n39860 = ~n39858;
  assign n39872 = n39906 & n39907;
  assign n39607 = ~n38339;
  assign n39567 = n39648 & n39649;
  assign n39611 = ~n39668;
  assign n39667 = n36047 & n39683;
  assign n39650 = n39686 & n39687;
  assign n39662 = ~n39698;
  assign n38354 = n37143 ^ n36047;
  assign n39661 = ~n39709;
  assign n36014 = ~n36047;
  assign n39747 = n39769 & n39770;
  assign n39655 = n39771 ^ n39772;
  assign n39693 = n39772 & n39771;
  assign n39733 = n39820 ^ n39821;
  assign n39806 = ~n39826;
  assign n39633 = n39848 & n39849;
  assign n39850 = n39860 & n39861;
  assign n38933 = ~n39862;
  assign n39828 = n39872 ^ n37617;
  assign n39873 = ~n39872;
  assign n39570 = ~n39567;
  assign n39609 = n39650 ^ n39651;
  assign n39542 = n38354 ^ n38344;
  assign n39645 = n39661 & n39662;
  assign n38377 = ~n39667;
  assign n39652 = ~n39650;
  assign n39629 = n39661 ^ n39682;
  assign n39684 = n36014 & n38374;
  assign n39730 = ~n39747;
  assign n39696 = ~n39693;
  assign n39778 = n39733 & n15109;
  assign n39773 = n39806 & n39807;
  assign n39779 = ~n39733;
  assign n39809 = n39633 & n39824;
  assign n39808 = ~n39633;
  assign n36333 = n39827 ^ n39828;
  assign n39822 = ~n39850;
  assign n39863 = n39873 & n39874;
  assign n39568 = n175 ^ n39609;
  assign n39572 = n39628 ^ n39629;
  assign n39619 = n39542 & n39630;
  assign n39618 = ~n39542;
  assign n39616 = ~n39645;
  assign n39627 = n39652 & n39653;
  assign n38392 = ~n39684;
  assign n39690 = n39730 & n39731;
  assign n39732 = n415 ^ n39773;
  assign n39748 = ~n39778;
  assign n39774 = n39779 & n415;
  assign n39749 = ~n39773;
  assign n39792 = n39808 & n39673;
  assign n39675 = ~n39809;
  assign n39793 = n36333 & n38878;
  assign n39780 = n39822 & n39823;
  assign n36394 = ~n36333;
  assign n39829 = ~n39863;
  assign n38303 = n39567 ^ n39568;
  assign n39569 = ~n39568;
  assign n39592 = n39572 & n174;
  assign n39591 = ~n39572;
  assign n39581 = n39616 & n39617;
  assign n39612 = n39618 & n39582;
  assign n39545 = ~n39619;
  assign n39610 = ~n39627;
  assign n39654 = n39690 ^ n37113;
  assign n39692 = n39690 & n37113;
  assign n39691 = ~n39690;
  assign n39694 = n39732 ^ n39733;
  assign n39740 = n39748 & n39749;
  assign n39711 = ~n39774;
  assign n39742 = n39780 ^ n39781;
  assign n39783 = n39780 & n39791;
  assign n39636 = ~n39792;
  assign n39784 = n36394 & n38837;
  assign n38899 = ~n39793;
  assign n39785 = n36394 & n39794;
  assign n39782 = ~n39780;
  assign n39795 = n39829 & n39830;
  assign n39522 = ~n38303;
  assign n39499 = n39569 & n39570;
  assign n39541 = n39581 ^ n39582;
  assign n39580 = n39591 & n17004;
  assign n39524 = ~n39592;
  assign n39571 = n39610 & n39611;
  assign n39584 = ~n39581;
  assign n39583 = ~n39612;
  assign n35969 = n39654 ^ n39655;
  assign n39669 = n39691 & n37110;
  assign n39663 = ~n39692;
  assign n39546 = n39693 ^ n39694;
  assign n39695 = ~n39694;
  assign n39710 = ~n39740;
  assign n39671 = n39741 ^ n39742;
  assign n39775 = n39782 & n39781;
  assign n39750 = ~n39783;
  assign n39752 = ~n39784;
  assign n38881 = ~n39785;
  assign n39755 = n39795 ^ n37567;
  assign n39796 = ~n39795;
  assign n39475 = n39541 ^ n39542;
  assign n39502 = ~n39499;
  assign n39535 = n39571 ^ n39572;
  assign n39552 = ~n39580;
  assign n39573 = n39583 & n39584;
  assign n39553 = ~n39571;
  assign n38322 = n37110 ^ n35969;
  assign n39608 = n35969 & n38339;
  assign n35994 = ~n35969;
  assign n39656 = n39663 & n39655;
  assign n39657 = n39546 & n37083;
  assign n39621 = ~n39669;
  assign n39658 = ~n39546;
  assign n39593 = n39695 & n39696;
  assign n39670 = n39710 & n39711;
  assign n39700 = n39671 & n414;
  assign n39699 = ~n39671;
  assign n39743 = n39750 & n39751;
  assign n39556 = n39752 & n39753;
  assign n36258 = n39754 ^ n39755;
  assign n39713 = ~n39775;
  assign n39786 = n39796 & n39797;
  assign n39513 = n39475 & n173;
  assign n39500 = n174 ^ n39535;
  assign n39512 = ~n39475;
  assign n39543 = n39552 & n39553;
  assign n39544 = ~n39573;
  assign n39474 = n38322 ^ n38270;
  assign n39590 = n35994 & n39607;
  assign n38341 = ~n39608;
  assign n39620 = ~n39656;
  assign n39588 = ~n39657;
  assign n39631 = n39658 & n37053;
  assign n39596 = ~n39593;
  assign n39632 = n39670 ^ n39671;
  assign n39665 = ~n39670;
  assign n39697 = n39699 & n15067;
  assign n39623 = ~n39700;
  assign n39715 = n39556 & n39734;
  assign n39716 = n36258 & n39735;
  assign n39712 = ~n39743;
  assign n39714 = ~n39556;
  assign n36331 = ~n36258;
  assign n39756 = ~n39786;
  assign n38264 = n39499 ^ n39500;
  assign n39504 = n39512 & n16960;
  assign n39450 = ~n39513;
  assign n39501 = ~n39500;
  assign n39523 = ~n39543;
  assign n39515 = n39544 & n39545;
  assign n38357 = ~n39590;
  assign n39589 = n39620 & n39621;
  assign n39549 = ~n39631;
  assign n39594 = n414 ^ n39632;
  assign n39664 = ~n39697;
  assign n39672 = n39712 & n39713;
  assign n39701 = n39714 & n39600;
  assign n39602 = ~n39715;
  assign n39702 = n36331 & n38848;
  assign n38864 = ~n39716;
  assign n39703 = n36331 & n38792;
  assign n39717 = n39756 & n39757;
  assign n39447 = ~n38264;
  assign n39419 = n39501 & n39502;
  assign n39471 = ~n39504;
  assign n39473 = n39515 ^ n39516;
  assign n39514 = n39523 & n39524;
  assign n39519 = n39515 & n39516;
  assign n39517 = ~n39515;
  assign n39547 = n39589 ^ n37053;
  assign n39477 = n39593 ^ n39594;
  assign n39587 = ~n39589;
  assign n39595 = ~n39594;
  assign n39659 = n39664 & n39665;
  assign n39634 = n39672 ^ n39673;
  assign n39674 = ~n39672;
  assign n39559 = ~n39701;
  assign n38851 = ~n39702;
  assign n39676 = ~n39703;
  assign n39678 = n39717 ^ n37553;
  assign n39718 = ~n39717;
  assign n39401 = n39473 ^ n39474;
  assign n39472 = ~n39514;
  assign n39505 = n39517 & n39518;
  assign n39483 = ~n39519;
  assign n35959 = n39546 ^ n39547;
  assign n39565 = n39477 & n37050;
  assign n39566 = ~n39477;
  assign n39579 = n39587 & n39588;
  assign n39494 = n39595 & n39596;
  assign n39574 = n39633 ^ n39634;
  assign n39622 = ~n39659;
  assign n39666 = n39674 & n39675;
  assign n39484 = n39676 & n39677;
  assign n36247 = n39678 ^ n39679;
  assign n39704 = n39718 & n39719;
  assign n39467 = n39471 & n39472;
  assign n39448 = n39472 ^ n39475;
  assign n39476 = n39483 & n39474;
  assign n39459 = ~n39505;
  assign n38282 = n35959 ^ n37053;
  assign n39511 = n35959 & n39522;
  assign n35927 = ~n35959;
  assign n39480 = ~n39565;
  assign n39540 = n39566 & n37029;
  assign n39548 = ~n39579;
  assign n39498 = ~n39494;
  assign n39598 = n39574 & n413;
  assign n39613 = n39622 & n39623;
  assign n39597 = ~n39574;
  assign n39638 = n39484 & n39660;
  assign n39639 = n36247 & n38757;
  assign n39640 = n36247 & n38811;
  assign n39635 = ~n39666;
  assign n39637 = ~n39484;
  assign n36186 = ~n36247;
  assign n39680 = ~n39704;
  assign n39420 = n173 ^ n39448;
  assign n39449 = ~n39467;
  assign n39458 = ~n39476;
  assign n39402 = n38282 ^ n38261;
  assign n39503 = n35927 & n38303;
  assign n38305 = ~n39511;
  assign n39509 = ~n39540;
  assign n39510 = n39548 & n39549;
  assign n39585 = n39597 & n15056;
  assign n39526 = ~n39598;
  assign n39555 = ~n39613;
  assign n39599 = n39635 & n39636;
  assign n39624 = n39637 & n39530;
  assign n39532 = ~n39638;
  assign n39614 = ~n39639;
  assign n38814 = ~n39640;
  assign n39625 = n36186 & n39641;
  assign n39642 = n39680 & n39681;
  assign n38223 = n39419 ^ n39420;
  assign n39351 = n39420 & n39419;
  assign n39431 = n39449 & n39450;
  assign n39432 = n39458 & n39459;
  assign n38325 = ~n39503;
  assign n39478 = n39510 ^ n37029;
  assign n39508 = ~n39510;
  assign n39536 = n39555 ^ n39574;
  assign n39554 = ~n39585;
  assign n39557 = n39599 ^ n39600;
  assign n39427 = n39614 & n39615;
  assign n39601 = ~n39599;
  assign n39487 = ~n39624;
  assign n38833 = ~n39625;
  assign n39604 = n39642 ^ n37446;
  assign n39643 = ~n39642;
  assign n39388 = ~n38223;
  assign n39354 = ~n39351;
  assign n39421 = n39431 & n16911;
  assign n39403 = n39432 ^ n39433;
  assign n39414 = ~n39431;
  assign n39436 = n39432 & n39433;
  assign n39434 = ~n39432;
  assign n35915 = n39477 ^ n39478;
  assign n39496 = n39508 & n39509;
  assign n39495 = n413 ^ n39536;
  assign n39550 = n39554 & n39555;
  assign n39493 = n39556 ^ n39557;
  assign n39577 = n39427 & n39464;
  assign n39586 = n39601 & n39602;
  assign n39575 = ~n39427;
  assign n36120 = n39603 ^ n39604;
  assign n39626 = n39643 & n39644;
  assign n39321 = n39402 ^ n39403;
  assign n39381 = n39414 ^ n39401;
  assign n39415 = n39414 & n172;
  assign n39400 = ~n39421;
  assign n39422 = n39434 & n39435;
  assign n39416 = ~n39436;
  assign n38244 = n35915 ^ n37050;
  assign n39446 = n35915 & n38264;
  assign n35883 = ~n35915;
  assign n39481 = n39494 ^ n39495;
  assign n39479 = ~n39496;
  assign n39497 = ~n39495;
  assign n39528 = n39493 & n412;
  assign n39525 = ~n39550;
  assign n39527 = ~n39493;
  assign n39560 = n39575 & n39576;
  assign n39561 = n36120 & n38724;
  assign n39466 = ~n39577;
  assign n39562 = n36120 & n39578;
  assign n39558 = ~n39586;
  assign n36180 = ~n36120;
  assign n39605 = ~n39626;
  assign n39352 = n172 ^ n39381;
  assign n39390 = n39400 & n39401;
  assign n39366 = ~n39415;
  assign n39404 = n39416 & n39402;
  assign n39383 = ~n39422;
  assign n39323 = n38244 ^ n38228;
  assign n38266 = ~n39446;
  assign n39443 = n35883 & n39447;
  assign n39451 = n39479 & n39480;
  assign n39468 = n39481 & n37000;
  assign n39423 = ~n39481;
  assign n39437 = n39497 & n39498;
  assign n39492 = n39525 & n39526;
  assign n39520 = n39527 & n14988;
  assign n39462 = ~n39528;
  assign n39529 = n39558 & n39559;
  assign n39442 = ~n39560;
  assign n39537 = ~n39561;
  assign n38803 = ~n39562;
  assign n39551 = n36180 & n38775;
  assign n39563 = n39605 & n39606;
  assign n39330 = n39351 ^ n39352;
  assign n39353 = ~n39352;
  assign n39365 = ~n39390;
  assign n39382 = ~n39404;
  assign n39391 = n39323 & n39405;
  assign n39392 = ~n39323;
  assign n38286 = ~n39443;
  assign n39424 = n39451 ^ n37000;
  assign n39452 = ~n39451;
  assign n39460 = n39423 & n37061;
  assign n39453 = ~n39468;
  assign n39457 = n39492 ^ n39493;
  assign n39491 = ~n39492;
  assign n39490 = ~n39520;
  assign n39485 = n39529 ^ n39530;
  assign n39376 = n39537 & n39538;
  assign n39531 = ~n39529;
  assign n38782 = ~n39551;
  assign n38748 = n39563 ^ n39564;
  assign n38184 = ~n39330;
  assign n39286 = n39353 & n39354;
  assign n39339 = n39365 & n39366;
  assign n39355 = n39382 & n39383;
  assign n39325 = ~n39391;
  assign n39384 = n39392 & n39356;
  assign n35869 = n39423 ^ n39424;
  assign n39444 = n39452 & n39453;
  assign n39438 = n412 ^ n39457;
  assign n39426 = ~n39460;
  assign n39440 = n39484 ^ n39485;
  assign n39482 = n39490 & n39491;
  assign n39521 = n39531 & n39532;
  assign n39379 = ~n39376;
  assign n39488 = n39533 ^ n38748;
  assign n39534 = n38748 & n39539;
  assign n36148 = ~n38748;
  assign n39309 = n39339 ^ n39321;
  assign n39341 = n39339 & n16887;
  assign n39322 = n39355 ^ n39356;
  assign n39340 = ~n39339;
  assign n39357 = ~n39355;
  assign n39358 = ~n39384;
  assign n38204 = n35869 ^ n37061;
  assign n39389 = n35869 & n38223;
  assign n35838 = ~n35869;
  assign n39394 = n39437 ^ n39438;
  assign n39425 = ~n39444;
  assign n39368 = n39438 & n39437;
  assign n39455 = n39440 & n411;
  assign n39461 = ~n39482;
  assign n39456 = ~n39440;
  assign n38767 = n39488 ^ n39489;
  assign n39486 = ~n39521;
  assign n39506 = ~n39534;
  assign n39287 = n171 ^ n39309;
  assign n39255 = n39322 ^ n39323;
  assign n39331 = n39340 & n171;
  assign n39320 = ~n39341;
  assign n39342 = n39357 & n39358;
  assign n39282 = n38204 ^ n38190;
  assign n39380 = n35838 & n39388;
  assign n38225 = ~n39389;
  assign n39407 = n39394 & n36960;
  assign n39393 = n39425 & n39426;
  assign n39406 = ~n39394;
  assign n39371 = ~n39368;
  assign n39410 = ~n39455;
  assign n39445 = n39456 & n14942;
  assign n39439 = n39461 & n39462;
  assign n39463 = n39486 & n39487;
  assign n39469 = n39506 & n39507;
  assign n39277 = n39286 ^ n39287;
  assign n39234 = n39287 & n39286;
  assign n39310 = n39320 & n39321;
  assign n39297 = ~n39331;
  assign n39324 = ~n39342;
  assign n39333 = n39282 & n39343;
  assign n39332 = ~n39282;
  assign n38248 = ~n39380;
  assign n38165 = n39393 ^ n39394;
  assign n39395 = n39406 & n36991;
  assign n39385 = ~n39407;
  assign n39386 = ~n39393;
  assign n39408 = n39439 ^ n39440;
  assign n39430 = ~n39445;
  assign n39429 = ~n39439;
  assign n39428 = n39463 ^ n39464;
  assign n39305 = n39469 ^ n39470;
  assign n39465 = ~n39463;
  assign n38146 = ~n39277;
  assign n39296 = ~n39310;
  assign n39298 = n39324 & n39325;
  assign n39326 = n39332 & n39299;
  assign n39284 = ~n39333;
  assign n39237 = n38112 ^ n38165;
  assign n35790 = n38165 ^ n36960;
  assign n39367 = n39385 & n39386;
  assign n39360 = ~n39395;
  assign n39369 = n411 ^ n39408;
  assign n39373 = n39427 ^ n39428;
  assign n39418 = n39429 & n39430;
  assign n39454 = n39465 & n39466;
  assign n39278 = n39296 & n39297;
  assign n39281 = n39298 ^ n39299;
  assign n39300 = ~n39298;
  assign n39301 = ~n39326;
  assign n39319 = n35790 & n39330;
  assign n39334 = n39237 & n39260;
  assign n39335 = ~n39237;
  assign n35818 = ~n35790;
  assign n39359 = ~n39367;
  assign n39303 = n39368 ^ n39369;
  assign n39370 = ~n39369;
  assign n39411 = n39373 & n14910;
  assign n39409 = ~n39418;
  assign n39412 = ~n39373;
  assign n39441 = ~n39454;
  assign n39254 = n170 ^ n39278;
  assign n39218 = n39281 ^ n39282;
  assign n39280 = n39278 & n16859;
  assign n39279 = ~n39278;
  assign n39288 = n39300 & n39301;
  assign n39308 = n35818 & n38184;
  assign n38208 = ~n39319;
  assign n39262 = ~n39334;
  assign n39327 = n39335 & n39336;
  assign n39328 = n39359 & n39360;
  assign n39344 = n39303 & n36904;
  assign n39345 = ~n39303;
  assign n39313 = n39370 & n39371;
  assign n39372 = n39409 & n39410;
  assign n39375 = ~n39411;
  assign n39396 = n39412 & n410;
  assign n39413 = n39441 & n39442;
  assign n39235 = n39254 ^ n39255;
  assign n39258 = n39218 & n169;
  assign n39257 = ~n39218;
  assign n39267 = n39279 & n170;
  assign n39264 = ~n39280;
  assign n39283 = ~n39288;
  assign n38187 = ~n39308;
  assign n39239 = ~n39327;
  assign n39302 = n39328 ^ n36978;
  assign n39311 = ~n39328;
  assign n39290 = ~n39344;
  assign n39337 = n39345 & n36978;
  assign n39346 = n39372 ^ n39373;
  assign n39374 = ~n39372;
  assign n39348 = ~n39396;
  assign n39377 = n39413 ^ n39399;
  assign n39397 = n39413 & n39417;
  assign n39398 = ~n39413;
  assign n38104 = n39234 ^ n39235;
  assign n39180 = n39235 & n39234;
  assign n39246 = n39257 & n16793;
  assign n39202 = ~n39258;
  assign n39256 = n39264 & n39255;
  assign n39244 = ~n39267;
  assign n39259 = n39283 & n39284;
  assign n35714 = n39302 ^ n39303;
  assign n39312 = ~n39337;
  assign n39314 = n410 ^ n39346;
  assign n39363 = n39374 & n39375;
  assign n39316 = n39376 ^ n39377;
  assign n39378 = ~n39397;
  assign n39387 = n39398 & n39399;
  assign n39208 = ~n38104;
  assign n39183 = ~n39180;
  assign n39220 = ~n39246;
  assign n39243 = ~n39256;
  assign n39236 = n39259 ^ n39260;
  assign n39263 = n35714 & n38146;
  assign n39261 = ~n39259;
  assign n38126 = n35714 ^ n36904;
  assign n35795 = ~n35714;
  assign n39306 = n39311 & n39312;
  assign n39269 = n39313 ^ n39314;
  assign n39272 = n39314 & n39313;
  assign n39350 = n39316 & n409;
  assign n39347 = ~n39363;
  assign n39349 = ~n39316;
  assign n39364 = n39378 & n39379;
  assign n39362 = ~n39387;
  assign n39185 = n39236 ^ n39237;
  assign n39217 = n39243 & n39244;
  assign n39247 = n39261 & n39262;
  assign n39214 = n38126 ^ n38073;
  assign n38148 = ~n39263;
  assign n39266 = n35795 & n39277;
  assign n39291 = n39269 & n36865;
  assign n39289 = ~n39306;
  assign n39292 = ~n39269;
  assign n39315 = n39347 & n39348;
  assign n39338 = n39349 & n14879;
  assign n39295 = ~n39350;
  assign n39361 = ~n39364;
  assign n39200 = n39217 ^ n39218;
  assign n39211 = n39185 & n16739;
  assign n39212 = ~n39185;
  assign n39219 = ~n39217;
  assign n39242 = n39214 & n39197;
  assign n39238 = ~n39247;
  assign n39240 = ~n39214;
  assign n38169 = ~n39266;
  assign n39268 = n39289 & n39290;
  assign n39249 = ~n39291;
  assign n39285 = n39292 & n36963;
  assign n39293 = n39315 ^ n39316;
  assign n39317 = ~n39315;
  assign n39318 = ~n39338;
  assign n39329 = n39361 & n39362;
  assign n39181 = n169 ^ n39200;
  assign n39187 = ~n39211;
  assign n39204 = n39212 & n168;
  assign n39210 = n39219 & n39220;
  assign n39213 = n39238 & n39239;
  assign n39224 = n39240 & n39241;
  assign n39216 = ~n39242;
  assign n38085 = n39268 ^ n39269;
  assign n39270 = ~n39268;
  assign n39271 = ~n39285;
  assign n39273 = n409 ^ n39293;
  assign n39307 = n39317 & n39318;
  assign n39304 = n408 ^ n39329;
  assign n38065 = n39180 ^ n39181;
  assign n39182 = ~n39181;
  assign n39166 = ~n39204;
  assign n39201 = ~n39210;
  assign n39196 = n39213 ^ n39214;
  assign n39215 = ~n39213;
  assign n39199 = ~n39224;
  assign n35648 = n38085 ^ n36963;
  assign n39177 = n38085 ^ n38015;
  assign n39265 = n39270 & n39271;
  assign n39229 = n39272 ^ n39273;
  assign n39274 = ~n39273;
  assign n39276 = n39304 ^ n39305;
  assign n39294 = ~n39307;
  assign n39163 = ~n38065;
  assign n39147 = n39182 & n39183;
  assign n39133 = n39196 ^ n39197;
  assign n39184 = n39201 & n39202;
  assign n39203 = n35648 & n39208;
  assign n39205 = n39215 & n39216;
  assign n39225 = n39177 & n39159;
  assign n35717 = ~n35648;
  assign n39226 = ~n39177;
  assign n39250 = n39229 & n36877;
  assign n39248 = ~n39265;
  assign n39251 = ~n39229;
  assign n39252 = n39274 & n39272;
  assign n39275 = n39294 & n39295;
  assign n39164 = n39184 ^ n39185;
  assign n39174 = n39133 & n16715;
  assign n39175 = ~n39133;
  assign n39186 = ~n39184;
  assign n38107 = ~n39203;
  assign n39198 = ~n39205;
  assign n39209 = n35717 & n38104;
  assign n39179 = ~n39225;
  assign n39221 = n39226 & n39227;
  assign n39228 = n39248 & n39249;
  assign n39231 = ~n39250;
  assign n39245 = n39251 & n36831;
  assign n39253 = n39275 ^ n39276;
  assign n39148 = n168 ^ n39164;
  assign n39151 = ~n39174;
  assign n39167 = n39175 & n183;
  assign n39173 = n39186 & n39187;
  assign n39176 = n39198 & n39199;
  assign n38131 = ~n39209;
  assign n39161 = ~n39221;
  assign n38047 = n39228 ^ n39229;
  assign n39230 = ~n39228;
  assign n39207 = ~n39245;
  assign n39169 = n39252 ^ n39253;
  assign n38029 = n39147 ^ n39148;
  assign n39107 = n39148 & n39147;
  assign n39135 = ~n39167;
  assign n39165 = ~n39173;
  assign n39158 = n39176 ^ n39177;
  assign n39178 = ~n39176;
  assign n35574 = n38047 ^ n36877;
  assign n39144 = n38047 ^ n38026;
  assign n39222 = n39230 & n39231;
  assign n39232 = n39169 & n36892;
  assign n39233 = ~n39169;
  assign n39131 = ~n38029;
  assign n39110 = n39158 ^ n39159;
  assign n39157 = n35574 & n39163;
  assign n39149 = n39165 & n39166;
  assign n39168 = n39178 & n39179;
  assign n39190 = n39144 & n39125;
  assign n35653 = ~n35574;
  assign n39191 = ~n39144;
  assign n39206 = ~n39222;
  assign n39172 = ~n39232;
  assign n39223 = n39233 & n36814;
  assign n39132 = n183 ^ n39149;
  assign n39141 = n39110 & n16633;
  assign n39142 = ~n39110;
  assign n38089 = ~n39157;
  assign n39150 = ~n39149;
  assign n39162 = n35653 & n38065;
  assign n39160 = ~n39168;
  assign n39146 = ~n39190;
  assign n39188 = n39191 & n39192;
  assign n39193 = n39206 & n39207;
  assign n39195 = ~n39223;
  assign n39108 = n39132 ^ n39133;
  assign n39112 = ~n39141;
  assign n39136 = n39142 & n182;
  assign n39140 = n39150 & n39151;
  assign n39143 = n39160 & n39161;
  assign n38068 = ~n39162;
  assign n39127 = ~n39188;
  assign n39170 = n39193 ^ n36892;
  assign n39194 = ~n39193;
  assign n37991 = n39107 ^ n39108;
  assign n39072 = n39108 & n39107;
  assign n39093 = ~n39136;
  assign n39134 = ~n39140;
  assign n39124 = n39143 ^ n39144;
  assign n39145 = ~n39143;
  assign n35538 = n39169 ^ n39170;
  assign n39189 = n39194 & n39195;
  assign n39089 = ~n37991;
  assign n39075 = ~n39072;
  assign n39077 = n39124 ^ n39125;
  assign n39123 = n35538 & n39131;
  assign n39109 = n39134 & n39135;
  assign n39137 = n39145 & n39146;
  assign n38009 = n36892 ^ n35538;
  assign n35586 = ~n35538;
  assign n39171 = ~n39189;
  assign n39091 = n39109 ^ n39110;
  assign n39102 = n39077 & n16558;
  assign n39103 = ~n39077;
  assign n38051 = ~n39123;
  assign n39111 = ~n39109;
  assign n39130 = n35586 & n38029;
  assign n39126 = ~n39137;
  assign n39086 = n38009 ^ n37959;
  assign n39153 = n39171 & n39172;
  assign n39073 = n182 ^ n39091;
  assign n39079 = ~n39102;
  assign n39096 = n39103 & n181;
  assign n39101 = n39111 & n39112;
  assign n39104 = n39126 & n39127;
  assign n39118 = n39086 & n39105;
  assign n38032 = ~n39130;
  assign n39116 = ~n39086;
  assign n37971 = n39153 ^ n39154;
  assign n39155 = ~n39153;
  assign n37952 = n39072 ^ n39073;
  assign n39074 = ~n39073;
  assign n39058 = ~n39096;
  assign n39092 = ~n39101;
  assign n39085 = n39104 ^ n39105;
  assign n39097 = ~n39104;
  assign n39113 = n39116 & n39117;
  assign n39083 = ~n39118;
  assign n35469 = n36812 ^ n37971;
  assign n39046 = n37971 ^ n37918;
  assign n39152 = n39155 & n39156;
  assign n39055 = ~n37952;
  assign n39038 = n39074 & n39075;
  assign n39041 = n39085 ^ n39086;
  assign n39084 = n35469 & n39089;
  assign n39076 = n39092 & n39093;
  assign n39098 = ~n39113;
  assign n39119 = n39046 & n39128;
  assign n35516 = ~n35469;
  assign n39120 = ~n39046;
  assign n39138 = ~n39152;
  assign n39044 = ~n39038;
  assign n39056 = n39076 ^ n39077;
  assign n39067 = n39041 & n16510;
  assign n39068 = ~n39041;
  assign n38013 = ~n39084;
  assign n39078 = ~n39076;
  assign n39090 = n35516 & n37991;
  assign n39094 = n39097 & n39098;
  assign n39048 = ~n39119;
  assign n39114 = n39120 & n39062;
  assign n39129 = n39138 & n39139;
  assign n39039 = n181 ^ n39056;
  assign n39043 = ~n39067;
  assign n39060 = n39068 & n180;
  assign n39066 = n39078 & n39079;
  assign n37994 = ~n39090;
  assign n39082 = ~n39094;
  assign n39064 = ~n39114;
  assign n39122 = n39129 & n36723;
  assign n39121 = ~n39129;
  assign n37935 = n39038 ^ n39039;
  assign n39002 = n39039 & n39044;
  assign n39024 = ~n39060;
  assign n39057 = ~n39066;
  assign n39061 = n39082 & n39083;
  assign n39115 = n39121 & n36769;
  assign n39100 = ~n39122;
  assign n39020 = ~n37935;
  assign n39005 = ~n39002;
  assign n39040 = n39057 & n39058;
  assign n39045 = n39061 ^ n39062;
  assign n39063 = ~n39061;
  assign n39099 = n39100 & n39106;
  assign n39088 = ~n39115;
  assign n39022 = n39040 ^ n39041;
  assign n39007 = n39045 ^ n39046;
  assign n39042 = ~n39040;
  assign n39059 = n39063 & n39064;
  assign n39087 = ~n39099;
  assign n39095 = n39088 & n39100;
  assign n39003 = n180 ^ n39022;
  assign n39030 = n39007 & n179;
  assign n39034 = n39042 & n39043;
  assign n39029 = ~n39007;
  assign n39047 = ~n39059;
  assign n39069 = n39087 & n39088;
  assign n39081 = ~n39095;
  assign n38988 = n39002 ^ n39003;
  assign n39004 = ~n39003;
  assign n39025 = n39029 & n16437;
  assign n38984 = ~n39030;
  assign n39023 = ~n39034;
  assign n39031 = n39047 & n39048;
  assign n39051 = n39069 ^ n36710;
  assign n35434 = n39080 ^ n39081;
  assign n39070 = ~n39069;
  assign n37874 = ~n38988;
  assign n38969 = n39004 & n39005;
  assign n39006 = n39023 & n39024;
  assign n39009 = ~n39025;
  assign n39012 = n39031 ^ n39028;
  assign n39010 = ~n39031;
  assign n35359 = n39051 ^ n39052;
  assign n39049 = n35434 & n39055;
  assign n37932 = n36723 ^ n35434;
  assign n39065 = n39070 & n39071;
  assign n35395 = ~n35434;
  assign n38982 = n39006 ^ n39007;
  assign n39008 = ~n39006;
  assign n39014 = n35359 & n39020;
  assign n37893 = n35359 ^ n36672;
  assign n39013 = n37932 ^ n37881;
  assign n35319 = ~n35359;
  assign n37955 = ~n39049;
  assign n39050 = n35395 & n37952;
  assign n39053 = ~n39065;
  assign n38970 = n179 ^ n38982;
  assign n38993 = n39008 & n39009;
  assign n38972 = n39012 ^ n39013;
  assign n37914 = ~n39014;
  assign n38944 = n37893 ^ n37879;
  assign n39021 = n35319 & n37935;
  assign n39026 = n39013 & n39032;
  assign n39027 = ~n39013;
  assign n37976 = ~n39050;
  assign n39035 = n39053 & n39054;
  assign n38956 = n38969 ^ n38970;
  assign n38934 = n38970 & n38969;
  assign n38983 = ~n38993;
  assign n38990 = n38972 & n178;
  assign n38989 = ~n38972;
  assign n38994 = n38944 & n38964;
  assign n38995 = ~n38944;
  assign n37937 = ~n39021;
  assign n38987 = ~n39026;
  assign n39015 = n39027 & n39028;
  assign n39017 = n39035 ^ n36613;
  assign n39036 = ~n39035;
  assign n37836 = ~n38956;
  assign n38971 = n38983 & n38984;
  assign n38985 = n38989 & n16378;
  assign n38952 = ~n38990;
  assign n38954 = ~n38994;
  assign n38991 = n38995 & n38996;
  assign n39011 = ~n39015;
  assign n35290 = n39016 ^ n39017;
  assign n39033 = n39036 & n39037;
  assign n38950 = n38971 ^ n38972;
  assign n38973 = ~n38971;
  assign n38977 = n35290 & n37874;
  assign n38974 = ~n38985;
  assign n38976 = ~n38991;
  assign n37855 = n35290 ^ n36613;
  assign n38997 = n39010 & n39011;
  assign n35239 = ~n35290;
  assign n39018 = ~n39033;
  assign n38935 = n178 ^ n38950;
  assign n38959 = n38973 & n38974;
  assign n37876 = ~n38977;
  assign n38916 = n37855 ^ n37841;
  assign n38981 = n35239 & n38988;
  assign n38986 = ~n38997;
  assign n38998 = n39018 & n39019;
  assign n38919 = n38934 ^ n38935;
  assign n38889 = n38935 & n38934;
  assign n38951 = ~n38959;
  assign n38961 = n38916 & n38975;
  assign n38960 = ~n38916;
  assign n37897 = ~n38981;
  assign n38978 = n38986 & n38987;
  assign n35119 = n38998 ^ n38999;
  assign n39000 = ~n38998;
  assign n37795 = ~n38919;
  assign n38942 = n35119 & n37836;
  assign n38923 = n38951 & n38952;
  assign n38957 = n38960 & n38937;
  assign n38918 = ~n38961;
  assign n38963 = ~n38978;
  assign n37816 = n35119 ^ n36509;
  assign n35213 = ~n35119;
  assign n38992 = n39000 & n39001;
  assign n37838 = ~n38942;
  assign n38910 = ~n38923;
  assign n38949 = n35213 & n38956;
  assign n38938 = ~n38957;
  assign n38903 = n37816 ^ n37792;
  assign n38943 = n38963 ^ n38964;
  assign n38962 = n38976 & n38963;
  assign n38979 = ~n38992;
  assign n38924 = n38943 ^ n38944;
  assign n37859 = ~n38949;
  assign n38946 = n38903 & n38955;
  assign n38945 = ~n38903;
  assign n38953 = ~n38962;
  assign n38965 = n38979 & n38980;
  assign n38909 = n38923 ^ n38924;
  assign n38926 = n38924 & n177;
  assign n38925 = ~n38924;
  assign n38941 = n38945 & n38884;
  assign n38905 = ~n38946;
  assign n38936 = n38953 & n38954;
  assign n37776 = n38965 ^ n38966;
  assign n38967 = ~n38965;
  assign n38890 = n177 ^ n38909;
  assign n38920 = n38925 & n16277;
  assign n38892 = ~n38926;
  assign n38915 = n38936 ^ n38937;
  assign n38886 = ~n38941;
  assign n38939 = ~n38936;
  assign n38868 = n37776 ^ n37761;
  assign n35040 = n37776 ^ n36439;
  assign n38958 = n38967 & n38968;
  assign n38882 = n38889 ^ n38890;
  assign n38843 = n38890 & n38889;
  assign n38908 = n35040 & n37795;
  assign n38875 = n38915 ^ n38916;
  assign n38911 = ~n38920;
  assign n38927 = n38938 & n38939;
  assign n38928 = n38868 & n38940;
  assign n38929 = ~n38868;
  assign n35135 = ~n35040;
  assign n38947 = ~n38958;
  assign n37755 = ~n38882;
  assign n38901 = n38875 & n176;
  assign n37798 = ~n38908;
  assign n38907 = n38910 & n38911;
  assign n38900 = ~n38875;
  assign n38914 = n35135 & n38919;
  assign n38917 = ~n38927;
  assign n38870 = ~n38928;
  assign n38921 = n38929 & n38853;
  assign n38930 = n38947 & n38948;
  assign n38893 = n38900 & n16229;
  assign n38859 = ~n38901;
  assign n38891 = ~n38907;
  assign n37821 = ~n38914;
  assign n38902 = n38917 & n38918;
  assign n38855 = ~n38921;
  assign n37734 = n38930 ^ n38931;
  assign n38932 = ~n38930;
  assign n38874 = n38891 & n38892;
  assign n38876 = ~n38893;
  assign n38883 = n38902 ^ n38903;
  assign n38904 = ~n38902;
  assign n38839 = n37734 ^ n37642;
  assign n34964 = n36468 ^ n37734;
  assign n38922 = n38932 & n38933;
  assign n38857 = n38874 ^ n38875;
  assign n38873 = n34964 & n38882;
  assign n38824 = n38883 ^ n38884;
  assign n38877 = ~n38874;
  assign n38894 = n38904 & n38905;
  assign n38895 = n38839 & n38906;
  assign n38896 = ~n38839;
  assign n35045 = ~n34964;
  assign n38912 = ~n38922;
  assign n38844 = n176 ^ n38857;
  assign n38866 = n38824 & n191;
  assign n38871 = n35045 & n37755;
  assign n37780 = ~n38873;
  assign n38872 = n38876 & n38877;
  assign n38865 = ~n38824;
  assign n38885 = ~n38894;
  assign n38841 = ~n38895;
  assign n38887 = n38896 & n38816;
  assign n38897 = n38912 & n38913;
  assign n38834 = n38843 ^ n38844;
  assign n38805 = n38844 & n38843;
  assign n38860 = n38865 & n16084;
  assign n38826 = ~n38866;
  assign n37758 = ~n38871;
  assign n38858 = ~n38872;
  assign n38867 = n38885 & n38886;
  assign n38818 = ~n38887;
  assign n38879 = n38897 ^ n36333;
  assign n38898 = ~n38897;
  assign n37708 = ~n38834;
  assign n38845 = n38858 & n38859;
  assign n38846 = ~n38860;
  assign n38852 = n38867 ^ n38868;
  assign n38869 = ~n38867;
  assign n34968 = n38878 ^ n38879;
  assign n38888 = n38898 & n38899;
  assign n38822 = n34968 & n38834;
  assign n38823 = n191 ^ n38845;
  assign n38808 = n38852 ^ n38853;
  assign n38847 = ~n38845;
  assign n37684 = n34968 ^ n36394;
  assign n38861 = n38869 & n38870;
  assign n34927 = ~n34968;
  assign n38880 = ~n38888;
  assign n37739 = ~n38822;
  assign n38819 = n34927 & n37708;
  assign n38806 = n38823 ^ n38824;
  assign n38836 = n38808 & n190;
  assign n38842 = n38846 & n38847;
  assign n38835 = ~n38808;
  assign n38778 = n37684 ^ n37617;
  assign n38854 = ~n38861;
  assign n38862 = n38880 & n38881;
  assign n38796 = n38805 ^ n38806;
  assign n38769 = n38806 & n38805;
  assign n37711 = ~n38819;
  assign n38827 = n38835 & n16051;
  assign n38788 = ~n38836;
  assign n38828 = n38778 & n38837;
  assign n38825 = ~n38842;
  assign n38829 = ~n38778;
  assign n38838 = n38854 & n38855;
  assign n38849 = n38862 ^ n36258;
  assign n38863 = ~n38862;
  assign n37661 = ~n38796;
  assign n38807 = n38825 & n38826;
  assign n38810 = ~n38827;
  assign n38780 = ~n38828;
  assign n38820 = n38829 & n38800;
  assign n38815 = n38838 ^ n38839;
  assign n38840 = ~n38838;
  assign n34891 = n38848 ^ n38849;
  assign n38856 = n38863 & n38864;
  assign n38783 = n34891 & n37661;
  assign n38786 = n38807 ^ n38808;
  assign n38772 = n38815 ^ n38816;
  assign n38809 = ~n38807;
  assign n38801 = ~n38820;
  assign n37634 = n34891 ^ n36331;
  assign n38830 = n38840 & n38841;
  assign n34846 = ~n34891;
  assign n38850 = ~n38856;
  assign n37663 = ~n38783;
  assign n38770 = n190 ^ n38786;
  assign n38785 = n34846 & n38796;
  assign n38798 = n38772 & n189;
  assign n38804 = n38809 & n38810;
  assign n38797 = ~n38772;
  assign n38744 = n37634 ^ n37605;
  assign n38817 = ~n38830;
  assign n38831 = n38850 & n38851;
  assign n38759 = n38769 ^ n38770;
  assign n38737 = n38770 & n38769;
  assign n37688 = ~n38785;
  assign n38789 = n38797 & n15951;
  assign n38755 = ~n38798;
  assign n38790 = n38744 & n38763;
  assign n38787 = ~n38804;
  assign n38791 = ~n38744;
  assign n38799 = n38817 & n38818;
  assign n38812 = n38831 ^ n36247;
  assign n38832 = ~n38831;
  assign n37608 = ~n38759;
  assign n38771 = n38787 & n38788;
  assign n38774 = ~n38789;
  assign n38765 = ~n38790;
  assign n38784 = n38791 & n38792;
  assign n38777 = n38799 ^ n38800;
  assign n38802 = ~n38799;
  assign n34757 = n38811 ^ n38812;
  assign n38821 = n38832 & n38833;
  assign n38752 = n34757 & n38759;
  assign n38753 = n38771 ^ n38772;
  assign n38740 = n38777 ^ n38778;
  assign n38773 = ~n38771;
  assign n38746 = ~n38784;
  assign n38793 = n38801 & n38802;
  assign n34824 = ~n34757;
  assign n38813 = ~n38821;
  assign n38749 = n34824 & n37608;
  assign n37639 = ~n38752;
  assign n38738 = n189 ^ n38753;
  assign n38761 = n38740 & n188;
  assign n38768 = n38773 & n38774;
  assign n38760 = ~n38740;
  assign n37586 = n34824 ^ n36247;
  assign n38779 = ~n38793;
  assign n38794 = n38813 & n38814;
  assign n38727 = n38737 ^ n38738;
  assign n38705 = n38738 & n38737;
  assign n37611 = ~n38749;
  assign n38756 = n38760 & n15860;
  assign n38721 = ~n38761;
  assign n38754 = ~n38768;
  assign n38712 = n37586 ^ n37507;
  assign n38762 = n38779 & n38780;
  assign n38776 = n38794 ^ n36120;
  assign n38795 = n38794 & n38803;
  assign n37556 = ~n38727;
  assign n38739 = n38754 & n38755;
  assign n38742 = ~n38756;
  assign n38750 = n38712 & n38757;
  assign n38743 = n38762 ^ n38763;
  assign n38751 = ~n38712;
  assign n38764 = ~n38762;
  assign n34691 = n38775 ^ n38776;
  assign n38781 = ~n38795;
  assign n38716 = n34691 & n37556;
  assign n38719 = n38739 ^ n38740;
  assign n38708 = n38743 ^ n38744;
  assign n38741 = ~n38739;
  assign n38715 = ~n38750;
  assign n38747 = n38751 & n38731;
  assign n37522 = n34691 ^ n36120;
  assign n38758 = n38764 & n38765;
  assign n34733 = ~n34691;
  assign n38766 = n38781 & n38782;
  assign n37558 = ~n38716;
  assign n38706 = n188 ^ n38719;
  assign n38718 = n34733 & n38727;
  assign n38728 = n38708 & n15777;
  assign n38736 = n38741 & n38742;
  assign n38729 = ~n38708;
  assign n38689 = n37522 ^ n37491;
  assign n38733 = ~n38747;
  assign n38745 = ~n38758;
  assign n36190 = n38766 ^ n38767;
  assign n38692 = n38705 ^ n38706;
  assign n38681 = n38706 & n38705;
  assign n37591 = ~n38718;
  assign n38709 = ~n38728;
  assign n38722 = n38729 & n187;
  assign n38725 = n38689 & n38701;
  assign n38720 = ~n38736;
  assign n38723 = ~n38689;
  assign n38730 = n38745 & n38746;
  assign n38735 = n38748 ^ n36190;
  assign n37526 = n38692 ^ n36190;
  assign n38707 = n38720 & n38721;
  assign n38695 = ~n38722;
  assign n38717 = n38723 & n38724;
  assign n38703 = ~n38725;
  assign n38711 = n38730 ^ n38731;
  assign n37493 = n38734 ^ n38735;
  assign n38732 = ~n38730;
  assign n38693 = n38707 ^ n38708;
  assign n38685 = n38711 ^ n38712;
  assign n38671 = n37493 ^ n38713;
  assign n38710 = ~n38707;
  assign n38691 = ~n38717;
  assign n38726 = n38732 & n38733;
  assign n38682 = n187 ^ n38693;
  assign n38699 = n38685 & n186;
  assign n38704 = n38709 & n38710;
  assign n38698 = ~n38685;
  assign n38714 = ~n38726;
  assign n36798 = n38681 ^ n38682;
  assign n38683 = ~n38682;
  assign n38696 = n38698 & n15671;
  assign n38675 = ~n38699;
  assign n38694 = ~n38704;
  assign n38700 = n38714 & n38715;
  assign n38661 = n38672 ^ n36798;
  assign n35914 = n36798 ^ n36790;
  assign n38639 = n36798 & n36790;
  assign n38664 = n38683 & n38681;
  assign n38684 = n38694 & n38695;
  assign n38687 = ~n38696;
  assign n38688 = n38700 ^ n38701;
  assign n38702 = ~n38700;
  assign n37160 = n263 ^ n38661;
  assign n38561 = n38661 & n263;
  assign n38662 = ~n38661;
  assign n38673 = n38684 ^ n38685;
  assign n38667 = n38688 ^ n38689;
  assign n38686 = ~n38684;
  assign n38697 = n38702 & n38703;
  assign n37186 = ~n37160;
  assign n38602 = n38662 & n38663;
  assign n38665 = n186 ^ n38673;
  assign n38677 = n38667 & n15638;
  assign n38680 = n38686 & n38687;
  assign n38678 = ~n38667;
  assign n38690 = ~n38697;
  assign n38659 = n38664 ^ n38665;
  assign n38648 = n38665 & n38664;
  assign n38668 = ~n38677;
  assign n38676 = n38678 & n185;
  assign n38674 = ~n38680;
  assign n38679 = n38690 & n38691;
  assign n38655 = n38659 & n36764;
  assign n38654 = ~n38659;
  assign n38666 = n38674 & n38675;
  assign n38658 = ~n38676;
  assign n38670 = n184 ^ n38679;
  assign n38653 = n38654 & n36621;
  assign n38647 = ~n38655;
  assign n38656 = n38666 ^ n38667;
  assign n38652 = n38670 ^ n38671;
  assign n38669 = ~n38666;
  assign n38646 = n38647 & n38639;
  assign n38645 = ~n38653;
  assign n38649 = n185 ^ n38656;
  assign n38660 = n38668 & n38669;
  assign n38644 = ~n38646;
  assign n38638 = n38647 & n38645;
  assign n38627 = n38648 ^ n38649;
  assign n38650 = ~n38649;
  assign n38657 = ~n38660;
  assign n35729 = n38638 ^ n38639;
  assign n38636 = n38644 & n38645;
  assign n38641 = n38627 & n36590;
  assign n38640 = ~n38627;
  assign n38642 = n38650 & n38648;
  assign n38651 = n38657 & n38658;
  assign n38625 = n38631 ^ n35729;
  assign n38628 = n38636 ^ n36588;
  assign n35891 = ~n35729;
  assign n38633 = ~n38636;
  assign n38637 = n38640 & n36588;
  assign n38624 = ~n38641;
  assign n38643 = n38651 ^ n38652;
  assign n38622 = n38625 & n38626;
  assign n35700 = n38627 ^ n38628;
  assign n38620 = ~n38625;
  assign n38632 = ~n38637;
  assign n38605 = n38642 ^ n38643;
  assign n38573 = n38618 ^ n35700;
  assign n38619 = n38620 & n38621;
  assign n38604 = ~n38622;
  assign n35722 = ~n35700;
  assign n38629 = n38632 & n38633;
  assign n38634 = n38605 & n36526;
  assign n38635 = ~n38605;
  assign n38609 = n38573 & n38611;
  assign n38610 = ~n38573;
  assign n38614 = ~n38619;
  assign n38623 = ~n38629;
  assign n38608 = ~n38634;
  assign n38630 = n38635 & n36491;
  assign n38591 = ~n38609;
  assign n38600 = n38610 & n38589;
  assign n38612 = n38614 & n38602;
  assign n38601 = n38614 & n38604;
  assign n38615 = n38623 & n38624;
  assign n38617 = ~n38630;
  assign n38577 = ~n38600;
  assign n38598 = n38601 ^ n38602;
  assign n38603 = ~n38612;
  assign n38606 = n38615 ^ n36491;
  assign n38616 = ~n38615;
  assign n38593 = n38598 & n262;
  assign n38592 = ~n38598;
  assign n38599 = n38603 & n38604;
  assign n35635 = n38605 ^ n38606;
  assign n38613 = n38616 & n38617;
  assign n38587 = n38592 & n11627;
  assign n38567 = ~n38593;
  assign n38543 = n38594 ^ n35635;
  assign n38588 = ~n38599;
  assign n35619 = ~n35635;
  assign n38607 = ~n38613;
  assign n38580 = n38543 & n38585;
  assign n38578 = ~n38587;
  assign n38579 = ~n38543;
  assign n38572 = n38588 ^ n38589;
  assign n38586 = n38591 & n38588;
  assign n38595 = n38607 & n38608;
  assign n38539 = n38572 ^ n38573;
  assign n38574 = n38578 & n38561;
  assign n38560 = n38578 & n38567;
  assign n38575 = n38579 & n38563;
  assign n38547 = ~n38580;
  assign n38576 = ~n38586;
  assign n38581 = n38595 ^ n36420;
  assign n38596 = ~n38595;
  assign n38555 = n38539 & n11492;
  assign n38544 = n38560 ^ n38561;
  assign n38556 = ~n38539;
  assign n38566 = ~n38574;
  assign n38564 = ~n38575;
  assign n38562 = n38576 & n38577;
  assign n35548 = n38581 ^ n38582;
  assign n38590 = n38596 & n38597;
  assign n37137 = n38544 ^ n37160;
  assign n38505 = n38544 & n37160;
  assign n38545 = ~n38555;
  assign n38553 = n38556 & n261;
  assign n38542 = n38562 ^ n38563;
  assign n38558 = n38566 & n38567;
  assign n38513 = n38568 ^ n35548;
  assign n38565 = ~n38562;
  assign n35561 = ~n35548;
  assign n38583 = ~n38590;
  assign n38292 = ~n37137;
  assign n38515 = n38542 ^ n38543;
  assign n38549 = n38513 & n38552;
  assign n38530 = ~n38553;
  assign n38538 = ~n38558;
  assign n38548 = ~n38513;
  assign n38557 = n38564 & n38565;
  assign n38571 = n38583 & n38584;
  assign n38528 = n38515 & n260;
  assign n38527 = ~n38515;
  assign n38523 = n38538 ^ n38539;
  assign n38537 = n38545 & n38538;
  assign n38540 = n38548 & n38532;
  assign n38517 = ~n38549;
  assign n38546 = ~n38557;
  assign n38570 = n38571 & n36346;
  assign n38569 = ~n38571;
  assign n38506 = n261 ^ n38523;
  assign n38522 = n38527 & n11437;
  assign n38496 = ~n38528;
  assign n38529 = ~n38537;
  assign n38534 = ~n38540;
  assign n38531 = n38546 & n38547;
  assign n38559 = n38569 & n36402;
  assign n38551 = ~n38570;
  assign n37104 = n38505 ^ n38506;
  assign n38508 = ~n38506;
  assign n38510 = ~n38522;
  assign n38514 = n38529 & n38530;
  assign n38512 = n38531 ^ n38532;
  assign n38533 = ~n38531;
  assign n38550 = n38551 & n38554;
  assign n38536 = ~n38559;
  assign n38253 = ~n37104;
  assign n38475 = n38508 & n38505;
  assign n38479 = n38512 ^ n38513;
  assign n38494 = n38514 ^ n38515;
  assign n38511 = ~n38514;
  assign n38524 = n38533 & n38534;
  assign n38535 = ~n38550;
  assign n38541 = n38536 & n38551;
  assign n38476 = n260 ^ n38494;
  assign n38498 = n38479 & n259;
  assign n38497 = ~n38479;
  assign n38507 = n38510 & n38511;
  assign n38516 = ~n38524;
  assign n38519 = n38535 & n38536;
  assign n38526 = ~n38541;
  assign n37086 = n38475 ^ n38476;
  assign n38477 = ~n38476;
  assign n38490 = n38497 & n11347;
  assign n38460 = ~n38498;
  assign n38495 = ~n38507;
  assign n38499 = n38516 & n38517;
  assign n38501 = n38519 ^ n36309;
  assign n35515 = n38525 ^ n38526;
  assign n38520 = ~n38519;
  assign n38213 = ~n37086;
  assign n38441 = n38477 & n38475;
  assign n38480 = ~n38490;
  assign n38478 = n38495 & n38496;
  assign n38482 = n38499 ^ n38500;
  assign n35419 = n38501 ^ n38502;
  assign n38474 = ~n38499;
  assign n38483 = n38509 ^ n35515;
  assign n38518 = n38520 & n38521;
  assign n35455 = ~n35515;
  assign n38458 = n38478 ^ n38479;
  assign n38445 = n38482 ^ n38483;
  assign n38420 = n38485 ^ n35419;
  assign n38481 = ~n38478;
  assign n38491 = n38483 & n38500;
  assign n35383 = ~n35419;
  assign n38492 = ~n38483;
  assign n38503 = ~n38518;
  assign n38442 = n259 ^ n38458;
  assign n38461 = n38445 & n11226;
  assign n38462 = ~n38445;
  assign n38466 = n38420 & n38435;
  assign n38472 = n38480 & n38481;
  assign n38464 = ~n38420;
  assign n38457 = ~n38491;
  assign n38486 = n38492 & n38493;
  assign n38487 = n38503 & n38504;
  assign n37037 = n38441 ^ n38442;
  assign n38443 = ~n38442;
  assign n38446 = ~n38461;
  assign n38455 = n38462 & n258;
  assign n38463 = n38464 & n38465;
  assign n38425 = ~n38466;
  assign n38459 = ~n38472;
  assign n38473 = ~n38486;
  assign n38467 = n38487 ^ n36201;
  assign n38488 = ~n38487;
  assign n38175 = ~n37037;
  assign n38415 = n38443 & n38441;
  assign n38428 = ~n38455;
  assign n38444 = n38459 & n38460;
  assign n38440 = ~n38463;
  assign n35365 = n38467 ^ n38468;
  assign n38469 = n38473 & n38474;
  assign n38484 = n38488 & n38489;
  assign n38426 = n38444 ^ n38445;
  assign n38394 = n38449 ^ n35365;
  assign n38447 = ~n38444;
  assign n35307 = ~n35365;
  assign n38456 = ~n38469;
  assign n38470 = ~n38484;
  assign n38416 = n258 ^ n38426;
  assign n38431 = n38394 & n38439;
  assign n38438 = n38446 & n38447;
  assign n38430 = ~n38394;
  assign n38450 = n38456 & n38457;
  assign n38451 = n38470 & n38471;
  assign n38136 = n38415 ^ n38416;
  assign n38364 = n38416 & n38415;
  assign n38429 = n38430 & n38412;
  assign n38396 = ~n38431;
  assign n38427 = ~n38438;
  assign n38434 = ~n38450;
  assign n38433 = n38451 ^ n38452;
  assign n38453 = ~n38451;
  assign n38128 = ~n38136;
  assign n38399 = n38427 & n38428;
  assign n38414 = ~n38429;
  assign n35217 = n36167 ^ n38433;
  assign n38419 = n38434 ^ n38435;
  assign n38432 = n38440 & n38434;
  assign n38448 = n38453 & n38454;
  assign n38359 = n38418 ^ n35217;
  assign n38400 = n38419 ^ n38420;
  assign n38388 = ~n38399;
  assign n35257 = ~n35217;
  assign n38424 = ~n38432;
  assign n38436 = ~n38448;
  assign n38386 = n38399 ^ n38400;
  assign n38404 = n38359 & n38381;
  assign n38405 = n38400 & n257;
  assign n38402 = ~n38359;
  assign n38401 = ~n38400;
  assign n38411 = n38424 & n38425;
  assign n38421 = n38436 & n38437;
  assign n38365 = n257 ^ n38386;
  assign n38397 = n38401 & n11154;
  assign n38398 = n38402 & n38403;
  assign n38361 = ~n38404;
  assign n38369 = ~n38405;
  assign n38393 = n38411 ^ n38412;
  assign n38413 = ~n38411;
  assign n38408 = n38421 ^ n36105;
  assign n38422 = ~n38421;
  assign n36994 = n38364 ^ n38365;
  assign n38366 = ~n38365;
  assign n38351 = n38393 ^ n38394;
  assign n38387 = ~n38397;
  assign n38383 = ~n38398;
  assign n35140 = n38407 ^ n38408;
  assign n38406 = n38413 & n38414;
  assign n38417 = n38422 & n38423;
  assign n38094 = ~n36994;
  assign n38312 = n38366 & n38364;
  assign n38379 = n38351 & n256;
  assign n38378 = ~n38351;
  assign n38384 = n38387 & n38388;
  assign n38327 = n38389 ^ n35140;
  assign n35180 = ~n35140;
  assign n38395 = ~n38406;
  assign n38409 = ~n38417;
  assign n38315 = ~n38312;
  assign n38367 = n38378 & n11085;
  assign n38333 = ~n38379;
  assign n38372 = n38327 & n38346;
  assign n38368 = ~n38384;
  assign n38370 = ~n38327;
  assign n38380 = n38395 & n38396;
  assign n38390 = n38409 & n38410;
  assign n38353 = ~n38367;
  assign n38362 = n38368 & n38369;
  assign n38363 = n38370 & n38371;
  assign n38347 = ~n38372;
  assign n38358 = n38380 ^ n38381;
  assign n38382 = ~n38380;
  assign n38375 = n38390 ^ n36047;
  assign n38391 = ~n38390;
  assign n38319 = n38358 ^ n38359;
  assign n38350 = ~n38362;
  assign n38329 = ~n38363;
  assign n35099 = n38374 ^ n38375;
  assign n38373 = n38382 & n38383;
  assign n38385 = n38391 & n38392;
  assign n38342 = n38319 & n10976;
  assign n38330 = n38350 ^ n38351;
  assign n38349 = n38353 & n38350;
  assign n38343 = ~n38319;
  assign n38289 = n38354 ^ n35099;
  assign n35052 = ~n35099;
  assign n38360 = ~n38373;
  assign n38376 = ~n38385;
  assign n38313 = n256 ^ n38330;
  assign n38320 = ~n38342;
  assign n38334 = n38343 & n271;
  assign n38336 = n38289 & n38344;
  assign n38332 = ~n38349;
  assign n38335 = ~n38289;
  assign n38345 = n38360 & n38361;
  assign n38355 = n38376 & n38377;
  assign n36935 = n38312 ^ n38313;
  assign n38314 = ~n38313;
  assign n38318 = n38332 & n38333;
  assign n38296 = ~n38334;
  assign n38331 = n38335 & n38309;
  assign n38291 = ~n38336;
  assign n38326 = n38345 ^ n38346;
  assign n38348 = ~n38345;
  assign n38338 = n38355 ^ n35994;
  assign n38356 = ~n38355;
  assign n38056 = ~n36935;
  assign n38276 = n38314 & n38315;
  assign n38294 = n38318 ^ n38319;
  assign n38279 = n38326 ^ n38327;
  assign n38321 = ~n38318;
  assign n38311 = ~n38331;
  assign n34998 = n38338 ^ n38339;
  assign n38337 = n38347 & n38348;
  assign n38352 = n38356 & n38357;
  assign n38277 = n271 ^ n38294;
  assign n38287 = ~n38276;
  assign n38306 = n38279 & n10896;
  assign n38316 = n38320 & n38321;
  assign n38307 = ~n38279;
  assign n38250 = n38322 ^ n34998;
  assign n34977 = ~n34998;
  assign n38328 = ~n38337;
  assign n38340 = ~n38352;
  assign n36917 = n38276 ^ n38277;
  assign n38236 = n38277 & n38287;
  assign n38280 = ~n38306;
  assign n38297 = n38307 & n270;
  assign n38300 = n38250 & n38270;
  assign n38295 = ~n38316;
  assign n38298 = ~n38250;
  assign n38308 = n38328 & n38329;
  assign n38323 = n38340 & n38341;
  assign n38018 = ~n36917;
  assign n38239 = ~n38236;
  assign n38278 = n38295 & n38296;
  assign n38257 = ~n38297;
  assign n38293 = n38298 & n38299;
  assign n38252 = ~n38300;
  assign n38288 = n38308 ^ n38309;
  assign n38310 = ~n38308;
  assign n38302 = n38323 ^ n35927;
  assign n38324 = ~n38323;
  assign n38255 = n38278 ^ n38279;
  assign n38241 = n38288 ^ n38289;
  assign n38281 = ~n38278;
  assign n38272 = ~n38293;
  assign n34902 = n38302 ^ n38303;
  assign n38301 = n38310 & n38311;
  assign n38317 = n38324 & n38325;
  assign n38237 = n270 ^ n38255;
  assign n38268 = n38241 & n269;
  assign n38273 = n38280 & n38281;
  assign n38267 = ~n38241;
  assign n38210 = n38282 ^ n34902;
  assign n38283 = n34902 & n38292;
  assign n34950 = ~n34902;
  assign n38290 = ~n38301;
  assign n38304 = ~n38317;
  assign n37972 = n38236 ^ n38237;
  assign n38238 = ~n38237;
  assign n38258 = n38267 & n10806;
  assign n38217 = ~n38268;
  assign n38259 = n38210 & n38230;
  assign n38256 = ~n38273;
  assign n38260 = ~n38210;
  assign n38274 = n34950 & n37137;
  assign n37152 = ~n38283;
  assign n38269 = n38290 & n38291;
  assign n38284 = n38304 & n38305;
  assign n36860 = ~n37972;
  assign n38198 = n38238 & n38239;
  assign n38240 = n38256 & n38257;
  assign n38243 = ~n38258;
  assign n38232 = ~n38259;
  assign n38254 = n38260 & n38261;
  assign n38249 = n38269 ^ n38270;
  assign n37139 = ~n38274;
  assign n38271 = ~n38269;
  assign n38263 = n38284 ^ n35883;
  assign n38285 = ~n38284;
  assign n38215 = n38240 ^ n38241;
  assign n38201 = n38249 ^ n38250;
  assign n38242 = ~n38240;
  assign n38212 = ~n38254;
  assign n34863 = n38263 ^ n38264;
  assign n38262 = n38271 & n38272;
  assign n38275 = n38285 & n38286;
  assign n38199 = n269 ^ n38215;
  assign n38226 = n38201 & n10723;
  assign n38233 = n38242 & n38243;
  assign n38227 = ~n38201;
  assign n38172 = n38244 ^ n34863;
  assign n38245 = n34863 & n38253;
  assign n34820 = ~n34863;
  assign n38251 = ~n38262;
  assign n38265 = ~n38275;
  assign n36825 = n38198 ^ n38199;
  assign n38159 = n38199 & n38198;
  assign n38202 = ~n38226;
  assign n38218 = n38227 & n268;
  assign n38219 = n38172 & n38228;
  assign n38216 = ~n38233;
  assign n38220 = ~n38172;
  assign n38234 = n34820 & n37104;
  assign n37106 = ~n38245;
  assign n38229 = n38251 & n38252;
  assign n38246 = n38265 & n38266;
  assign n37942 = ~n36825;
  assign n38170 = ~n38159;
  assign n38200 = n38216 & n38217;
  assign n38179 = ~n38218;
  assign n38174 = ~n38219;
  assign n38214 = n38220 & n38192;
  assign n38209 = n38229 ^ n38230;
  assign n37120 = ~n38234;
  assign n38231 = ~n38229;
  assign n38222 = n38246 ^ n35838;
  assign n38247 = ~n38246;
  assign n38177 = n38200 ^ n38201;
  assign n38162 = n38209 ^ n38210;
  assign n38203 = ~n38200;
  assign n38194 = ~n38214;
  assign n34724 = n38222 ^ n38223;
  assign n38221 = n38231 & n38232;
  assign n38235 = n38247 & n38248;
  assign n38160 = n268 ^ n38177;
  assign n38188 = n38162 & n10627;
  assign n38195 = n38202 & n38203;
  assign n38189 = ~n38162;
  assign n38133 = n38204 ^ n34724;
  assign n38205 = n34724 & n38213;
  assign n34749 = ~n34724;
  assign n38211 = ~n38221;
  assign n38224 = ~n38235;
  assign n36786 = n38159 ^ n38160;
  assign n38118 = n38160 & n38170;
  assign n38164 = ~n38188;
  assign n38180 = n38189 & n267;
  assign n38181 = n38133 & n38190;
  assign n38178 = ~n38195;
  assign n38182 = ~n38133;
  assign n38196 = n34749 & n37086;
  assign n37071 = ~n38205;
  assign n38191 = n38211 & n38212;
  assign n38206 = n38224 & n38225;
  assign n37902 = ~n36786;
  assign n38121 = ~n38118;
  assign n38161 = n38178 & n38179;
  assign n38140 = ~n38180;
  assign n38135 = ~n38181;
  assign n38176 = n38182 & n38153;
  assign n38171 = n38191 ^ n38192;
  assign n37088 = ~n38196;
  assign n38193 = ~n38191;
  assign n38185 = n38206 ^ n35790;
  assign n38207 = ~n38206;
  assign n38138 = n38161 ^ n38162;
  assign n38123 = n38171 ^ n38172;
  assign n38163 = ~n38161;
  assign n38155 = ~n38176;
  assign n34697 = n38184 ^ n38185;
  assign n38183 = n38193 & n38194;
  assign n38197 = n38207 & n38208;
  assign n38119 = n267 ^ n38138;
  assign n38150 = n38123 & n266;
  assign n38156 = n38163 & n38164;
  assign n38149 = ~n38123;
  assign n38091 = n34697 ^ n38165;
  assign n38166 = n34697 & n38175;
  assign n34647 = ~n34697;
  assign n38173 = ~n38183;
  assign n38186 = ~n38197;
  assign n36737 = n38118 ^ n38119;
  assign n38120 = ~n38119;
  assign n38141 = n38149 & n10589;
  assign n38099 = ~n38150;
  assign n38142 = n38091 & n38151;
  assign n38139 = ~n38156;
  assign n38143 = ~n38091;
  assign n38157 = n34647 & n37037;
  assign n37039 = ~n38166;
  assign n38152 = n38173 & n38174;
  assign n38167 = n38186 & n38187;
  assign n37864 = ~n36737;
  assign n38079 = n38120 & n38121;
  assign n38122 = n38139 & n38140;
  assign n38125 = ~n38141;
  assign n38093 = ~n38142;
  assign n38137 = n38143 & n38112;
  assign n38132 = n38152 ^ n38153;
  assign n37058 = ~n38157;
  assign n38154 = ~n38152;
  assign n38145 = n38167 ^ n35795;
  assign n38168 = ~n38167;
  assign n38097 = n38122 ^ n38123;
  assign n38082 = n38132 ^ n38133;
  assign n38124 = ~n38122;
  assign n38114 = ~n38137;
  assign n34663 = n38145 ^ n38146;
  assign n38144 = n38154 & n38155;
  assign n38158 = n38168 & n38169;
  assign n38080 = n266 ^ n38097;
  assign n38109 = n38082 & n265;
  assign n38115 = n38124 & n38125;
  assign n38108 = ~n38082;
  assign n38053 = n38126 ^ n34663;
  assign n38127 = n34663 & n38136;
  assign n34589 = ~n34663;
  assign n38134 = ~n38144;
  assign n38147 = ~n38158;
  assign n37818 = n38079 ^ n38080;
  assign n38042 = n38080 & n38079;
  assign n38100 = n38108 & n10522;
  assign n38060 = ~n38109;
  assign n38102 = n38053 & n38110;
  assign n38098 = ~n38115;
  assign n38101 = ~n38053;
  assign n37011 = ~n38127;
  assign n38116 = n34589 & n38128;
  assign n38111 = n38134 & n38135;
  assign n38129 = n38147 & n38148;
  assign n37826 = ~n37818;
  assign n38081 = n38098 & n38099;
  assign n38084 = ~n38100;
  assign n38095 = n38101 & n38073;
  assign n38055 = ~n38102;
  assign n38090 = n38111 ^ n38112;
  assign n37027 = ~n38116;
  assign n38113 = ~n38111;
  assign n38105 = n38129 ^ n35648;
  assign n38130 = ~n38129;
  assign n38058 = n38081 ^ n38082;
  assign n38021 = n38090 ^ n38091;
  assign n38083 = ~n38081;
  assign n38075 = ~n38095;
  assign n38096 = n37011 & n37027;
  assign n34525 = n38104 ^ n38105;
  assign n38103 = n38113 & n38114;
  assign n38117 = n38130 & n38131;
  assign n38043 = n265 ^ n38058;
  assign n38070 = n38021 & n264;
  assign n38076 = n38083 & n38084;
  assign n38069 = ~n38021;
  assign n38036 = n38085 ^ n34525;
  assign n38086 = n34525 & n38094;
  assign n37025 = ~n38096;
  assign n34619 = ~n34525;
  assign n38092 = ~n38103;
  assign n38106 = ~n38117;
  assign n37785 = n38042 ^ n38043;
  assign n38004 = n38043 & n38042;
  assign n38061 = n38069 & n10470;
  assign n38023 = ~n38070;
  assign n38063 = n38036 & n38071;
  assign n38059 = ~n38076;
  assign n38062 = ~n38036;
  assign n36973 = ~n38086;
  assign n38077 = n34619 & n36994;
  assign n38072 = n38092 & n38093;
  assign n38087 = n38106 & n38107;
  assign n36664 = ~n37785;
  assign n38044 = n38059 & n38060;
  assign n38046 = ~n38061;
  assign n38057 = n38062 & n38015;
  assign n38038 = ~n38063;
  assign n38052 = n38072 ^ n38073;
  assign n36996 = ~n38077;
  assign n38074 = ~n38072;
  assign n38066 = n38087 ^ n35574;
  assign n38088 = ~n38087;
  assign n38020 = n264 ^ n38044;
  assign n37983 = n38052 ^ n38053;
  assign n38045 = ~n38044;
  assign n38017 = ~n38057;
  assign n34489 = n38065 ^ n38066;
  assign n38064 = n38074 & n38075;
  assign n38078 = n38088 & n38089;
  assign n38005 = n38020 ^ n38021;
  assign n38034 = n37983 & n279;
  assign n38039 = n38045 & n38046;
  assign n38033 = ~n37983;
  assign n37998 = n38047 ^ n34489;
  assign n38048 = n34489 & n38056;
  assign n34536 = ~n34489;
  assign n38054 = ~n38064;
  assign n38067 = ~n38078;
  assign n37736 = n38004 ^ n38005;
  assign n37965 = n38005 & n38004;
  assign n38024 = n38033 & n10418;
  assign n37985 = ~n38034;
  assign n38027 = n37998 & n37978;
  assign n38022 = ~n38039;
  assign n38025 = ~n37998;
  assign n38040 = n34536 & n36935;
  assign n36938 = ~n38048;
  assign n38035 = n38054 & n38055;
  assign n38049 = n38067 & n38068;
  assign n36571 = ~n37736;
  assign n38006 = n38022 & n38023;
  assign n38008 = ~n38024;
  assign n38019 = n38025 & n38026;
  assign n37980 = ~n38027;
  assign n38014 = n38035 ^ n38036;
  assign n36956 = ~n38040;
  assign n38037 = ~n38035;
  assign n38030 = n38049 ^ n35538;
  assign n38050 = ~n38049;
  assign n37982 = n279 ^ n38006;
  assign n37968 = n38014 ^ n38015;
  assign n38007 = ~n38006;
  assign n38000 = ~n38019;
  assign n34462 = n38029 ^ n38030;
  assign n38028 = n38037 & n38038;
  assign n38041 = n38050 & n38051;
  assign n37966 = n37982 ^ n37983;
  assign n37996 = n37968 & n278;
  assign n38001 = n38007 & n38008;
  assign n37995 = ~n37968;
  assign n37939 = n38009 ^ n34462;
  assign n38010 = n34462 & n38018;
  assign n34474 = ~n34462;
  assign n38016 = ~n38028;
  assign n38031 = ~n38041;
  assign n36505 = n37965 ^ n37966;
  assign n37924 = n37966 & n37965;
  assign n37986 = n37995 & n10398;
  assign n37946 = ~n37996;
  assign n37987 = n37939 & n37959;
  assign n37984 = ~n38001;
  assign n37988 = ~n37939;
  assign n38002 = n34474 & n36917;
  assign n36902 = ~n38010;
  assign n37997 = n38016 & n38017;
  assign n38011 = n38031 & n38032;
  assign n37693 = ~n36505;
  assign n37927 = ~n37924;
  assign n37967 = n37984 & n37985;
  assign n37970 = ~n37986;
  assign n37961 = ~n37987;
  assign n37981 = n37988 & n37989;
  assign n37977 = n37997 ^ n37998;
  assign n36919 = ~n38002;
  assign n37999 = ~n37997;
  assign n37992 = n38011 ^ n35469;
  assign n38012 = ~n38011;
  assign n37944 = n37967 ^ n37968;
  assign n37929 = n37977 ^ n37978;
  assign n37969 = ~n37967;
  assign n37941 = ~n37981;
  assign n34419 = n37991 ^ n37992;
  assign n37990 = n37999 & n38000;
  assign n38003 = n38012 & n38013;
  assign n37925 = n278 ^ n37944;
  assign n37956 = n37929 & n10372;
  assign n37962 = n37969 & n37970;
  assign n37957 = ~n37929;
  assign n37899 = n37971 ^ n34419;
  assign n37973 = n34419 & n36860;
  assign n34434 = ~n34419;
  assign n37979 = ~n37990;
  assign n37993 = ~n38003;
  assign n36435 = n37924 ^ n37925;
  assign n37926 = ~n37925;
  assign n37931 = ~n37956;
  assign n37947 = n37957 & n277;
  assign n37950 = n37899 & n37918;
  assign n37945 = ~n37962;
  assign n37948 = ~n37899;
  assign n37963 = n34434 & n37972;
  assign n36862 = ~n37973;
  assign n37958 = n37979 & n37980;
  assign n37974 = n37993 & n37994;
  assign n37636 = ~n36435;
  assign n37887 = n37926 & n37927;
  assign n37928 = n37945 & n37946;
  assign n37906 = ~n37947;
  assign n37943 = n37948 & n37949;
  assign n37920 = ~n37950;
  assign n37938 = n37958 ^ n37959;
  assign n36885 = ~n37963;
  assign n37960 = ~n37958;
  assign n37953 = n37974 ^ n35434;
  assign n37975 = ~n37974;
  assign n37904 = n37928 ^ n37929;
  assign n37890 = n37938 ^ n37939;
  assign n37930 = ~n37928;
  assign n37901 = ~n37943;
  assign n34409 = n37952 ^ n37953;
  assign n37951 = n37960 & n37961;
  assign n37964 = n37975 & n37976;
  assign n37888 = n277 ^ n37904;
  assign n37915 = n37890 & n10334;
  assign n37921 = n37930 & n37931;
  assign n37916 = ~n37890;
  assign n37861 = n37932 ^ n34409;
  assign n37933 = n34409 & n37942;
  assign n34379 = ~n34409;
  assign n37940 = ~n37951;
  assign n37954 = ~n37964;
  assign n36360 = n37887 ^ n37888;
  assign n37849 = n37888 & n37887;
  assign n37891 = ~n37915;
  assign n37907 = n37916 & n276;
  assign n37910 = n37861 & n37881;
  assign n37905 = ~n37921;
  assign n37908 = ~n37861;
  assign n36828 = ~n37933;
  assign n37922 = n34379 & n36825;
  assign n37917 = n37940 & n37941;
  assign n37934 = n37954 & n37955;
  assign n37588 = ~n36360;
  assign n37889 = n37905 & n37906;
  assign n37868 = ~n37907;
  assign n37903 = n37908 & n37909;
  assign n37883 = ~n37910;
  assign n37898 = n37917 ^ n37918;
  assign n36845 = ~n37922;
  assign n37919 = ~n37917;
  assign n37912 = n37934 ^ n37935;
  assign n37936 = ~n37934;
  assign n37866 = n37889 ^ n37890;
  assign n37852 = n37898 ^ n37899;
  assign n37892 = ~n37889;
  assign n37863 = ~n37903;
  assign n34345 = n35359 ^ n37912;
  assign n37911 = n37919 & n37920;
  assign n37923 = n37936 & n37937;
  assign n37850 = n276 ^ n37866;
  assign n37877 = n37852 & n10269;
  assign n37884 = n37891 & n37892;
  assign n37878 = ~n37852;
  assign n37823 = n37893 ^ n34345;
  assign n37894 = n34345 & n37902;
  assign n34368 = ~n34345;
  assign n37900 = ~n37911;
  assign n37913 = ~n37923;
  assign n36287 = n37849 ^ n37850;
  assign n37808 = n37850 & n37849;
  assign n37854 = ~n37877;
  assign n37869 = n37878 & n275;
  assign n37870 = n37823 & n37879;
  assign n37867 = ~n37884;
  assign n37871 = ~n37823;
  assign n37885 = n34368 & n36786;
  assign n36788 = ~n37894;
  assign n37880 = n37900 & n37901;
  assign n37895 = n37913 & n37914;
  assign n37524 = ~n36287;
  assign n37811 = ~n37808;
  assign n37851 = n37867 & n37868;
  assign n37830 = ~n37869;
  assign n37825 = ~n37870;
  assign n37865 = n37871 & n37843;
  assign n37860 = n37880 ^ n37881;
  assign n36809 = ~n37885;
  assign n37882 = ~n37880;
  assign n37873 = n37895 ^ n35239;
  assign n37896 = ~n37895;
  assign n37828 = n37851 ^ n37852;
  assign n37813 = n37860 ^ n37861;
  assign n37853 = ~n37851;
  assign n37845 = ~n37865;
  assign n34311 = n37873 ^ n37874;
  assign n37872 = n37882 & n37883;
  assign n37886 = n37896 & n37897;
  assign n37809 = n275 ^ n37828;
  assign n37839 = n37813 & n10216;
  assign n37846 = n37853 & n37854;
  assign n37840 = ~n37813;
  assign n37782 = n37855 ^ n34311;
  assign n37856 = n34311 & n37864;
  assign n34333 = ~n34311;
  assign n37862 = ~n37872;
  assign n37875 = ~n37886;
  assign n37494 = n37808 ^ n37809;
  assign n37810 = ~n37809;
  assign n37814 = ~n37839;
  assign n37831 = n37840 & n274;
  assign n37833 = n37782 & n37841;
  assign n37829 = ~n37846;
  assign n37832 = ~n37782;
  assign n37847 = n34333 & n36737;
  assign n36740 = ~n37856;
  assign n37842 = n37862 & n37863;
  assign n37857 = n37875 & n37876;
  assign n37769 = n37810 & n37811;
  assign n37812 = n37829 & n37830;
  assign n37789 = ~n37831;
  assign n37827 = n37832 & n37802;
  assign n37784 = ~n37833;
  assign n37822 = n37842 ^ n37843;
  assign n36762 = ~n37847;
  assign n37844 = ~n37842;
  assign n37835 = n37857 ^ n35213;
  assign n37858 = ~n37857;
  assign n37787 = n37812 ^ n37813;
  assign n37773 = n37822 ^ n37823;
  assign n37815 = ~n37812;
  assign n37804 = ~n37827;
  assign n34253 = n37835 ^ n37836;
  assign n37834 = n37844 & n37845;
  assign n37848 = n37858 & n37859;
  assign n37770 = n274 ^ n37787;
  assign n37800 = n37773 & n273;
  assign n37805 = n37814 & n37815;
  assign n37799 = ~n37773;
  assign n37743 = n37816 ^ n34253;
  assign n37817 = n34253 & n37826;
  assign n34303 = ~n34253;
  assign n37824 = ~n37834;
  assign n37837 = ~n37848;
  assign n35920 = n37769 ^ n37770;
  assign n37771 = ~n37770;
  assign n37790 = n37799 & n10199;
  assign n37750 = ~n37800;
  assign n37793 = n37743 & n37763;
  assign n37788 = ~n37805;
  assign n37791 = ~n37743;
  assign n36691 = ~n37817;
  assign n37806 = n34303 & n37818;
  assign n37801 = n37824 & n37825;
  assign n37819 = n37837 & n37838;
  assign n37740 = n36790 ^ n35920;
  assign n37728 = n35920 ^ n37747;
  assign n34029 = n35914 ^ n35920;
  assign n37648 = n35920 & n35914;
  assign n37729 = n37771 & n37769;
  assign n37772 = n37788 & n37789;
  assign n37775 = ~n37790;
  assign n37786 = n37791 & n37792;
  assign n37745 = ~n37793;
  assign n37781 = n37801 ^ n37802;
  assign n36718 = ~n37806;
  assign n37803 = ~n37801;
  assign n37796 = n37819 ^ n35040;
  assign n37820 = ~n37819;
  assign n37016 = n359 ^ n37728;
  assign n37574 = n37740 & n37741;
  assign n37512 = n37728 & n359;
  assign n37748 = n37772 ^ n37773;
  assign n37701 = n37781 ^ n37782;
  assign n37774 = ~n37772;
  assign n37765 = ~n37786;
  assign n36715 = n36691 & n36718;
  assign n34216 = n37795 ^ n37796;
  assign n37794 = n37803 & n37804;
  assign n37807 = n37820 & n37821;
  assign n37715 = n37574 & n37542;
  assign n37716 = n37512 & n358;
  assign n37009 = ~n37016;
  assign n37713 = ~n37574;
  assign n37712 = ~n37512;
  assign n37730 = n273 ^ n37748;
  assign n37760 = n37701 & n272;
  assign n37766 = n37774 & n37775;
  assign n37759 = ~n37701;
  assign n37722 = n37776 ^ n34216;
  assign n37777 = n34216 & n37785;
  assign n34296 = ~n34216;
  assign n37783 = ~n37794;
  assign n37797 = ~n37807;
  assign n37696 = n37712 & n4928;
  assign n37697 = n37713 & n37714;
  assign n37560 = ~n37715;
  assign n37496 = ~n37716;
  assign n37717 = n37729 ^ n37730;
  assign n37677 = n37730 & n37729;
  assign n37751 = n37759 & n10140;
  assign n37703 = ~n37760;
  assign n37753 = n37722 & n37761;
  assign n37749 = ~n37766;
  assign n37752 = ~n37722;
  assign n37767 = n34296 & n36664;
  assign n36666 = ~n37777;
  assign n37762 = n37783 & n37784;
  assign n37778 = n37797 & n37798;
  assign n37527 = ~n37696;
  assign n37592 = ~n37697;
  assign n37698 = n37717 & n35891;
  assign n37699 = ~n37717;
  assign n37680 = ~n37677;
  assign n37731 = n37749 & n37750;
  assign n37733 = ~n37751;
  assign n37746 = n37752 & n37690;
  assign n37724 = ~n37753;
  assign n37742 = n37762 ^ n37763;
  assign n36636 = ~n37767;
  assign n37764 = ~n37762;
  assign n37756 = n37778 ^ n34964;
  assign n37779 = ~n37778;
  assign n37676 = ~n37698;
  assign n37694 = n37699 & n35729;
  assign n37700 = n272 ^ n37731;
  assign n37652 = n37742 ^ n37743;
  assign n37732 = ~n37731;
  assign n37692 = ~n37746;
  assign n34174 = n37755 ^ n37756;
  assign n37754 = n37764 & n37765;
  assign n37768 = n37779 & n37780;
  assign n37675 = n37676 & n37648;
  assign n37665 = ~n37694;
  assign n37678 = n37700 ^ n37701;
  assign n37718 = n37652 & n10097;
  assign n37725 = n37732 & n37733;
  assign n37719 = ~n37652;
  assign n37669 = n37734 ^ n34174;
  assign n37735 = n34174 & n36571;
  assign n34221 = ~n34174;
  assign n37744 = ~n37754;
  assign n37757 = ~n37768;
  assign n37664 = ~n37675;
  assign n37647 = n37665 & n37676;
  assign n37613 = n37677 ^ n37678;
  assign n37679 = ~n37678;
  assign n37683 = ~n37718;
  assign n37704 = n37719 & n287;
  assign n37705 = n37669 & n37720;
  assign n37702 = ~n37725;
  assign n37706 = ~n37669;
  assign n36574 = ~n37735;
  assign n37726 = n34221 & n37736;
  assign n37721 = n37744 & n37745;
  assign n37737 = n37757 & n37758;
  assign n33982 = n37647 ^ n37648;
  assign n37640 = n37664 & n37665;
  assign n37649 = n37613 & n35700;
  assign n37650 = ~n37613;
  assign n37626 = n37679 & n37680;
  assign n37681 = n37702 & n37703;
  assign n37654 = ~n37704;
  assign n37671 = ~n37705;
  assign n37695 = n37706 & n37642;
  assign n37689 = n37721 ^ n37722;
  assign n36608 = ~n37726;
  assign n37723 = ~n37721;
  assign n37709 = n37737 ^ n34968;
  assign n37738 = ~n37737;
  assign n36678 = n33982 ^ n35729;
  assign n37612 = n37640 ^ n35722;
  assign n33978 = ~n33982;
  assign n37624 = ~n37640;
  assign n37599 = ~n37649;
  assign n37645 = n37650 & n35722;
  assign n37629 = ~n37626;
  assign n37651 = n287 ^ n37681;
  assign n37631 = n37689 ^ n37690;
  assign n37682 = ~n37681;
  assign n37644 = ~n37695;
  assign n34181 = n37708 ^ n37709;
  assign n37707 = n37723 & n37724;
  assign n37727 = n37738 & n37739;
  assign n37575 = n36678 ^ n36621;
  assign n33929 = n37612 ^ n37613;
  assign n37625 = ~n37645;
  assign n37627 = n37651 ^ n37652;
  assign n37667 = n37631 & n286;
  assign n37672 = n37682 & n37683;
  assign n37666 = ~n37631;
  assign n37594 = n37684 ^ n34181;
  assign n37685 = n34181 & n37693;
  assign n34157 = ~n34181;
  assign n37691 = ~n37707;
  assign n37710 = ~n37727;
  assign n37541 = n37574 ^ n37575;
  assign n37576 = n37575 & n37592;
  assign n36622 = n33929 ^ n35700;
  assign n33967 = ~n33929;
  assign n37620 = n37624 & n37625;
  assign n37544 = n37626 ^ n37627;
  assign n37628 = ~n37627;
  assign n37655 = n37666 & n10065;
  assign n37602 = ~n37667;
  assign n37658 = n37594 & n37617;
  assign n37653 = ~n37672;
  assign n37656 = ~n37594;
  assign n36507 = ~n37685;
  assign n37673 = n34157 & n36505;
  assign n37668 = n37691 & n37692;
  assign n37686 = n37710 & n37711;
  assign n37513 = n37541 ^ n37542;
  assign n37497 = n36622 ^ n36590;
  assign n37559 = ~n37576;
  assign n37598 = ~n37620;
  assign n37562 = ~n37544;
  assign n37580 = n37628 & n37629;
  assign n37630 = n37653 & n37654;
  assign n37633 = ~n37655;
  assign n37646 = n37656 & n37657;
  assign n37619 = ~n37658;
  assign n37641 = n37668 ^ n37669;
  assign n36542 = ~n37673;
  assign n37670 = ~n37668;
  assign n37660 = n37686 ^ n34846;
  assign n37687 = ~n37686;
  assign n37480 = n37512 ^ n37513;
  assign n37514 = n37513 & n37527;
  assign n37528 = n37497 & n37532;
  assign n37529 = ~n37497;
  assign n37531 = n37559 & n37560;
  assign n37577 = n37598 & n37599;
  assign n37600 = n37630 ^ n37631;
  assign n37583 = n37641 ^ n37642;
  assign n37632 = ~n37630;
  assign n37596 = ~n37646;
  assign n34125 = n37660 ^ n37661;
  assign n37659 = n37670 & n37671;
  assign n37674 = n37687 & n37688;
  assign n35797 = n358 ^ n37480;
  assign n37495 = ~n37514;
  assign n37468 = ~n37528;
  assign n37515 = n37529 & n37530;
  assign n37498 = n37531 ^ n37532;
  assign n37500 = ~n37531;
  assign n37543 = n37577 ^ n35619;
  assign n37579 = n37577 & n35619;
  assign n37578 = ~n37577;
  assign n37581 = n286 ^ n37600;
  assign n37615 = n37583 & n285;
  assign n37621 = n37632 & n37633;
  assign n37614 = ~n37583;
  assign n37536 = n37634 ^ n34125;
  assign n37635 = n34125 & n36435;
  assign n34185 = ~n34125;
  assign n37643 = ~n37659;
  assign n37662 = ~n37674;
  assign n36964 = ~n35797;
  assign n37463 = n37495 & n37496;
  assign n37464 = n37497 ^ n37498;
  assign n37499 = ~n37515;
  assign n33917 = n37543 ^ n37544;
  assign n37570 = n37578 & n35635;
  assign n37561 = ~n37579;
  assign n37563 = n37580 ^ n37581;
  assign n37516 = n37581 & n37580;
  assign n37603 = n37614 & n10044;
  assign n37549 = ~n37615;
  assign n37606 = n37536 & n37567;
  assign n37601 = ~n37621;
  assign n37604 = ~n37536;
  assign n36437 = ~n37635;
  assign n37622 = n34185 & n37636;
  assign n37616 = n37643 & n37644;
  assign n37637 = n37662 & n37663;
  assign n37434 = n37463 ^ n37464;
  assign n37465 = n37464 & n4867;
  assign n37450 = ~n37463;
  assign n37466 = ~n37464;
  assign n37481 = n37499 & n37500;
  assign n36559 = n35635 ^ n33917;
  assign n33941 = ~n33917;
  assign n37545 = n37561 & n37562;
  assign n37546 = n37563 & n35561;
  assign n37534 = ~n37570;
  assign n37470 = ~n37563;
  assign n37582 = n37601 & n37602;
  assign n37585 = ~n37603;
  assign n37597 = n37604 & n37605;
  assign n37538 = ~n37606;
  assign n37593 = n37616 ^ n37617;
  assign n36473 = ~n37622;
  assign n37618 = ~n37616;
  assign n37609 = n37637 ^ n34757;
  assign n37638 = ~n37637;
  assign n37409 = n357 ^ n37434;
  assign n37449 = ~n37465;
  assign n37453 = n37466 & n357;
  assign n37467 = ~n37481;
  assign n37410 = n36559 ^ n36526;
  assign n37533 = ~n37545;
  assign n37539 = n37470 & n35548;
  assign n37503 = ~n37546;
  assign n37547 = n37582 ^ n37583;
  assign n37519 = n37593 ^ n37594;
  assign n37584 = ~n37582;
  assign n37569 = ~n37597;
  assign n34107 = n37608 ^ n37609;
  assign n37607 = n37618 & n37619;
  assign n37623 = n37638 & n37639;
  assign n35747 = n37409 ^ n35797;
  assign n37343 = n37409 & n35797;
  assign n37435 = n37449 & n37450;
  assign n37423 = ~n37453;
  assign n37436 = n37467 & n37468;
  assign n37456 = n37410 & n37437;
  assign n37454 = ~n37410;
  assign n37501 = n37533 & n37534;
  assign n37472 = ~n37539;
  assign n37517 = n285 ^ n37547;
  assign n37564 = n37519 & n9976;
  assign n37571 = n37584 & n37585;
  assign n37565 = ~n37519;
  assign n37475 = n34107 ^ n37586;
  assign n37587 = n34107 & n36360;
  assign n34087 = ~n34107;
  assign n37595 = ~n37607;
  assign n37610 = ~n37623;
  assign n36914 = ~n35747;
  assign n37422 = ~n37435;
  assign n37411 = n37436 ^ n37437;
  assign n37439 = ~n37436;
  assign n37451 = n37454 & n37455;
  assign n37438 = ~n37456;
  assign n37469 = n37501 ^ n35561;
  assign n37502 = ~n37501;
  assign n37414 = n37516 ^ n37517;
  assign n37457 = n37517 & n37516;
  assign n37521 = ~n37564;
  assign n37550 = n37565 & n284;
  assign n37551 = n37475 & n37507;
  assign n37548 = ~n37571;
  assign n37552 = ~n37475;
  assign n36362 = ~n37587;
  assign n37572 = n34087 & n37588;
  assign n37566 = n37595 & n37596;
  assign n37589 = n37610 & n37611;
  assign n37389 = n37410 ^ n37411;
  assign n37388 = n37422 & n37423;
  assign n37425 = n37438 & n37439;
  assign n37413 = ~n37451;
  assign n33910 = n37469 ^ n37470;
  assign n37482 = n37502 & n37503;
  assign n37483 = n37414 & n35455;
  assign n37484 = ~n37414;
  assign n37473 = ~n37457;
  assign n37518 = n37548 & n37549;
  assign n37487 = ~n37550;
  assign n37477 = ~n37551;
  assign n37540 = n37552 & n37553;
  assign n37535 = n37566 ^ n37567;
  assign n36399 = ~n37572;
  assign n37568 = ~n37566;
  assign n37555 = n37589 ^ n34733;
  assign n37590 = ~n37589;
  assign n37365 = n37388 ^ n37389;
  assign n37390 = n37389 & n4824;
  assign n37391 = ~n37389;
  assign n37376 = ~n37388;
  assign n37412 = ~n37425;
  assign n36494 = n33910 ^ n35548;
  assign n33886 = ~n33910;
  assign n37471 = ~n37482;
  assign n37442 = ~n37483;
  assign n37478 = n37484 & n35515;
  assign n37485 = n37518 ^ n37519;
  assign n37460 = n37535 ^ n37536;
  assign n37520 = ~n37518;
  assign n37509 = ~n37540;
  assign n34116 = n37555 ^ n37556;
  assign n37554 = n37568 & n37569;
  assign n37573 = n37590 & n37591;
  assign n37344 = n356 ^ n37365;
  assign n37375 = ~n37390;
  assign n37378 = n37391 & n356;
  assign n37402 = n37412 & n37413;
  assign n37357 = n36494 ^ n36474;
  assign n37440 = n37471 & n37472;
  assign n37417 = ~n37478;
  assign n37458 = n284 ^ n37485;
  assign n37504 = n37460 & n9936;
  assign n37510 = n37520 & n37521;
  assign n37505 = ~n37460;
  assign n37419 = n34116 ^ n37522;
  assign n37523 = n34116 & n36287;
  assign n34057 = ~n34116;
  assign n37537 = ~n37554;
  assign n37557 = ~n37573;
  assign n35654 = n37343 ^ n37344;
  assign n37290 = n37344 & n37343;
  assign n37366 = n37375 & n37376;
  assign n37353 = ~n37378;
  assign n37392 = n37357 & n37379;
  assign n37368 = ~n37402;
  assign n37393 = ~n37357;
  assign n37415 = n37440 ^ n35515;
  assign n37441 = ~n37440;
  assign n37370 = n37457 ^ n37458;
  assign n37403 = n37458 & n37473;
  assign n37462 = ~n37504;
  assign n37488 = n37505 & n283;
  assign n37489 = n37419 & n37446;
  assign n37486 = ~n37510;
  assign n37490 = ~n37419;
  assign n36336 = ~n37523;
  assign n37511 = n34057 & n37524;
  assign n37506 = n37537 & n37538;
  assign n37525 = n37557 & n37558;
  assign n36893 = ~n35654;
  assign n37352 = ~n37366;
  assign n37356 = n37368 ^ n37379;
  assign n37346 = ~n37392;
  assign n37380 = n37393 & n37394;
  assign n33853 = n37414 ^ n37415;
  assign n37426 = n37441 & n37442;
  assign n37427 = n37370 & n35383;
  assign n37428 = ~n37370;
  assign n37459 = n37486 & n37487;
  assign n37431 = ~n37488;
  assign n37421 = ~n37489;
  assign n37479 = n37490 & n37491;
  assign n37474 = n37506 ^ n37507;
  assign n36295 = ~n37511;
  assign n37508 = ~n37506;
  assign n34060 = n37525 ^ n37526;
  assign n37330 = n37352 & n37353;
  assign n37331 = n37356 ^ n37357;
  assign n37367 = ~n37380;
  assign n36423 = n33853 ^ n35515;
  assign n33871 = ~n33853;
  assign n37416 = ~n37426;
  assign n37397 = ~n37427;
  assign n37424 = n37428 & n35419;
  assign n37429 = n37459 ^ n37460;
  assign n37406 = n37474 ^ n37475;
  assign n37461 = ~n37459;
  assign n37448 = ~n37479;
  assign n37374 = n37493 ^ n34060;
  assign n36263 = n37494 ^ n34060;
  assign n37492 = n37508 & n37509;
  assign n37313 = n37330 ^ n37331;
  assign n37316 = ~n37330;
  assign n37335 = n37331 & n355;
  assign n37334 = ~n37331;
  assign n37358 = n37367 & n37368;
  assign n37306 = n36423 ^ n36402;
  assign n37395 = n37416 & n37417;
  assign n37372 = ~n37424;
  assign n37404 = n283 ^ n37429;
  assign n37443 = n37406 & n9908;
  assign n37452 = n37461 & n37462;
  assign n37444 = ~n37406;
  assign n37476 = ~n37492;
  assign n37291 = n355 ^ n37313;
  assign n37332 = n37334 & n4762;
  assign n37297 = ~n37335;
  assign n37347 = n37306 & n37354;
  assign n37345 = ~n37358;
  assign n37348 = ~n37306;
  assign n37369 = n37395 ^ n35383;
  assign n37396 = ~n37395;
  assign n37327 = n37403 ^ n37404;
  assign n37359 = n37404 & n37403;
  assign n37408 = ~n37443;
  assign n37432 = n37444 & n282;
  assign n37430 = ~n37452;
  assign n37445 = n37476 & n37477;
  assign n35615 = n37290 ^ n37291;
  assign n37292 = ~n37291;
  assign n37315 = ~n37332;
  assign n37322 = n37345 & n37346;
  assign n37308 = ~n37347;
  assign n37336 = n37348 & n37323;
  assign n33816 = n37369 ^ n37370;
  assign n37381 = n37396 & n37397;
  assign n37383 = n37327 & n35365;
  assign n37382 = ~n37327;
  assign n37405 = n37430 & n37431;
  assign n37386 = ~n37432;
  assign n37418 = n37445 ^ n37446;
  assign n37447 = ~n37445;
  assign n36852 = ~n35615;
  assign n37240 = n37292 & n37290;
  assign n37314 = n37315 & n37316;
  assign n37305 = n37322 ^ n37323;
  assign n37324 = ~n37322;
  assign n37325 = ~n37336;
  assign n33820 = ~n33816;
  assign n37371 = ~n37381;
  assign n37377 = n37382 & n35307;
  assign n37329 = ~n37383;
  assign n37384 = n37405 ^ n37406;
  assign n37362 = n37418 ^ n37419;
  assign n37407 = ~n37405;
  assign n37433 = n37447 & n37448;
  assign n37243 = ~n37240;
  assign n37274 = n37305 ^ n37306;
  assign n37296 = ~n37314;
  assign n37317 = n37324 & n37325;
  assign n36349 = n33820 ^ n35419;
  assign n37349 = n37371 & n37372;
  assign n37351 = ~n37377;
  assign n37360 = n282 ^ n37384;
  assign n37398 = n37362 & n9894;
  assign n37401 = n37407 & n37408;
  assign n37399 = ~n37362;
  assign n37420 = ~n37433;
  assign n37283 = n37274 & n354;
  assign n37293 = n37296 & n37297;
  assign n37282 = ~n37274;
  assign n37307 = ~n37317;
  assign n37267 = n36349 ^ n36273;
  assign n37326 = n37349 ^ n35307;
  assign n37350 = ~n37349;
  assign n37287 = n37359 ^ n37360;
  assign n37318 = n37360 & n37359;
  assign n37364 = ~n37398;
  assign n37387 = n37399 & n281;
  assign n37385 = ~n37401;
  assign n37400 = n37420 & n37421;
  assign n37277 = n37282 & n4727;
  assign n37251 = ~n37283;
  assign n37265 = ~n37293;
  assign n37284 = n37307 & n37308;
  assign n37299 = n37267 & n37309;
  assign n37298 = ~n37267;
  assign n33754 = n37326 ^ n37327;
  assign n37337 = n37350 & n37351;
  assign n37339 = n37287 & n35217;
  assign n37338 = ~n37287;
  assign n37361 = n37385 & n37386;
  assign n37342 = ~n37387;
  assign n37373 = n280 ^ n37400;
  assign n37258 = n37265 ^ n37274;
  assign n37264 = ~n37277;
  assign n37266 = n37284 ^ n37285;
  assign n37278 = ~n37284;
  assign n37294 = n37298 & n37285;
  assign n37261 = ~n37299;
  assign n36276 = n35365 ^ n33754;
  assign n33799 = ~n33754;
  assign n37328 = ~n37337;
  assign n37333 = n37338 & n35257;
  assign n37289 = ~n37339;
  assign n37340 = n37361 ^ n37362;
  assign n37321 = n37373 ^ n37374;
  assign n37363 = ~n37361;
  assign n37241 = n354 ^ n37258;
  assign n37259 = n37264 & n37265;
  assign n37231 = n37266 ^ n37267;
  assign n37225 = n36276 ^ n36254;
  assign n37279 = ~n37294;
  assign n37310 = n37328 & n37329;
  assign n37312 = ~n37333;
  assign n37319 = n281 ^ n37340;
  assign n37355 = n37363 & n37364;
  assign n35509 = n37240 ^ n37241;
  assign n37242 = ~n37241;
  assign n37253 = n37231 & n353;
  assign n37250 = ~n37259;
  assign n37252 = ~n37231;
  assign n37268 = n37225 & n37247;
  assign n37275 = n37278 & n37279;
  assign n37269 = ~n37225;
  assign n37286 = n37310 ^ n35257;
  assign n37311 = ~n37310;
  assign n37254 = n37318 ^ n37319;
  assign n37303 = n37319 & n37318;
  assign n37341 = ~n37355;
  assign n36817 = ~n35509;
  assign n37194 = n37242 & n37243;
  assign n37230 = n37250 & n37251;
  assign n37245 = n37252 & n4683;
  assign n37218 = ~n37253;
  assign n37227 = ~n37268;
  assign n37262 = n37269 & n37270;
  assign n37260 = ~n37275;
  assign n33765 = n37286 ^ n37287;
  assign n37300 = n37311 & n37312;
  assign n37302 = n37254 & n35180;
  assign n37301 = ~n37254;
  assign n37320 = n37341 & n37342;
  assign n37197 = ~n37194;
  assign n37216 = n37230 ^ n37231;
  assign n37232 = ~n37230;
  assign n37233 = ~n37245;
  assign n37246 = n37260 & n37261;
  assign n37249 = ~n37262;
  assign n36204 = n33765 ^ n35257;
  assign n33732 = ~n33765;
  assign n37288 = ~n37300;
  assign n37295 = n37301 & n35140;
  assign n37257 = ~n37302;
  assign n37304 = n37320 ^ n37321;
  assign n37195 = n353 ^ n37216;
  assign n37223 = n37232 & n37233;
  assign n37224 = n37246 ^ n37247;
  assign n37188 = n36204 ^ n36133;
  assign n37248 = ~n37246;
  assign n37271 = n37288 & n37289;
  assign n37273 = ~n37295;
  assign n37220 = n37303 ^ n37304;
  assign n35436 = n37194 ^ n37195;
  assign n37196 = ~n37195;
  assign n37217 = ~n37223;
  assign n37199 = n37224 ^ n37225;
  assign n37234 = n37188 & n37213;
  assign n37244 = n37248 & n37249;
  assign n37235 = ~n37188;
  assign n37255 = n37271 ^ n35140;
  assign n37272 = ~n37271;
  assign n37280 = n37220 & n35099;
  assign n37281 = ~n37220;
  assign n36774 = ~n35436;
  assign n37161 = n37196 & n37197;
  assign n37198 = n37217 & n37218;
  assign n37210 = n37199 & n4635;
  assign n37211 = ~n37199;
  assign n37191 = ~n37234;
  assign n37228 = n37235 & n37236;
  assign n37226 = ~n37244;
  assign n33730 = n37254 ^ n37255;
  assign n37263 = n37272 & n37273;
  assign n37222 = ~n37280;
  assign n37276 = n37281 & n35052;
  assign n37181 = n37198 ^ n37199;
  assign n37201 = ~n37198;
  assign n37200 = ~n37210;
  assign n37207 = n37211 & n352;
  assign n37212 = n37226 & n37227;
  assign n37215 = ~n37228;
  assign n36136 = n33730 ^ n35180;
  assign n33697 = ~n33730;
  assign n37256 = ~n37263;
  assign n37239 = ~n37276;
  assign n37162 = n352 ^ n37181;
  assign n37187 = n37200 & n37201;
  assign n37183 = ~n37207;
  assign n37189 = n37212 ^ n37213;
  assign n37155 = n36136 ^ n36071;
  assign n37214 = ~n37212;
  assign n37237 = n37256 & n37257;
  assign n35362 = n37161 ^ n37162;
  assign n37126 = n37162 & n37161;
  assign n37182 = ~n37187;
  assign n37164 = n37188 ^ n37189;
  assign n37204 = n37155 & n37177;
  assign n37208 = n37214 & n37215;
  assign n37202 = ~n37155;
  assign n37219 = n37237 ^ n35052;
  assign n37238 = ~n37237;
  assign n36714 = ~n35362;
  assign n37129 = ~n37126;
  assign n37163 = n37182 & n37183;
  assign n37174 = n37164 & n4592;
  assign n37175 = ~n37164;
  assign n37192 = n37202 & n37203;
  assign n37179 = ~n37204;
  assign n37190 = ~n37208;
  assign n33695 = n37219 ^ n37220;
  assign n37229 = n37238 & n37239;
  assign n37146 = n37163 ^ n37164;
  assign n37165 = ~n37163;
  assign n37166 = ~n37174;
  assign n37170 = n37175 & n367;
  assign n37176 = n37190 & n37191;
  assign n37157 = ~n37192;
  assign n36074 = n35099 ^ n33695;
  assign n33661 = ~n33695;
  assign n37221 = ~n37229;
  assign n37127 = n367 ^ n37146;
  assign n37153 = n37165 & n37166;
  assign n37148 = ~n37170;
  assign n37154 = n37176 ^ n37177;
  assign n37123 = n36074 ^ n36047;
  assign n37178 = ~n37176;
  assign n37209 = n37221 & n37222;
  assign n35283 = n37126 ^ n37127;
  assign n37128 = ~n37127;
  assign n37147 = ~n37153;
  assign n37131 = n37154 ^ n37155;
  assign n37169 = n37123 & n37143;
  assign n37171 = n37178 & n37179;
  assign n37167 = ~n37123;
  assign n37206 = n37209 & n34977;
  assign n37205 = ~n37209;
  assign n36688 = ~n35283;
  assign n37094 = n37128 & n37129;
  assign n37130 = n37147 & n37148;
  assign n37140 = n37131 & n4556;
  assign n37141 = ~n37131;
  assign n37158 = n37167 & n37168;
  assign n37125 = ~n37169;
  assign n37156 = ~n37171;
  assign n37193 = n37205 & n34998;
  assign n37185 = ~n37206;
  assign n37100 = ~n37094;
  assign n37114 = n37130 ^ n37131;
  assign n37132 = ~n37130;
  assign n37133 = ~n37140;
  assign n37134 = n37141 & n366;
  assign n37142 = n37156 & n37157;
  assign n37145 = ~n37158;
  assign n37184 = n37185 & n37186;
  assign n37173 = ~n37193;
  assign n37095 = n366 ^ n37114;
  assign n37121 = n37132 & n37133;
  assign n37116 = ~n37134;
  assign n37122 = n37142 ^ n37143;
  assign n37144 = ~n37142;
  assign n37172 = ~n37184;
  assign n37180 = n37173 & n37185;
  assign n35246 = n37094 ^ n37095;
  assign n37062 = n37095 & n37100;
  assign n37115 = ~n37121;
  assign n37097 = n37122 ^ n37123;
  assign n37135 = n37144 & n37145;
  assign n37150 = n37172 & n37173;
  assign n37159 = ~n37180;
  assign n36616 = ~n35246;
  assign n37096 = n37115 & n37116;
  assign n37107 = n37097 & n4506;
  assign n37108 = ~n37097;
  assign n37124 = ~n37135;
  assign n37136 = n37150 ^ n34902;
  assign n33659 = n37159 ^ n37160;
  assign n37151 = ~n37150;
  assign n37076 = n37096 ^ n37097;
  assign n37098 = ~n37096;
  assign n37099 = ~n37107;
  assign n37101 = n37108 & n365;
  assign n37109 = n37124 & n37125;
  assign n33621 = n37136 ^ n37137;
  assign n36017 = n34998 ^ n33659;
  assign n37149 = n37151 & n37152;
  assign n33623 = ~n33659;
  assign n37063 = n365 ^ n37076;
  assign n37089 = n37098 & n37099;
  assign n37078 = ~n37101;
  assign n37090 = n37109 ^ n37110;
  assign n37093 = ~n37109;
  assign n35972 = n34950 ^ n33621;
  assign n37091 = n36017 ^ n35969;
  assign n33585 = ~n33621;
  assign n37138 = ~n37149;
  assign n35124 = n37062 ^ n37063;
  assign n37032 = n37063 & n37062;
  assign n37077 = ~n37089;
  assign n37065 = n37090 ^ n37091;
  assign n37035 = n35972 ^ n35959;
  assign n37111 = n37091 & n37110;
  assign n37112 = ~n37091;
  assign n37118 = n37138 & n37139;
  assign n36549 = ~n35124;
  assign n37064 = n37077 & n37078;
  assign n37072 = n37065 & n4471;
  assign n37073 = ~n37065;
  assign n37081 = n37035 & n37053;
  assign n37082 = ~n37035;
  assign n37075 = ~n37111;
  assign n37102 = n37112 & n37113;
  assign n37103 = n37118 ^ n34820;
  assign n37119 = ~n37118;
  assign n37043 = n37064 ^ n37065;
  assign n37066 = ~n37064;
  assign n37067 = ~n37072;
  assign n37068 = n37073 & n364;
  assign n37041 = ~n37081;
  assign n37079 = n37082 & n37083;
  assign n37092 = ~n37102;
  assign n33547 = n37103 ^ n37104;
  assign n37117 = n37119 & n37120;
  assign n37033 = n364 ^ n37043;
  assign n37059 = n37066 & n37067;
  assign n37045 = ~n37068;
  assign n37060 = ~n37079;
  assign n37084 = n37092 & n37093;
  assign n33572 = ~n33547;
  assign n37105 = ~n37117;
  assign n35046 = n37032 ^ n37033;
  assign n36983 = n37033 & n37032;
  assign n37044 = ~n37059;
  assign n35930 = n34863 ^ n33572;
  assign n37074 = ~n37084;
  assign n37085 = n37105 & n37106;
  assign n36481 = ~n35046;
  assign n37019 = n37044 & n37045;
  assign n37013 = n35930 ^ n35915;
  assign n37069 = n37074 & n37075;
  assign n35886 = n37085 ^ n37086;
  assign n37087 = ~n37085;
  assign n37007 = ~n37019;
  assign n37047 = n37013 & n37050;
  assign n37046 = ~n37013;
  assign n37052 = ~n37069;
  assign n36975 = n35869 ^ n35886;
  assign n33507 = n35886 ^ n34749;
  assign n37080 = n37087 & n37088;
  assign n37042 = n37046 & n37029;
  assign n37015 = ~n37047;
  assign n37034 = n37052 ^ n37053;
  assign n37051 = n37060 & n37052;
  assign n37055 = n36975 & n37061;
  assign n37054 = ~n36975;
  assign n33534 = ~n33507;
  assign n37070 = ~n37080;
  assign n37020 = n37034 ^ n37035;
  assign n37031 = ~n37042;
  assign n37040 = ~n37051;
  assign n37048 = n37054 & n37000;
  assign n36977 = ~n37055;
  assign n37056 = n37070 & n37071;
  assign n37005 = n37019 ^ n37020;
  assign n37022 = n37020 & n363;
  assign n37021 = ~n37020;
  assign n37028 = n37040 & n37041;
  assign n37002 = ~n37048;
  assign n37036 = n37056 ^ n34647;
  assign n37057 = ~n37056;
  assign n36984 = n363 ^ n37005;
  assign n37017 = n37021 & n4427;
  assign n36988 = ~n37022;
  assign n37012 = n37028 ^ n37029;
  assign n37030 = ~n37028;
  assign n33463 = n37036 ^ n37037;
  assign n37049 = n37057 & n37058;
  assign n34971 = n36983 ^ n36984;
  assign n36985 = ~n36984;
  assign n36967 = n37012 ^ n37013;
  assign n37006 = ~n37017;
  assign n35841 = n34697 ^ n33463;
  assign n37023 = n37030 & n37031;
  assign n33505 = ~n33463;
  assign n37038 = ~n37049;
  assign n36410 = ~n34971;
  assign n36926 = n36985 & n36983;
  assign n36998 = n36967 & n362;
  assign n36997 = ~n36967;
  assign n37003 = n37006 & n37007;
  assign n36939 = n35841 ^ n35818;
  assign n37014 = ~n37023;
  assign n37024 = n37038 & n37039;
  assign n36929 = ~n36926;
  assign n36986 = n36997 & n4376;
  assign n36948 = ~n36998;
  assign n36989 = n36939 & n36960;
  assign n36987 = ~n37003;
  assign n36990 = ~n36939;
  assign n36999 = n37014 & n37015;
  assign n33410 = n37024 ^ n37025;
  assign n37026 = ~n37024;
  assign n36969 = ~n36986;
  assign n36979 = n36987 & n36988;
  assign n36962 = ~n36989;
  assign n36980 = n36990 & n36991;
  assign n36974 = n36999 ^ n37000;
  assign n37001 = ~n36999;
  assign n35820 = n33410 ^ n34663;
  assign n37008 = n33410 & n37016;
  assign n33488 = ~n33410;
  assign n37018 = n37026 & n37027;
  assign n36932 = n36974 ^ n36975;
  assign n36966 = ~n36979;
  assign n36942 = ~n36980;
  assign n36923 = n35820 ^ n35795;
  assign n36992 = n37001 & n37002;
  assign n35822 = ~n37008;
  assign n37004 = n33488 & n37009;
  assign n37010 = ~n37018;
  assign n36958 = n36932 & n361;
  assign n36943 = n36966 ^ n36967;
  assign n36965 = n36969 & n36966;
  assign n36957 = ~n36932;
  assign n36971 = n36923 & n36978;
  assign n36970 = ~n36923;
  assign n36976 = ~n36992;
  assign n35845 = ~n37004;
  assign n36993 = n37010 & n37011;
  assign n36927 = n362 ^ n36943;
  assign n36949 = n36957 & n4334;
  assign n36911 = ~n36958;
  assign n36947 = ~n36965;
  assign n36968 = n36970 & n36904;
  assign n36925 = ~n36971;
  assign n36959 = n36976 & n36977;
  assign n36981 = n35845 & n35822;
  assign n35726 = n36993 ^ n36994;
  assign n36995 = ~n36993;
  assign n36324 = n36926 ^ n36927;
  assign n36928 = ~n36927;
  assign n36931 = n36947 & n36948;
  assign n36933 = ~n36949;
  assign n36940 = n36959 ^ n36960;
  assign n36906 = ~n36968;
  assign n36961 = ~n36959;
  assign n36889 = n35726 ^ n35717;
  assign n33371 = n34525 ^ n35726;
  assign n35843 = ~n36981;
  assign n36982 = n36995 & n36996;
  assign n34893 = ~n36324;
  assign n36895 = n36928 & n36929;
  assign n36909 = n36931 ^ n36932;
  assign n36898 = n36939 ^ n36940;
  assign n36934 = ~n36931;
  assign n36950 = n36961 & n36962;
  assign n36951 = n36889 & n36963;
  assign n36953 = n33371 & n36964;
  assign n36952 = ~n36889;
  assign n33418 = ~n33371;
  assign n36972 = ~n36982;
  assign n36896 = n361 ^ n36909;
  assign n36920 = n36898 & n4295;
  assign n36930 = n36933 & n36934;
  assign n36921 = ~n36898;
  assign n36941 = ~n36950;
  assign n36891 = ~n36951;
  assign n36944 = n36952 & n36865;
  assign n36945 = n33418 & n35797;
  assign n35772 = ~n36953;
  assign n36954 = n36972 & n36973;
  assign n34808 = n36895 ^ n36896;
  assign n36854 = n36896 & n36895;
  assign n36900 = ~n36920;
  assign n36912 = n36921 & n360;
  assign n36910 = ~n36930;
  assign n36922 = n36941 & n36942;
  assign n36867 = ~n36944;
  assign n35799 = ~n36945;
  assign n36936 = n36954 ^ n34489;
  assign n36955 = ~n36954;
  assign n36261 = ~n34808;
  assign n36863 = ~n36854;
  assign n36897 = n36910 & n36911;
  assign n36874 = ~n36912;
  assign n36903 = n36922 ^ n36923;
  assign n36924 = ~n36922;
  assign n33332 = n36935 ^ n36936;
  assign n36946 = n36955 & n36956;
  assign n36872 = n36897 ^ n36898;
  assign n36837 = n36903 ^ n36904;
  assign n36899 = ~n36897;
  assign n35684 = n33332 ^ n34489;
  assign n36913 = n36924 & n36925;
  assign n36915 = n33332 & n35747;
  assign n33388 = ~n33332;
  assign n36937 = ~n36946;
  assign n36855 = n360 ^ n36872;
  assign n36887 = n36837 & n375;
  assign n36894 = n36899 & n36900;
  assign n36886 = ~n36837;
  assign n36849 = n35653 ^ n35684;
  assign n36905 = ~n36913;
  assign n36907 = n33388 & n36914;
  assign n35720 = ~n36915;
  assign n36916 = n36937 & n36938;
  assign n34735 = n36854 ^ n36855;
  assign n36819 = n36855 & n36863;
  assign n36875 = n36886 & n4257;
  assign n36839 = ~n36887;
  assign n36878 = n36849 & n36831;
  assign n36873 = ~n36894;
  assign n36876 = ~n36849;
  assign n36888 = n36905 & n36906;
  assign n35749 = ~n36907;
  assign n35613 = n36916 ^ n36917;
  assign n36918 = ~n36916;
  assign n36829 = ~n36819;
  assign n36856 = n36873 & n36874;
  assign n36858 = ~n36875;
  assign n36868 = n36876 & n36877;
  assign n36833 = ~n36878;
  assign n36864 = n36888 ^ n36889;
  assign n36890 = ~n36888;
  assign n36792 = n35613 ^ n35586;
  assign n33312 = n35613 ^ n34474;
  assign n36908 = n36918 & n36919;
  assign n36836 = n375 ^ n36856;
  assign n36822 = n36864 ^ n36865;
  assign n36857 = ~n36856;
  assign n36851 = ~n36868;
  assign n36879 = n36890 & n36891;
  assign n36880 = n36792 & n36892;
  assign n36882 = n33312 & n36893;
  assign n36881 = ~n36792;
  assign n33351 = ~n33312;
  assign n36901 = ~n36908;
  assign n36820 = n36836 ^ n36837;
  assign n36847 = n36822 & n374;
  assign n36853 = n36857 & n36858;
  assign n36846 = ~n36822;
  assign n36866 = ~n36879;
  assign n36794 = ~n36880;
  assign n36869 = n36881 & n36814;
  assign n35687 = ~n36882;
  assign n36870 = n33351 & n35654;
  assign n36883 = n36901 & n36902;
  assign n34031 = n36819 ^ n36820;
  assign n36777 = n36820 & n36829;
  assign n36840 = n36846 & n4218;
  assign n36801 = ~n36847;
  assign n36838 = ~n36853;
  assign n36848 = n36866 & n36867;
  assign n36816 = ~n36869;
  assign n35657 = ~n36870;
  assign n36859 = n36883 ^ n34434;
  assign n36884 = ~n36883;
  assign n36789 = n35914 ^ n34031;
  assign n36776 = n36798 ^ n34031;
  assign n33088 = n34029 ^ n34031;
  assign n36701 = n34031 & n34029;
  assign n36780 = ~n36777;
  assign n36821 = n36838 & n36839;
  assign n36823 = ~n36840;
  assign n36830 = n36848 ^ n36849;
  assign n36850 = ~n36848;
  assign n33272 = n36859 ^ n36860;
  assign n36871 = n36884 & n36885;
  assign n34386 = n455 ^ n36776;
  assign n36647 = n36789 & n36790;
  assign n36518 = n36776 & n455;
  assign n36799 = n36821 ^ n36822;
  assign n36782 = n36830 ^ n36831;
  assign n36824 = ~n36821;
  assign n35541 = n34419 ^ n33272;
  assign n36841 = n36850 & n36851;
  assign n36842 = n33272 & n36852;
  assign n33300 = ~n33272;
  assign n36861 = ~n36871;
  assign n36765 = n36647 & n36621;
  assign n35323 = ~n34386;
  assign n36763 = ~n36647;
  assign n36778 = n374 ^ n36799;
  assign n36810 = n36782 & n4169;
  assign n36818 = n36823 & n36824;
  assign n36811 = ~n36782;
  assign n36742 = n35541 ^ n35516;
  assign n36832 = ~n36841;
  assign n36834 = n33300 & n35615;
  assign n35581 = ~n36842;
  assign n36843 = n36861 & n36862;
  assign n36749 = n36763 & n36764;
  assign n36638 = ~n36765;
  assign n36766 = n36777 ^ n36778;
  assign n36779 = ~n36778;
  assign n36784 = ~n36810;
  assign n36802 = n36811 & n373;
  assign n36803 = n36742 & n36812;
  assign n36800 = ~n36818;
  assign n36804 = ~n36742;
  assign n36813 = n36832 & n36833;
  assign n35617 = ~n36834;
  assign n36826 = n36843 ^ n34409;
  assign n36844 = ~n36843;
  assign n36667 = ~n36749;
  assign n36750 = n36766 & n33982;
  assign n36751 = ~n36766;
  assign n36729 = n36779 & n36780;
  assign n36781 = n36800 & n36801;
  assign n36754 = ~n36802;
  assign n36744 = ~n36803;
  assign n36795 = n36804 & n36771;
  assign n36791 = n36813 ^ n36814;
  assign n36815 = ~n36813;
  assign n33270 = n36825 ^ n36826;
  assign n36835 = n36844 & n36845;
  assign n36703 = ~n36750;
  assign n36745 = n36751 & n33978;
  assign n36732 = ~n36729;
  assign n36752 = n36781 ^ n36782;
  assign n36734 = n36791 ^ n36792;
  assign n36783 = ~n36781;
  assign n36773 = ~n36795;
  assign n35472 = n33270 ^ n34409;
  assign n36805 = n36815 & n36816;
  assign n36806 = n33270 & n36817;
  assign n33234 = ~n33270;
  assign n36827 = ~n36835;
  assign n36728 = ~n36745;
  assign n36730 = n373 ^ n36752;
  assign n36768 = n36734 & n372;
  assign n36775 = n36783 & n36784;
  assign n36767 = ~n36734;
  assign n36693 = n35472 ^ n35434;
  assign n36793 = ~n36805;
  assign n36796 = n33234 & n35509;
  assign n35511 = ~n36806;
  assign n36807 = n36827 & n36828;
  assign n36726 = n36728 & n36701;
  assign n36700 = n36728 & n36703;
  assign n36719 = n36729 ^ n36730;
  assign n36731 = ~n36730;
  assign n36755 = n36767 & n4120;
  assign n36707 = ~n36768;
  assign n36757 = n36693 & n36769;
  assign n36753 = ~n36775;
  assign n36756 = ~n36693;
  assign n36770 = n36793 & n36794;
  assign n35544 = ~n36796;
  assign n36785 = n36807 ^ n34368;
  assign n36808 = ~n36807;
  assign n32951 = n36700 ^ n36701;
  assign n36704 = n36719 & n33967;
  assign n36702 = ~n36726;
  assign n36651 = ~n36719;
  assign n36682 = n36731 & n36732;
  assign n36733 = n36753 & n36754;
  assign n36736 = ~n36755;
  assign n36746 = n36756 & n36723;
  assign n36695 = ~n36757;
  assign n36741 = n36770 ^ n36771;
  assign n36772 = ~n36770;
  assign n33194 = n36785 ^ n36786;
  assign n36797 = n36808 & n36809;
  assign n36648 = n32951 ^ n36678;
  assign n32935 = ~n32951;
  assign n36679 = n36702 & n36703;
  assign n36696 = n36651 & n33929;
  assign n36680 = ~n36704;
  assign n36705 = n36733 ^ n36734;
  assign n36685 = n36741 ^ n36742;
  assign n36735 = ~n36733;
  assign n36725 = ~n36746;
  assign n35398 = n33194 ^ n34345;
  assign n36758 = n36772 & n36773;
  assign n36759 = n33194 & n36774;
  assign n33221 = ~n33194;
  assign n36787 = ~n36797;
  assign n36620 = n36647 ^ n36648;
  assign n36649 = n36648 & n36667;
  assign n36650 = n36679 ^ n33967;
  assign n36681 = ~n36679;
  assign n36653 = ~n36696;
  assign n36683 = n372 ^ n36705;
  assign n36721 = n36685 & n371;
  assign n36727 = n36735 & n36736;
  assign n36720 = ~n36685;
  assign n36640 = n35398 ^ n35319;
  assign n36743 = ~n36758;
  assign n36747 = n33221 & n35436;
  assign n35475 = ~n36759;
  assign n36760 = n36787 & n36788;
  assign n36609 = n36620 ^ n36621;
  assign n36637 = ~n36649;
  assign n32841 = n36650 ^ n36651;
  assign n36675 = n36680 & n36681;
  assign n36668 = n36682 ^ n36683;
  assign n36627 = n36683 & n36682;
  assign n36708 = n36720 & n4067;
  assign n36657 = ~n36721;
  assign n36711 = n36640 & n36672;
  assign n36706 = ~n36727;
  assign n36709 = ~n36640;
  assign n36722 = n36743 & n36744;
  assign n35439 = ~n36747;
  assign n36738 = n36760 ^ n34311;
  assign n36761 = ~n36760;
  assign n36586 = n36609 & n454;
  assign n36585 = ~n36609;
  assign n36556 = n36622 ^ n32841;
  assign n36623 = n36637 & n36638;
  assign n32893 = ~n32841;
  assign n36654 = n36668 & n33917;
  assign n36652 = ~n36675;
  assign n36591 = ~n36668;
  assign n36684 = n36706 & n36707;
  assign n36687 = ~n36708;
  assign n36697 = n36709 & n36710;
  assign n36642 = ~n36711;
  assign n36692 = n36722 ^ n36723;
  assign n36724 = ~n36722;
  assign n33192 = n36737 ^ n36738;
  assign n36748 = n36761 & n36762;
  assign n36579 = n36585 & n18650;
  assign n36520 = ~n36586;
  assign n36589 = n36556 & n36590;
  assign n36587 = ~n36556;
  assign n36558 = ~n36623;
  assign n36624 = n36652 & n36653;
  assign n36626 = ~n36654;
  assign n36644 = n36591 & n33941;
  assign n36655 = n36684 ^ n36685;
  assign n36630 = n36692 ^ n36693;
  assign n36686 = ~n36684;
  assign n36674 = ~n36697;
  assign n35322 = n33192 ^ n34311;
  assign n36712 = n36724 & n36725;
  assign n36713 = n33192 & n35362;
  assign n33155 = ~n33192;
  assign n36739 = ~n36748;
  assign n36554 = ~n36579;
  assign n36580 = n36587 & n36588;
  assign n36524 = ~n36589;
  assign n36555 = n36558 ^ n36590;
  assign n36592 = n36624 ^ n33917;
  assign n36625 = ~n36624;
  assign n36594 = ~n36644;
  assign n36628 = n371 ^ n36655;
  assign n36670 = n36630 & n370;
  assign n36676 = n36686 & n36687;
  assign n36669 = ~n36630;
  assign n36576 = n35322 ^ n35290;
  assign n36694 = ~n36712;
  assign n35364 = ~n36713;
  assign n36698 = n33155 & n36714;
  assign n36716 = n36739 & n36740;
  assign n36550 = n36554 & n36518;
  assign n36517 = n36554 & n36520;
  assign n36487 = n36555 ^ n36556;
  assign n36557 = ~n36580;
  assign n32831 = n36591 ^ n36592;
  assign n36617 = n36625 & n36626;
  assign n36528 = n36627 ^ n36628;
  assign n36563 = n36628 & n36627;
  assign n36658 = n36669 & n4032;
  assign n36599 = ~n36670;
  assign n36661 = n36576 & n36613;
  assign n36656 = ~n36676;
  assign n36659 = ~n36576;
  assign n36671 = n36694 & n36695;
  assign n35401 = ~n36698;
  assign n33163 = n36715 ^ n36716;
  assign n36717 = ~n36716;
  assign n34350 = n36517 ^ n36518;
  assign n36522 = n36487 & n453;
  assign n36519 = ~n36550;
  assign n36521 = ~n36487;
  assign n36551 = n36557 & n36558;
  assign n36449 = n36559 ^ n32831;
  assign n32785 = ~n32831;
  assign n36596 = n36528 & n33886;
  assign n36593 = ~n36617;
  assign n36595 = ~n36528;
  assign n36566 = ~n36563;
  assign n36629 = n36656 & n36657;
  assign n36632 = ~n36658;
  assign n36645 = n36659 & n36660;
  assign n36578 = ~n36661;
  assign n36639 = n36671 ^ n36672;
  assign n36673 = ~n36671;
  assign n35242 = n33163 ^ n34253;
  assign n36689 = n33163 & n35283;
  assign n33098 = ~n33163;
  assign n36699 = n36717 & n36718;
  assign n35244 = ~n34350;
  assign n36486 = n36519 & n36520;
  assign n36512 = n36521 & n18542;
  assign n36451 = ~n36522;
  assign n36527 = n36449 & n36491;
  assign n36523 = ~n36551;
  assign n36525 = ~n36449;
  assign n36560 = n36593 & n36594;
  assign n36581 = n36595 & n33910;
  assign n36561 = ~n36596;
  assign n36597 = n36629 ^ n36630;
  assign n36568 = n36639 ^ n36640;
  assign n36631 = ~n36629;
  assign n36615 = ~n36645;
  assign n36546 = n35242 ^ n35119;
  assign n36662 = n36673 & n36674;
  assign n36677 = n33098 & n36688;
  assign n35327 = ~n36689;
  assign n36690 = ~n36699;
  assign n36447 = n36486 ^ n36487;
  assign n36488 = ~n36486;
  assign n36489 = ~n36512;
  assign n36490 = n36523 & n36524;
  assign n36513 = n36525 & n36526;
  assign n36492 = ~n36527;
  assign n36529 = n36560 ^ n33910;
  assign n36562 = ~n36560;
  assign n36531 = ~n36581;
  assign n36564 = n370 ^ n36597;
  assign n36610 = n36568 & n3990;
  assign n36618 = n36631 & n36632;
  assign n36611 = ~n36568;
  assign n36633 = n36546 & n36643;
  assign n36634 = ~n36546;
  assign n36641 = ~n36662;
  assign n35285 = ~n36677;
  assign n36663 = n36690 & n36691;
  assign n34335 = n453 ^ n36447;
  assign n36482 = n36488 & n36489;
  assign n36448 = n36490 ^ n36491;
  assign n36493 = ~n36490;
  assign n36453 = ~n36513;
  assign n32731 = n36528 ^ n36529;
  assign n36552 = n36561 & n36562;
  assign n36457 = n36563 ^ n36564;
  assign n36565 = ~n36564;
  assign n36570 = ~n36610;
  assign n36600 = n36611 & n369;
  assign n36598 = ~n36618;
  assign n36548 = ~n36633;
  assign n36619 = n36634 & n36509;
  assign n36612 = n36641 & n36642;
  assign n35163 = n36663 ^ n36664;
  assign n36665 = ~n36663;
  assign n35164 = ~n34335;
  assign n36416 = n36448 ^ n36449;
  assign n36450 = ~n36482;
  assign n36483 = n36492 & n36493;
  assign n36379 = n36494 ^ n32731;
  assign n32775 = ~n32731;
  assign n36533 = n36457 & n33853;
  assign n36530 = ~n36552;
  assign n36532 = ~n36457;
  assign n36498 = n36565 & n36566;
  assign n36567 = n36598 & n36599;
  assign n36536 = ~n36600;
  assign n36575 = n36612 ^ n36613;
  assign n36511 = ~n36619;
  assign n36614 = ~n36612;
  assign n36478 = n35163 ^ n35135;
  assign n33047 = n34216 ^ n35163;
  assign n36646 = n36665 & n36666;
  assign n36417 = n36416 & n18500;
  assign n36418 = ~n36416;
  assign n36415 = n36450 & n36451;
  assign n36455 = n36379 & n36474;
  assign n36452 = ~n36483;
  assign n36454 = ~n36379;
  assign n36495 = n36530 & n36531;
  assign n36514 = n36532 & n33871;
  assign n36459 = ~n36533;
  assign n36534 = n36567 ^ n36568;
  assign n36501 = n36575 ^ n36576;
  assign n36569 = ~n36567;
  assign n36601 = n36614 & n36615;
  assign n36604 = n36478 & n36439;
  assign n36605 = n33047 & n36616;
  assign n36602 = ~n36478;
  assign n33116 = ~n33047;
  assign n36635 = ~n36646;
  assign n36376 = n36415 ^ n36416;
  assign n36400 = ~n36417;
  assign n36411 = n36418 & n452;
  assign n36401 = ~n36415;
  assign n36419 = n36452 & n36453;
  assign n36442 = n36454 & n36420;
  assign n36381 = ~n36455;
  assign n36456 = n36495 ^ n33871;
  assign n36496 = ~n36495;
  assign n36497 = ~n36514;
  assign n36499 = n369 ^ n36534;
  assign n36543 = n36501 & n3965;
  assign n36553 = n36569 & n36570;
  assign n36544 = ~n36501;
  assign n36577 = ~n36601;
  assign n36582 = n36602 & n36603;
  assign n36441 = ~n36604;
  assign n35207 = ~n36605;
  assign n36583 = n33116 & n35246;
  assign n36606 = n36635 & n36636;
  assign n36341 = n452 ^ n36376;
  assign n36377 = n36400 & n36401;
  assign n36364 = ~n36411;
  assign n36378 = n36419 ^ n36420;
  assign n36421 = ~n36419;
  assign n36422 = ~n36442;
  assign n32684 = n36456 ^ n36457;
  assign n36484 = n36496 & n36497;
  assign n36384 = n36498 ^ n36499;
  assign n36427 = n36499 & n36498;
  assign n36503 = ~n36543;
  assign n36537 = n36544 & n368;
  assign n36535 = ~n36553;
  assign n36545 = n36577 & n36578;
  assign n36480 = ~n36582;
  assign n35248 = ~n36583;
  assign n36572 = n36606 ^ n34174;
  assign n36607 = ~n36606;
  assign n34273 = n36341 ^ n35164;
  assign n36342 = ~n36341;
  assign n36363 = ~n36377;
  assign n36328 = n36378 ^ n36379;
  assign n36412 = n36421 & n36422;
  assign n36304 = n36423 ^ n32684;
  assign n32721 = ~n32684;
  assign n36460 = n36384 & n33820;
  assign n36458 = ~n36484;
  assign n36461 = ~n36384;
  assign n36430 = ~n36427;
  assign n36500 = n36535 & n36536;
  assign n36464 = ~n36537;
  assign n36508 = n36545 ^ n36546;
  assign n36547 = ~n36545;
  assign n33069 = n36571 ^ n36572;
  assign n36584 = n36607 & n36608;
  assign n35095 = ~n34273;
  assign n36250 = n36342 & n34335;
  assign n36327 = n36363 & n36364;
  assign n36344 = n36328 & n451;
  assign n36343 = ~n36328;
  assign n36382 = n36304 & n36402;
  assign n36380 = ~n36412;
  assign n36383 = ~n36304;
  assign n36424 = n36458 & n36459;
  assign n36387 = ~n36460;
  assign n36443 = n36461 & n33816;
  assign n36462 = n36500 ^ n36501;
  assign n36390 = n36508 ^ n36509;
  assign n36502 = ~n36500;
  assign n35083 = n33069 ^ n34174;
  assign n36538 = n36547 & n36548;
  assign n36539 = n33069 & n36549;
  assign n32998 = ~n33069;
  assign n36573 = ~n36584;
  assign n36288 = n36327 ^ n36328;
  assign n36253 = ~n36250;
  assign n36302 = ~n36327;
  assign n36337 = n36343 & n18450;
  assign n36269 = ~n36344;
  assign n36345 = n36380 & n36381;
  assign n36306 = ~n36382;
  assign n36370 = n36383 & n36346;
  assign n36385 = n36424 ^ n33816;
  assign n36425 = ~n36424;
  assign n36426 = ~n36443;
  assign n36428 = n368 ^ n36462;
  assign n36476 = n36390 & n383;
  assign n36485 = n36502 & n36503;
  assign n36475 = ~n36390;
  assign n36407 = n35045 ^ n35083;
  assign n36510 = ~n36538;
  assign n36515 = n32998 & n35124;
  assign n35168 = ~n36539;
  assign n36540 = n36573 & n36574;
  assign n36251 = n451 ^ n36288;
  assign n36301 = ~n36337;
  assign n36303 = n36345 ^ n36346;
  assign n36348 = ~n36345;
  assign n36347 = ~n36370;
  assign n32644 = n36384 ^ n36385;
  assign n36413 = n36425 & n36426;
  assign n36403 = n36427 ^ n36428;
  assign n36429 = ~n36428;
  assign n36465 = n36475 & n3911;
  assign n36392 = ~n36476;
  assign n36466 = n36407 & n36366;
  assign n36463 = ~n36485;
  assign n36467 = ~n36407;
  assign n36477 = n36510 & n36511;
  assign n35127 = ~n36515;
  assign n36504 = n36540 ^ n34157;
  assign n36541 = ~n36540;
  assign n34242 = n36250 ^ n36251;
  assign n36252 = ~n36251;
  assign n36296 = n36301 & n36302;
  assign n36226 = n36303 ^ n36304;
  assign n36338 = n36347 & n36348;
  assign n36230 = n36349 ^ n32644;
  assign n32667 = ~n32644;
  assign n36388 = n36403 & n33799;
  assign n36386 = ~n36413;
  assign n36311 = ~n36403;
  assign n36353 = n36429 & n36430;
  assign n36431 = n36463 & n36464;
  assign n36433 = ~n36465;
  assign n36409 = ~n36466;
  assign n36444 = n36467 & n36468;
  assign n36438 = n36477 ^ n36478;
  assign n36479 = ~n36477;
  assign n32974 = n36504 ^ n36505;
  assign n36516 = n36541 & n36542;
  assign n35013 = ~n34242;
  assign n36155 = n36252 & n36253;
  assign n36271 = n36226 & n450;
  assign n36268 = ~n36296;
  assign n36270 = ~n36226;
  assign n36307 = n36230 & n36273;
  assign n36305 = ~n36338;
  assign n36308 = ~n36230;
  assign n36350 = n36386 & n36387;
  assign n36371 = n36311 & n33754;
  assign n36352 = ~n36388;
  assign n36389 = n383 ^ n36431;
  assign n36356 = n36438 ^ n36439;
  assign n36432 = ~n36431;
  assign n36368 = ~n36444;
  assign n36469 = n36479 & n36480;
  assign n36470 = n32974 & n36481;
  assign n33008 = ~n32974;
  assign n36506 = ~n36516;
  assign n36225 = n36268 & n36269;
  assign n36264 = n36270 & n18410;
  assign n36197 = ~n36271;
  assign n36272 = n36305 & n36306;
  assign n36232 = ~n36307;
  assign n36297 = n36308 & n36309;
  assign n36310 = n36350 ^ n33799;
  assign n36351 = ~n36350;
  assign n36313 = ~n36371;
  assign n36354 = n36389 ^ n36390;
  assign n36404 = n36356 & n3849;
  assign n36414 = n36432 & n36433;
  assign n36405 = ~n36356;
  assign n35011 = n34181 ^ n33008;
  assign n36440 = ~n36469;
  assign n35087 = ~n36470;
  assign n36445 = n33008 & n35046;
  assign n36471 = n36506 & n36507;
  assign n36195 = n36225 ^ n36226;
  assign n36228 = ~n36225;
  assign n36227 = ~n36264;
  assign n36229 = n36272 ^ n36273;
  assign n36274 = ~n36272;
  assign n36275 = ~n36297;
  assign n32632 = n36310 ^ n36311;
  assign n36339 = n36351 & n36352;
  assign n36235 = n36353 ^ n36354;
  assign n36280 = n36354 & n36353;
  assign n36358 = ~n36404;
  assign n36393 = n36405 & n382;
  assign n36391 = ~n36414;
  assign n36291 = n35011 ^ n34927;
  assign n36406 = n36440 & n36441;
  assign n35049 = ~n36445;
  assign n36434 = n36471 ^ n34185;
  assign n36472 = ~n36471;
  assign n36156 = n450 ^ n36195;
  assign n36220 = n36227 & n36228;
  assign n36159 = n36229 ^ n36230;
  assign n36265 = n36274 & n36275;
  assign n36163 = n36276 ^ n32632;
  assign n32606 = ~n32632;
  assign n36315 = n36235 & n33732;
  assign n36312 = ~n36339;
  assign n36314 = ~n36235;
  assign n36289 = ~n36280;
  assign n36355 = n36391 & n36392;
  assign n36318 = ~n36393;
  assign n36372 = n36291 & n36394;
  assign n36365 = n36406 ^ n36407;
  assign n36373 = ~n36291;
  assign n36408 = ~n36406;
  assign n32972 = n36434 ^ n36435;
  assign n36446 = n36472 & n36473;
  assign n34224 = n36155 ^ n36156;
  assign n36157 = ~n36156;
  assign n36198 = n36159 & n18389;
  assign n36196 = ~n36220;
  assign n36199 = ~n36159;
  assign n36234 = n36163 & n36254;
  assign n36231 = ~n36265;
  assign n36233 = ~n36163;
  assign n36277 = n36312 & n36313;
  assign n36298 = n36314 & n33765;
  assign n36278 = ~n36315;
  assign n36316 = n36355 ^ n36356;
  assign n36283 = n36365 ^ n36366;
  assign n36357 = ~n36355;
  assign n36293 = ~n36372;
  assign n36369 = n36373 & n36333;
  assign n34915 = n32972 ^ n34125;
  assign n36395 = n36408 & n36409;
  assign n36396 = n32972 & n36410;
  assign n32918 = ~n32972;
  assign n36436 = ~n36446;
  assign n34931 = ~n34224;
  assign n36093 = n36157 & n36155;
  assign n36158 = n36196 & n36197;
  assign n36160 = ~n36198;
  assign n36191 = n36199 & n449;
  assign n36200 = n36231 & n36232;
  assign n36221 = n36233 & n36201;
  assign n36165 = ~n36234;
  assign n36236 = n36277 ^ n33765;
  assign n36279 = ~n36277;
  assign n36238 = ~n36298;
  assign n36281 = n382 ^ n36316;
  assign n36329 = n36283 & n3787;
  assign n36340 = n36357 & n36358;
  assign n36330 = ~n36283;
  assign n36217 = n34915 ^ n34891;
  assign n36335 = ~n36369;
  assign n36367 = ~n36395;
  assign n36374 = n32918 & n34971;
  assign n34973 = ~n36396;
  assign n36397 = n36436 & n36437;
  assign n36127 = n36158 ^ n36159;
  assign n36161 = ~n36158;
  assign n36129 = ~n36191;
  assign n36162 = n36200 ^ n36201;
  assign n36202 = ~n36200;
  assign n36203 = ~n36221;
  assign n32594 = n36235 ^ n36236;
  assign n36266 = n36278 & n36279;
  assign n36170 = n36280 ^ n36281;
  assign n36208 = n36281 & n36289;
  assign n36285 = ~n36329;
  assign n36319 = n36330 & n381;
  assign n36320 = n36217 & n36331;
  assign n36317 = ~n36340;
  assign n36321 = ~n36217;
  assign n36332 = n36367 & n36368;
  assign n35016 = ~n36374;
  assign n36359 = n36397 ^ n34087;
  assign n36398 = ~n36397;
  assign n36094 = n449 ^ n36127;
  assign n36151 = n36160 & n36161;
  assign n36096 = n36162 ^ n36163;
  assign n36192 = n36202 & n36203;
  assign n36100 = n36204 ^ n32594;
  assign n32576 = ~n32594;
  assign n36239 = n36170 & n33697;
  assign n36237 = ~n36266;
  assign n36240 = ~n36170;
  assign n36211 = ~n36208;
  assign n36282 = n36317 & n36318;
  assign n36243 = ~n36319;
  assign n36219 = ~n36320;
  assign n36299 = n36321 & n36258;
  assign n36290 = n36332 ^ n36333;
  assign n36334 = ~n36332;
  assign n32857 = n36359 ^ n36360;
  assign n36375 = n36398 & n36399;
  assign n34161 = n36093 ^ n36094;
  assign n36034 = n36094 & n36093;
  assign n36131 = n36096 & n448;
  assign n36128 = ~n36151;
  assign n36130 = ~n36096;
  assign n36168 = n36100 & n36133;
  assign n36164 = ~n36192;
  assign n36166 = ~n36100;
  assign n36205 = n36237 & n36238;
  assign n36207 = ~n36239;
  assign n36222 = n36240 & n33730;
  assign n36241 = n36282 ^ n36283;
  assign n36213 = n36290 ^ n36291;
  assign n36284 = ~n36282;
  assign n36259 = ~n36299;
  assign n34847 = n34107 ^ n32857;
  assign n36322 = n36334 & n36335;
  assign n36323 = n32857 & n34893;
  assign n32905 = ~n32857;
  assign n36361 = ~n36375;
  assign n34848 = ~n34161;
  assign n36095 = n36128 & n36129;
  assign n36123 = n36130 & n18335;
  assign n36067 = ~n36131;
  assign n36132 = n36164 & n36165;
  assign n36152 = n36166 & n36167;
  assign n36135 = ~n36168;
  assign n36169 = n36205 ^ n33697;
  assign n36206 = ~n36205;
  assign n36172 = ~n36222;
  assign n36209 = n381 ^ n36241;
  assign n36256 = n36213 & n380;
  assign n36267 = n36284 & n36285;
  assign n36255 = ~n36213;
  assign n36147 = n34847 ^ n34757;
  assign n36292 = ~n36322;
  assign n34895 = ~n36323;
  assign n36300 = n32905 & n36324;
  assign n36325 = n36361 & n36362;
  assign n36065 = n36095 ^ n36096;
  assign n36098 = ~n36095;
  assign n36097 = ~n36123;
  assign n36099 = n36132 ^ n36133;
  assign n36134 = ~n36132;
  assign n36102 = ~n36152;
  assign n32541 = n36169 ^ n36170;
  assign n36193 = n36206 & n36207;
  assign n36107 = n36208 ^ n36209;
  assign n36210 = ~n36209;
  assign n36244 = n36255 & n3736;
  assign n36177 = ~n36256;
  assign n36245 = n36147 & n36186;
  assign n36242 = ~n36267;
  assign n36246 = ~n36147;
  assign n36257 = n36292 & n36293;
  assign n34934 = ~n36300;
  assign n36286 = n36325 ^ n34057;
  assign n36326 = n36325 & n36336;
  assign n36035 = n448 ^ n36065;
  assign n36090 = n36097 & n36098;
  assign n36038 = n36099 ^ n36100;
  assign n36124 = n36134 & n36135;
  assign n36042 = n36136 ^ n32541;
  assign n32564 = ~n32541;
  assign n36173 = n36107 & n33661;
  assign n36171 = ~n36193;
  assign n36174 = ~n36107;
  assign n36140 = n36210 & n36211;
  assign n36212 = n36242 & n36243;
  assign n36215 = ~n36244;
  assign n36188 = ~n36245;
  assign n36223 = n36246 & n36247;
  assign n36216 = n36257 ^ n36258;
  assign n36260 = ~n36257;
  assign n32855 = n36286 ^ n36287;
  assign n36294 = ~n36326;
  assign n34143 = n36034 ^ n36035;
  assign n36036 = ~n36035;
  assign n36068 = n36038 & n18294;
  assign n36066 = ~n36090;
  assign n36069 = ~n36038;
  assign n36103 = n36042 & n36071;
  assign n36101 = ~n36124;
  assign n36104 = ~n36042;
  assign n36137 = n36171 & n36172;
  assign n36139 = ~n36173;
  assign n36153 = n36174 & n33695;
  assign n36175 = n36212 ^ n36213;
  assign n36143 = n36216 ^ n36217;
  assign n36214 = ~n36212;
  assign n36150 = ~n36223;
  assign n34770 = n34116 ^ n32855;
  assign n36248 = n36259 & n36260;
  assign n36249 = n32855 & n36261;
  assign n32798 = ~n32855;
  assign n36262 = n36294 & n36295;
  assign n34785 = ~n34143;
  assign n34702 = n36036 & n36034;
  assign n36037 = n36066 & n36067;
  assign n36040 = ~n36068;
  assign n36061 = n36069 & n463;
  assign n36070 = n36101 & n36102;
  assign n36072 = ~n36103;
  assign n36091 = n36104 & n36105;
  assign n36106 = n36137 ^ n33661;
  assign n36138 = ~n36137;
  assign n36109 = ~n36153;
  assign n36141 = n380 ^ n36175;
  assign n36184 = n36143 & n379;
  assign n36194 = n36214 & n36215;
  assign n36183 = ~n36143;
  assign n36087 = n34770 ^ n34691;
  assign n36218 = ~n36248;
  assign n34811 = ~n36249;
  assign n36224 = n32798 & n34808;
  assign n34074 = n36262 ^ n36263;
  assign n36008 = n36037 ^ n36038;
  assign n36039 = ~n36037;
  assign n36010 = ~n36061;
  assign n36041 = n36070 ^ n36071;
  assign n36073 = ~n36070;
  assign n36044 = ~n36091;
  assign n32504 = n36106 ^ n36107;
  assign n36125 = n36138 & n36139;
  assign n36048 = n36140 ^ n36141;
  assign n36078 = n36141 & n36140;
  assign n36178 = n36183 & n3634;
  assign n36114 = ~n36184;
  assign n36181 = n36087 & n36120;
  assign n36176 = ~n36194;
  assign n36179 = ~n36087;
  assign n36185 = n36218 & n36219;
  assign n36189 = n34074 ^ n34060;
  assign n34852 = ~n36224;
  assign n34669 = n463 ^ n36008;
  assign n36031 = n36039 & n36040;
  assign n35985 = n36041 ^ n36042;
  assign n36062 = n36072 & n36073;
  assign n35989 = n36074 ^ n32504;
  assign n32523 = ~n32504;
  assign n36111 = n36048 & n33623;
  assign n36108 = ~n36125;
  assign n36110 = ~n36048;
  assign n36081 = ~n36078;
  assign n36142 = n36176 & n36177;
  assign n36145 = ~n36178;
  assign n36154 = n36179 & n36180;
  assign n36089 = ~n36181;
  assign n36146 = n36185 ^ n36186;
  assign n34701 = n36189 ^ n36190;
  assign n36187 = ~n36185;
  assign n35939 = n34669 & n34702;
  assign n36011 = n35985 & n18263;
  assign n36009 = ~n36031;
  assign n36012 = ~n35985;
  assign n36045 = n35989 & n36014;
  assign n36043 = ~n36062;
  assign n36046 = ~n35989;
  assign n36075 = n36108 & n36109;
  assign n36092 = n36110 & n33659;
  assign n36076 = ~n36111;
  assign n36112 = n36142 ^ n36143;
  assign n36083 = n36146 ^ n36147;
  assign n36030 = n36148 ^ n34701;
  assign n36144 = ~n36142;
  assign n36122 = ~n36154;
  assign n36182 = n36187 & n36188;
  assign n35984 = n36009 & n36010;
  assign n35987 = ~n36011;
  assign n36004 = n36012 & n462;
  assign n36013 = n36043 & n36044;
  assign n36016 = ~n36045;
  assign n36032 = n36046 & n36047;
  assign n36049 = n36075 ^ n33659;
  assign n36077 = ~n36075;
  assign n36051 = ~n36092;
  assign n36079 = n379 ^ n36112;
  assign n36117 = n36083 & n3578;
  assign n36126 = n36144 & n36145;
  assign n36118 = ~n36083;
  assign n36149 = ~n36182;
  assign n35963 = n35984 ^ n35985;
  assign n35986 = ~n35984;
  assign n35965 = ~n36004;
  assign n35988 = n36013 ^ n36014;
  assign n36015 = ~n36013;
  assign n35991 = ~n36032;
  assign n32468 = n36048 ^ n36049;
  assign n36063 = n36076 & n36077;
  assign n35996 = n36078 ^ n36079;
  assign n36080 = ~n36079;
  assign n36084 = ~n36117;
  assign n36115 = n36118 & n378;
  assign n36113 = ~n36126;
  assign n36119 = n36149 & n36150;
  assign n35940 = n462 ^ n35963;
  assign n35981 = n35986 & n35987;
  assign n35942 = n35988 ^ n35989;
  assign n36005 = n36015 & n36016;
  assign n35946 = n36017 ^ n32468;
  assign n32473 = ~n32468;
  assign n36053 = n35996 & n33621;
  assign n36050 = ~n36063;
  assign n36052 = ~n35996;
  assign n36021 = n36080 & n36081;
  assign n36082 = n36113 & n36114;
  assign n36056 = ~n36115;
  assign n36086 = n36119 ^ n36120;
  assign n36121 = ~n36119;
  assign n33110 = n35939 ^ n35940;
  assign n35897 = n35940 & n35939;
  assign n35966 = n35942 & n18218;
  assign n35964 = ~n35981;
  assign n35967 = ~n35942;
  assign n35992 = n35946 & n35969;
  assign n35990 = ~n36005;
  assign n35993 = ~n35946;
  assign n36018 = n36050 & n36051;
  assign n36033 = n36052 & n33585;
  assign n35998 = ~n36053;
  assign n36024 = ~n36021;
  assign n36054 = n36082 ^ n36083;
  assign n36026 = n36086 ^ n36087;
  assign n36085 = ~n36082;
  assign n36116 = n36121 & n36122;
  assign n35913 = n34029 ^ n33110;
  assign n32155 = n33088 ^ n33110;
  assign n35896 = n35920 ^ n33110;
  assign n35828 = n33110 & n33088;
  assign n35941 = n35964 & n35965;
  assign n35944 = ~n35966;
  assign n35960 = n35967 & n461;
  assign n35968 = n35990 & n35991;
  assign n35948 = ~n35992;
  assign n35982 = n35993 & n35994;
  assign n35995 = n36018 ^ n33585;
  assign n36019 = ~n36018;
  assign n36020 = ~n36033;
  assign n36022 = n378 ^ n36054;
  assign n36058 = n36026 & n3502;
  assign n36064 = n36084 & n36085;
  assign n36059 = ~n36026;
  assign n36088 = ~n36116;
  assign n33938 = n39 ^ n35896;
  assign n35754 = n35913 & n35914;
  assign n35629 = n35896 & n39;
  assign n35921 = n35941 ^ n35942;
  assign n35943 = ~n35941;
  assign n35923 = ~n35960;
  assign n35945 = n35968 ^ n35969;
  assign n35970 = ~n35968;
  assign n35971 = ~n35982;
  assign n32444 = n35995 ^ n35996;
  assign n36006 = n36019 & n36020;
  assign n36003 = n36021 ^ n36022;
  assign n36023 = ~n36022;
  assign n36028 = ~n36058;
  assign n36057 = n36059 & n377;
  assign n36055 = ~n36064;
  assign n36060 = n36088 & n36089;
  assign n35892 = n35754 & n35729;
  assign n35637 = ~n33938;
  assign n35890 = ~n35754;
  assign n35898 = n461 ^ n35921;
  assign n35936 = n35943 & n35944;
  assign n35900 = n35945 ^ n35946;
  assign n35961 = n35970 & n35971;
  assign n35904 = n35972 ^ n32444;
  assign n32423 = ~n32444;
  assign n35999 = n36003 & n33547;
  assign n35997 = ~n36006;
  assign n35951 = ~n36003;
  assign n35976 = n36023 & n36024;
  assign n36025 = n36055 & n36056;
  assign n36002 = ~n36057;
  assign n36029 = n376 ^ n36060;
  assign n35874 = n35890 & n35891;
  assign n35751 = ~n35892;
  assign n35893 = n35897 ^ n35898;
  assign n35851 = n35898 & n35897;
  assign n35924 = n35900 & n18199;
  assign n35922 = ~n35936;
  assign n35925 = ~n35900;
  assign n35949 = n35904 & n35959;
  assign n35947 = ~n35961;
  assign n35950 = ~n35904;
  assign n35973 = n35997 & n35998;
  assign n35975 = ~n35999;
  assign n35983 = n35951 & n33572;
  assign n36000 = n36025 ^ n36026;
  assign n35980 = n36029 ^ n36030;
  assign n36027 = ~n36025;
  assign n35773 = ~n35874;
  assign n35875 = n35893 & n32951;
  assign n35876 = ~n35893;
  assign n35854 = ~n35851;
  assign n35899 = n35922 & n35923;
  assign n35902 = ~n35924;
  assign n35916 = n35925 & n460;
  assign n35926 = n35947 & n35948;
  assign n35906 = ~n35949;
  assign n35937 = n35950 & n35927;
  assign n35952 = n35973 ^ n33547;
  assign n35974 = ~n35973;
  assign n35954 = ~n35983;
  assign n35977 = n377 ^ n36000;
  assign n36007 = n36027 & n36028;
  assign n35830 = ~n35875;
  assign n35870 = n35876 & n32935;
  assign n35877 = n35899 ^ n35900;
  assign n35901 = ~n35899;
  assign n35879 = ~n35916;
  assign n35903 = n35926 ^ n35927;
  assign n35929 = ~n35926;
  assign n35928 = ~n35937;
  assign n32420 = n35951 ^ n35952;
  assign n35962 = n35974 & n35975;
  assign n35909 = n35976 ^ n35977;
  assign n35978 = ~n35977;
  assign n36001 = ~n36007;
  assign n35850 = ~n35870;
  assign n35852 = n460 ^ n35877;
  assign n35894 = n35901 & n35902;
  assign n35856 = n35903 ^ n35904;
  assign n35917 = n35928 & n35929;
  assign n35860 = n35930 ^ n32420;
  assign n32391 = ~n32420;
  assign n35955 = n35909 & n33534;
  assign n35953 = ~n35962;
  assign n35956 = ~n35909;
  assign n35957 = n35978 & n35976;
  assign n35979 = n36001 & n36002;
  assign n35847 = n35850 & n35828;
  assign n35827 = n35850 & n35830;
  assign n35846 = n35851 ^ n35852;
  assign n35853 = ~n35852;
  assign n35881 = n35856 & n459;
  assign n35878 = ~n35894;
  assign n35880 = ~n35856;
  assign n35908 = n35860 & n35915;
  assign n35905 = ~n35917;
  assign n35907 = ~n35860;
  assign n35931 = n35953 & n35954;
  assign n35912 = ~n35955;
  assign n35938 = n35956 & n33507;
  assign n35958 = n35979 ^ n35980;
  assign n31985 = n35827 ^ n35828;
  assign n35831 = n35846 & n32893;
  assign n35829 = ~n35847;
  assign n35780 = ~n35846;
  assign n35807 = n35853 & n35854;
  assign n35855 = n35878 & n35879;
  assign n35871 = n35880 & n18144;
  assign n35834 = ~n35881;
  assign n35882 = n35905 & n35906;
  assign n35895 = n35907 & n35883;
  assign n35862 = ~n35908;
  assign n35910 = n35931 ^ n33507;
  assign n35932 = ~n35931;
  assign n35933 = ~n35938;
  assign n35865 = n35957 ^ n35958;
  assign n33987 = n32951 ^ n31985;
  assign n32133 = ~n31985;
  assign n35804 = n35829 & n35830;
  assign n35805 = ~n35831;
  assign n35823 = n35780 & n32841;
  assign n35832 = n35855 ^ n35856;
  assign n35857 = ~n35855;
  assign n35858 = ~n35871;
  assign n35859 = n35882 ^ n35883;
  assign n35884 = ~n35882;
  assign n35885 = ~n35895;
  assign n32355 = n35909 ^ n35910;
  assign n35918 = n35932 & n35933;
  assign n35934 = n35865 & n33505;
  assign n35935 = ~n35865;
  assign n35755 = n33987 ^ n33982;
  assign n35779 = n35804 ^ n32893;
  assign n35806 = ~n35804;
  assign n35782 = ~n35823;
  assign n35808 = n459 ^ n35832;
  assign n35848 = n35857 & n35858;
  assign n35810 = n35859 ^ n35860;
  assign n35872 = n35884 & n35885;
  assign n35814 = n35886 ^ n32355;
  assign n32374 = ~n32355;
  assign n35911 = ~n35918;
  assign n35868 = ~n35934;
  assign n35919 = n35935 & n33463;
  assign n35728 = n35754 ^ n35755;
  assign n35756 = n35755 & n35773;
  assign n31956 = n35779 ^ n35780;
  assign n35801 = n35805 & n35806;
  assign n35800 = n35807 ^ n35808;
  assign n35760 = n35808 & n35807;
  assign n35836 = n35810 & n458;
  assign n35833 = ~n35848;
  assign n35835 = ~n35810;
  assign n35864 = n35814 & n35869;
  assign n35861 = ~n35872;
  assign n35863 = ~n35814;
  assign n35887 = n35911 & n35912;
  assign n35889 = ~n35919;
  assign n35721 = n35728 ^ n35729;
  assign n35750 = ~n35756;
  assign n33974 = n31956 ^ n32841;
  assign n31975 = ~n31956;
  assign n35783 = n35800 & n32785;
  assign n35781 = ~n35801;
  assign n35732 = ~n35800;
  assign n35809 = n35833 & n35834;
  assign n35824 = n35835 & n18124;
  assign n35786 = ~n35836;
  assign n35837 = n35861 & n35862;
  assign n35849 = n35863 & n35838;
  assign n35816 = ~n35864;
  assign n35866 = n35887 ^ n33463;
  assign n35888 = ~n35887;
  assign n35698 = n35721 & n38;
  assign n35697 = ~n35721;
  assign n35666 = n33974 ^ n33967;
  assign n35730 = n35750 & n35751;
  assign n35757 = n35781 & n35782;
  assign n35758 = ~n35783;
  assign n35774 = n35732 & n32831;
  assign n35784 = n35809 ^ n35810;
  assign n35811 = ~n35809;
  assign n35812 = ~n35824;
  assign n35813 = n35837 ^ n35838;
  assign n35839 = ~n35837;
  assign n35840 = ~n35849;
  assign n32342 = n35865 ^ n35866;
  assign n35873 = n35888 & n35889;
  assign n35691 = n35697 & n12610;
  assign n35631 = ~n35698;
  assign n35701 = n35666 & n35722;
  assign n35699 = ~n35666;
  assign n35689 = ~n35730;
  assign n35731 = n35757 ^ n32785;
  assign n35759 = ~n35757;
  assign n35734 = ~n35774;
  assign n35761 = n458 ^ n35784;
  assign n35802 = n35811 & n35812;
  assign n35763 = n35813 ^ n35814;
  assign n35825 = n35839 & n35840;
  assign n35767 = n35841 ^ n32342;
  assign n32317 = ~n32342;
  assign n35867 = ~n35873;
  assign n35665 = ~n35691;
  assign n35692 = n35699 & n35700;
  assign n35688 = ~n35701;
  assign n35667 = n35689 ^ n35700;
  assign n31910 = n35731 ^ n35732;
  assign n35752 = n35758 & n35759;
  assign n35669 = n35760 ^ n35761;
  assign n35705 = n35761 & n35760;
  assign n35788 = n35763 & n457;
  assign n35785 = ~n35802;
  assign n35787 = ~n35763;
  assign n35819 = n35767 & n35790;
  assign n35815 = ~n35825;
  assign n35817 = ~n35767;
  assign n35842 = n35867 & n35868;
  assign n35660 = n35665 & n35629;
  assign n35628 = n35665 & n35631;
  assign n35593 = n35666 ^ n35667;
  assign n35668 = n35688 & n35689;
  assign n35659 = ~n35692;
  assign n33950 = n32831 ^ n31910;
  assign n31874 = ~n31910;
  assign n35735 = n35669 & n32775;
  assign n35733 = ~n35752;
  assign n35736 = ~n35669;
  assign n35708 = ~n35705;
  assign n35762 = n35785 & n35786;
  assign n35775 = n35787 & n18059;
  assign n35739 = ~n35788;
  assign n35789 = n35815 & n35816;
  assign n35803 = n35817 & n35818;
  assign n35792 = ~n35819;
  assign n32262 = n35842 ^ n35843;
  assign n35844 = ~n35842;
  assign n33906 = n35628 ^ n35629;
  assign n35632 = n35593 & n12533;
  assign n35630 = ~n35660;
  assign n35633 = ~n35593;
  assign n35658 = ~n35668;
  assign n35583 = n33950 ^ n33917;
  assign n35702 = n35733 & n35734;
  assign n35703 = ~n35735;
  assign n35723 = n35736 & n32731;
  assign n35737 = n35762 ^ n35763;
  assign n35764 = ~n35762;
  assign n35765 = ~n35775;
  assign n35766 = n35789 ^ n35790;
  assign n35791 = ~n35789;
  assign n35769 = ~n35803;
  assign n35743 = n35820 ^ n32262;
  assign n32328 = ~n32262;
  assign n35826 = n35844 & n35845;
  assign n35558 = ~n33906;
  assign n35592 = n35630 & n35631;
  assign n35595 = ~n35632;
  assign n35622 = n35633 & n37;
  assign n35618 = n35658 & n35659;
  assign n35636 = n35583 & n35619;
  assign n35634 = ~n35583;
  assign n35670 = n35702 ^ n32731;
  assign n35704 = ~n35702;
  assign n35672 = ~n35723;
  assign n35706 = n457 ^ n35737;
  assign n35753 = n35764 & n35765;
  assign n35710 = n35766 ^ n35767;
  assign n35776 = n35791 & n35792;
  assign n35793 = n35743 & n35714;
  assign n35794 = ~n35743;
  assign n35821 = ~n35826;
  assign n35554 = n35592 ^ n35593;
  assign n35582 = n35618 ^ n35619;
  assign n35594 = ~n35592;
  assign n35556 = ~n35622;
  assign n35621 = ~n35618;
  assign n35623 = n35634 & n35635;
  assign n35620 = ~n35636;
  assign n31786 = n35669 ^ n35670;
  assign n35693 = n35703 & n35704;
  assign n35598 = n35705 ^ n35706;
  assign n35707 = ~n35706;
  assign n35740 = n35710 & n18051;
  assign n35738 = ~n35753;
  assign n35741 = ~n35710;
  assign n35768 = ~n35776;
  assign n35716 = ~n35793;
  assign n35777 = n35794 & n35795;
  assign n35796 = n35821 & n35822;
  assign n33848 = n37 ^ n35554;
  assign n35524 = n35582 ^ n35583;
  assign n35587 = n35594 & n35595;
  assign n35596 = n35620 & n35621;
  assign n35585 = ~n35623;
  assign n33924 = n31786 ^ n32731;
  assign n35638 = n31786 & n33938;
  assign n31784 = ~n31786;
  assign n35673 = n35598 & n32684;
  assign n35671 = ~n35693;
  assign n35674 = ~n35598;
  assign n35642 = n35707 & n35708;
  assign n35709 = n35738 & n35739;
  assign n35711 = ~n35740;
  assign n35724 = n35741 & n456;
  assign n35742 = n35768 & n35769;
  assign n35745 = ~n35777;
  assign n35770 = n35796 ^ n35797;
  assign n35798 = ~n35796;
  assign n35545 = n35524 & n12419;
  assign n33876 = ~n33848;
  assign n35546 = ~n35524;
  assign n35555 = ~n35587;
  assign n35584 = ~n35596;
  assign n35514 = n33924 ^ n33910;
  assign n35624 = n31784 & n35637;
  assign n33940 = ~n35638;
  assign n35639 = n35671 & n35672;
  assign n35600 = ~n35673;
  assign n35661 = n35674 & n32721;
  assign n35675 = n35709 ^ n35710;
  assign n35712 = ~n35709;
  assign n35677 = ~n35724;
  assign n35713 = n35742 ^ n35743;
  assign n35744 = ~n35742;
  assign n32222 = n35770 ^ n33371;
  assign n35778 = n35798 & n35799;
  assign n35517 = ~n35545;
  assign n35525 = n35546 & n36;
  assign n35523 = n35555 & n35556;
  assign n35547 = n35584 & n35585;
  assign n35559 = n35514 & n35548;
  assign n35560 = ~n35514;
  assign n33953 = ~n35624;
  assign n35597 = n35639 ^ n32721;
  assign n35640 = ~n35639;
  assign n35641 = ~n35661;
  assign n35643 = n456 ^ n35675;
  assign n35694 = n35711 & n35712;
  assign n35604 = n35713 ^ n35714;
  assign n35725 = n35744 & n35745;
  assign n32311 = ~n32222;
  assign n35771 = ~n35778;
  assign n35486 = n35523 ^ n35524;
  assign n35481 = ~n35525;
  assign n35513 = n35547 ^ n35548;
  assign n35518 = ~n35523;
  assign n35527 = ~n35547;
  assign n35488 = ~n35559;
  assign n35550 = n35560 & n35561;
  assign n31705 = n35597 ^ n35598;
  assign n35625 = n35640 & n35641;
  assign n35529 = n35642 ^ n35643;
  assign n35565 = n35643 & n35642;
  assign n35678 = n35604 & n17983;
  assign n35676 = ~n35694;
  assign n35679 = ~n35604;
  assign n35715 = ~n35725;
  assign n35681 = n35726 ^ n32311;
  assign n35746 = n35771 & n35772;
  assign n35452 = n36 ^ n35486;
  assign n35444 = n35513 ^ n35514;
  assign n35512 = n35517 & n35518;
  assign n35526 = ~n35550;
  assign n33889 = n31705 ^ n32684;
  assign n35557 = n31705 & n33906;
  assign n31703 = ~n31705;
  assign n35601 = n35529 & n32644;
  assign n35599 = ~n35625;
  assign n35602 = ~n35529;
  assign n35568 = ~n35565;
  assign n35644 = n35676 & n35677;
  assign n35646 = ~n35678;
  assign n35662 = n35679 & n471;
  assign n35680 = n35715 & n35716;
  assign n35696 = n35681 & n35717;
  assign n35695 = ~n35681;
  assign n35718 = n35746 ^ n35747;
  assign n35748 = ~n35746;
  assign n33827 = n35452 ^ n33848;
  assign n35370 = n35452 & n33848;
  assign n35476 = n35444 & n12343;
  assign n35477 = ~n35444;
  assign n35480 = ~n35512;
  assign n35519 = n35526 & n35527;
  assign n35415 = n33889 ^ n33853;
  assign n33908 = ~n35557;
  assign n35549 = n31703 & n35558;
  assign n35562 = n35599 & n35600;
  assign n35531 = ~n35601;
  assign n35588 = n35602 & n32667;
  assign n35603 = n471 ^ n35644;
  assign n35645 = ~n35644;
  assign n35606 = ~n35662;
  assign n35647 = n35680 ^ n35681;
  assign n35682 = ~n35680;
  assign n35690 = n35695 & n35648;
  assign n35683 = ~n35696;
  assign n32237 = n35718 ^ n33332;
  assign n35727 = n35748 & n35749;
  assign n35413 = ~n33827;
  assign n35445 = ~n35476;
  assign n35453 = n35477 & n35;
  assign n35443 = n35480 & n35481;
  assign n35490 = n35415 & n35515;
  assign n35487 = ~n35519;
  assign n35489 = ~n35415;
  assign n33927 = ~n35549;
  assign n35528 = n35562 ^ n32667;
  assign n35563 = ~n35562;
  assign n35564 = ~n35588;
  assign n35566 = n35603 ^ n35604;
  assign n35626 = n35645 & n35646;
  assign n35570 = n35647 ^ n35648;
  assign n35663 = n35682 & n35683;
  assign n35610 = n35684 ^ n32237;
  assign n35650 = ~n35690;
  assign n32186 = ~n32237;
  assign n35719 = ~n35727;
  assign n35407 = n35443 ^ n35444;
  assign n35409 = ~n35453;
  assign n35446 = ~n35443;
  assign n35454 = n35487 & n35488;
  assign n35482 = n35489 & n35455;
  assign n35417 = ~n35490;
  assign n31706 = n35528 ^ n35529;
  assign n35551 = n35563 & n35564;
  assign n35459 = n35565 ^ n35566;
  assign n35567 = ~n35566;
  assign n35608 = n35570 & n470;
  assign n35605 = ~n35626;
  assign n35607 = ~n35570;
  assign n35651 = n35610 & n35574;
  assign n35649 = ~n35663;
  assign n35652 = ~n35610;
  assign n35685 = n35719 & n35720;
  assign n35371 = n35 ^ n35407;
  assign n35440 = n35445 & n35446;
  assign n35414 = n35454 ^ n35455;
  assign n35457 = ~n35454;
  assign n35456 = ~n35482;
  assign n33834 = n31706 ^ n32644;
  assign n31605 = ~n31706;
  assign n35530 = ~n35551;
  assign n35479 = ~n35459;
  assign n35494 = n35567 & n35568;
  assign n35569 = n35605 & n35606;
  assign n35589 = n35607 & n17956;
  assign n35534 = ~n35608;
  assign n35609 = n35649 & n35650;
  assign n35612 = ~n35651;
  assign n35627 = n35652 & n35653;
  assign n35655 = n35685 ^ n33312;
  assign n35686 = ~n35685;
  assign n33787 = n35370 ^ n35371;
  assign n35291 = n35371 & n35370;
  assign n35373 = n35414 ^ n35415;
  assign n35408 = ~n35440;
  assign n35447 = n35456 & n35457;
  assign n35341 = n33834 ^ n33816;
  assign n35491 = n35530 & n35531;
  assign n35497 = ~n35494;
  assign n35532 = n35569 ^ n35570;
  assign n35571 = ~n35569;
  assign n35572 = ~n35589;
  assign n35573 = n35609 ^ n35610;
  assign n35611 = ~n35609;
  assign n35576 = ~n35627;
  assign n32194 = n35654 ^ n35655;
  assign n35664 = n35686 & n35687;
  assign n35328 = ~n33787;
  assign n35381 = n35373 & n34;
  assign n35372 = n35408 & n35409;
  assign n35380 = ~n35373;
  assign n35420 = n35341 & n35383;
  assign n35416 = ~n35447;
  assign n35418 = ~n35341;
  assign n35458 = n35491 ^ n32606;
  assign n35493 = n35491 & n32606;
  assign n35492 = ~n35491;
  assign n35495 = n470 ^ n35532;
  assign n35552 = n35571 & n35572;
  assign n35499 = n35573 ^ n35574;
  assign n35590 = n35611 & n35612;
  assign n35503 = n35613 ^ n32194;
  assign n32172 = ~n32194;
  assign n35656 = ~n35664;
  assign n35333 = n35372 ^ n35373;
  assign n35374 = n35380 & n12231;
  assign n35303 = ~n35381;
  assign n35339 = ~n35372;
  assign n35382 = n35416 & n35417;
  assign n35410 = n35418 & n35419;
  assign n35385 = ~n35420;
  assign n31542 = n35458 ^ n35459;
  assign n35483 = n35492 & n32632;
  assign n35478 = ~n35493;
  assign n35367 = n35494 ^ n35495;
  assign n35496 = ~n35495;
  assign n35535 = n35499 & n17901;
  assign n35533 = ~n35552;
  assign n35536 = ~n35499;
  assign n35578 = n35503 & n35586;
  assign n35575 = ~n35590;
  assign n35577 = ~n35503;
  assign n35614 = n35656 & n35657;
  assign n35292 = n34 ^ n35333;
  assign n35338 = ~n35374;
  assign n35340 = n35382 ^ n35383;
  assign n35384 = ~n35382;
  assign n35343 = ~n35410;
  assign n35405 = n31542 & n35413;
  assign n33805 = n32632 ^ n31542;
  assign n31616 = ~n31542;
  assign n35460 = n35478 & n35479;
  assign n35462 = n35367 & n32594;
  assign n35442 = ~n35483;
  assign n35461 = ~n35367;
  assign n35421 = n35496 & n35497;
  assign n35498 = n35533 & n35534;
  assign n35500 = ~n35535;
  assign n35520 = n35536 & n469;
  assign n35537 = n35575 & n35576;
  assign n35553 = n35577 & n35538;
  assign n35505 = ~n35578;
  assign n35579 = n35614 ^ n35615;
  assign n35616 = ~n35614;
  assign n33771 = n35291 ^ n35292;
  assign n35293 = ~n35292;
  assign n35334 = n35338 & n35339;
  assign n35262 = n35340 ^ n35341;
  assign n35375 = n35384 & n35385;
  assign n35266 = n33805 ^ n33799;
  assign n33843 = ~n35405;
  assign n35406 = n31616 & n33827;
  assign n35441 = ~n35460;
  assign n35448 = n35461 & n32576;
  assign n35369 = ~n35462;
  assign n35424 = ~n35421;
  assign n35463 = n35498 ^ n35499;
  assign n35501 = ~n35498;
  assign n35465 = ~n35520;
  assign n35502 = n35537 ^ n35538;
  assign n35539 = ~n35537;
  assign n35540 = ~n35553;
  assign n32162 = n35579 ^ n33272;
  assign n35591 = n35616 & n35617;
  assign n35255 = ~n33771;
  assign n35183 = n35293 & n35291;
  assign n35304 = n35262 & n12170;
  assign n35302 = ~n35334;
  assign n35305 = ~n35262;
  assign n35345 = n35266 & n35365;
  assign n35342 = ~n35375;
  assign n35344 = ~n35266;
  assign n33829 = ~n35406;
  assign n35402 = n35441 & n35442;
  assign n35404 = ~n35448;
  assign n35422 = n469 ^ n35463;
  assign n35484 = n35500 & n35501;
  assign n35426 = n35502 ^ n35503;
  assign n35521 = n35539 & n35540;
  assign n35430 = n35541 ^ n32162;
  assign n32129 = ~n32162;
  assign n35580 = ~n35591;
  assign n35186 = ~n35183;
  assign n35261 = n35302 & n35303;
  assign n35263 = ~n35304;
  assign n35294 = n35305 & n33;
  assign n35306 = n35342 & n35343;
  assign n35335 = n35344 & n35307;
  assign n35268 = ~n35345;
  assign n35366 = n35402 ^ n32576;
  assign n35403 = ~n35402;
  assign n35286 = n35421 ^ n35422;
  assign n35423 = ~n35422;
  assign n35467 = n35426 & n468;
  assign n35464 = ~n35484;
  assign n35466 = ~n35426;
  assign n35506 = n35430 & n35516;
  assign n35504 = ~n35521;
  assign n35507 = ~n35430;
  assign n35542 = n35580 & n35581;
  assign n35224 = n35261 ^ n35262;
  assign n35264 = ~n35261;
  assign n35226 = ~n35294;
  assign n35265 = n35306 ^ n35307;
  assign n35308 = ~n35306;
  assign n35309 = ~n35335;
  assign n31552 = n35366 ^ n35367;
  assign n35386 = n35403 & n35404;
  assign n35388 = n35286 & n32541;
  assign n35387 = ~n35286;
  assign n35346 = n35423 & n35424;
  assign n35425 = n35464 & n35465;
  assign n35449 = n35466 & n17859;
  assign n35391 = ~n35467;
  assign n35468 = n35504 & n35505;
  assign n35432 = ~n35506;
  assign n35485 = n35507 & n35469;
  assign n35508 = n35542 ^ n33234;
  assign n35543 = ~n35542;
  assign n35184 = n33 ^ n35224;
  assign n35256 = n35263 & n35264;
  assign n35188 = n35265 ^ n35266;
  assign n35295 = n35308 & n35309;
  assign n33768 = n31552 ^ n32594;
  assign n35329 = n31552 & n33787;
  assign n31473 = ~n31552;
  assign n35368 = ~n35386;
  assign n35376 = n35387 & n32564;
  assign n35332 = ~n35388;
  assign n35349 = ~n35346;
  assign n35389 = n35425 ^ n35426;
  assign n35428 = ~n35425;
  assign n35427 = ~n35449;
  assign n35429 = n35468 ^ n35469;
  assign n35470 = ~n35468;
  assign n35471 = ~n35485;
  assign n32082 = n35508 ^ n35509;
  assign n35522 = n35543 & n35544;
  assign n33722 = n35183 ^ n35184;
  assign n35185 = ~n35184;
  assign n35228 = n35188 & n32;
  assign n35225 = ~n35256;
  assign n35227 = ~n35188;
  assign n35177 = n33768 ^ n33732;
  assign n35267 = ~n35295;
  assign n35301 = n31473 & n35328;
  assign n33790 = ~n35329;
  assign n35330 = n35368 & n35369;
  assign n35289 = ~n35376;
  assign n35347 = n468 ^ n35389;
  assign n35411 = n35427 & n35428;
  assign n35351 = n35429 ^ n35430;
  assign n35450 = n35470 & n35471;
  assign n35355 = n35472 ^ n32082;
  assign n32111 = ~n32082;
  assign n35510 = ~n35522;
  assign n35146 = ~n33722;
  assign n35102 = n35185 & n35186;
  assign n35187 = n35225 & n35226;
  assign n35214 = n35227 & n12118;
  assign n35150 = ~n35228;
  assign n35250 = n35177 & n35257;
  assign n35258 = n35267 & n35268;
  assign n35251 = ~n35177;
  assign n33809 = ~n35301;
  assign n35287 = n35330 ^ n32564;
  assign n35331 = ~n35330;
  assign n35209 = n35346 ^ n35347;
  assign n35348 = ~n35347;
  assign n35393 = n35351 & n467;
  assign n35390 = ~n35411;
  assign n35392 = ~n35351;
  assign n35435 = n35355 & n35395;
  assign n35431 = ~n35450;
  assign n35433 = ~n35355;
  assign n35473 = n35510 & n35511;
  assign n35105 = ~n35102;
  assign n35148 = n35187 ^ n35188;
  assign n35190 = ~n35187;
  assign n35189 = ~n35214;
  assign n35215 = ~n35250;
  assign n35229 = n35251 & n35217;
  assign n35216 = ~n35258;
  assign n31418 = n35286 ^ n35287;
  assign n35310 = n35331 & n35332;
  assign n35312 = n35209 & n32523;
  assign n35311 = ~n35209;
  assign n35269 = n35348 & n35349;
  assign n35350 = n35390 & n35391;
  assign n35377 = n35392 & n17816;
  assign n35315 = ~n35393;
  assign n35394 = n35431 & n35432;
  assign n35412 = n35433 & n35434;
  assign n35397 = ~n35435;
  assign n35437 = n35473 ^ n33194;
  assign n35474 = ~n35473;
  assign n35103 = n32 ^ n35148;
  assign n35175 = n35189 & n35190;
  assign n35208 = n35215 & n35216;
  assign n35176 = n35216 ^ n35217;
  assign n35179 = ~n35229;
  assign n33736 = n32564 ^ n31418;
  assign n35249 = n31418 & n35255;
  assign n31484 = ~n31418;
  assign n35288 = ~n35310;
  assign n35296 = n35311 & n32504;
  assign n35212 = ~n35312;
  assign n35313 = n35350 ^ n35351;
  assign n35352 = ~n35350;
  assign n35353 = ~n35377;
  assign n35354 = n35394 ^ n35395;
  assign n35396 = ~n35394;
  assign n35357 = ~n35412;
  assign n32069 = n35436 ^ n35437;
  assign n35451 = n35474 & n35475;
  assign n33687 = n35102 ^ n35103;
  assign n35104 = ~n35103;
  assign n35149 = ~n35175;
  assign n35107 = n35176 ^ n35177;
  assign n35178 = ~n35208;
  assign n35097 = n33736 ^ n33730;
  assign n33756 = ~n35249;
  assign n35223 = n31484 & n33771;
  assign n35252 = n35288 & n35289;
  assign n35254 = ~n35296;
  assign n35270 = n467 ^ n35313;
  assign n35336 = n35352 & n35353;
  assign n35273 = n35354 ^ n35355;
  assign n35378 = n35396 & n35397;
  assign n35277 = n35398 ^ n32069;
  assign n32027 = ~n32069;
  assign n35438 = ~n35451;
  assign n35067 = ~n33687;
  assign n35031 = n35104 & n35105;
  assign n35106 = n35149 & n35150;
  assign n35137 = n35107 & n12057;
  assign n35138 = ~n35107;
  assign n35139 = n35178 & n35179;
  assign n35170 = n35097 & n35180;
  assign n35169 = ~n35097;
  assign n33773 = ~n35223;
  assign n35210 = n35252 ^ n32504;
  assign n35253 = ~n35252;
  assign n35132 = n35269 ^ n35270;
  assign n35271 = ~n35270;
  assign n35316 = n35273 & n17747;
  assign n35314 = ~n35336;
  assign n35317 = ~n35273;
  assign n35360 = n35277 & n35319;
  assign n35356 = ~n35378;
  assign n35358 = ~n35277;
  assign n35399 = n35438 & n35439;
  assign n35069 = n35106 ^ n35107;
  assign n35108 = ~n35106;
  assign n35109 = ~n35137;
  assign n35128 = n35138 & n47;
  assign n35096 = n35139 ^ n35140;
  assign n35129 = ~n35139;
  assign n35151 = n35169 & n35140;
  assign n35089 = ~n35170;
  assign n31427 = n35209 ^ n35210;
  assign n35230 = n35253 & n35254;
  assign n35232 = n35132 & n32473;
  assign n35231 = ~n35132;
  assign n35191 = n35271 & n35269;
  assign n35272 = n35314 & n35315;
  assign n35275 = ~n35316;
  assign n35297 = n35317 & n466;
  assign n35318 = n35356 & n35357;
  assign n35337 = n35358 & n35359;
  assign n35321 = ~n35360;
  assign n35361 = n35399 ^ n33155;
  assign n35400 = ~n35399;
  assign n35032 = n47 ^ n35069;
  assign n35028 = n35096 ^ n35097;
  assign n35098 = n35108 & n35109;
  assign n35071 = ~n35128;
  assign n35136 = n31427 & n35146;
  assign n35130 = ~n35151;
  assign n33703 = n32523 ^ n31427;
  assign n31370 = ~n31427;
  assign n35211 = ~n35230;
  assign n35218 = n35231 & n32468;
  assign n35173 = ~n35232;
  assign n35194 = ~n35191;
  assign n35233 = n35272 ^ n35273;
  assign n35274 = ~n35272;
  assign n35235 = ~n35297;
  assign n35276 = n35318 ^ n35319;
  assign n35320 = ~n35318;
  assign n35279 = ~n35337;
  assign n31968 = n35361 ^ n35362;
  assign n35379 = n35400 & n35401;
  assign n33651 = n35031 ^ n35032;
  assign n34944 = n35032 & n35031;
  assign n35061 = n35028 & n46;
  assign n35060 = ~n35028;
  assign n35070 = ~n35098;
  assign n35110 = n35129 & n35130;
  assign n35019 = n33703 ^ n33695;
  assign n33725 = ~n35136;
  assign n35147 = n31370 & n33722;
  assign n35171 = n35211 & n35212;
  assign n35134 = ~n35218;
  assign n35192 = n466 ^ n35233;
  assign n35259 = n35274 & n35275;
  assign n35196 = n35276 ^ n35277;
  assign n35298 = n35320 & n35321;
  assign n35200 = n35322 ^ n31968;
  assign n35324 = n31968 & n34386;
  assign n32007 = ~n31968;
  assign n35363 = ~n35379;
  assign n34995 = ~n33651;
  assign n34947 = ~n34944;
  assign n35050 = n35060 & n12021;
  assign n34986 = ~n35061;
  assign n35062 = n35070 & n35071;
  assign n35090 = n35019 & n35099;
  assign n35088 = ~n35110;
  assign n35091 = ~n35019;
  assign n33741 = ~n35147;
  assign n35131 = n35171 ^ n32473;
  assign n35172 = ~n35171;
  assign n35174 = n35191 ^ n35192;
  assign n35193 = ~n35192;
  assign n35236 = n35196 & n17696;
  assign n35234 = ~n35259;
  assign n35237 = ~n35196;
  assign n35280 = n35200 & n35290;
  assign n35278 = ~n35298;
  assign n35281 = ~n35200;
  assign n35299 = n32007 & n35323;
  assign n34388 = ~n35324;
  assign n35325 = n35363 & n35364;
  assign n35026 = ~n35050;
  assign n35027 = ~n35062;
  assign n35051 = n35088 & n35089;
  assign n35021 = ~n35090;
  assign n35072 = n35091 & n35052;
  assign n31330 = n35131 ^ n35132;
  assign n35152 = n35172 & n35173;
  assign n35153 = n35174 & n32423;
  assign n35056 = ~n35174;
  assign n35111 = n35193 & n35194;
  assign n35195 = n35234 & n35235;
  assign n35198 = ~n35236;
  assign n35219 = n35237 & n465;
  assign n35238 = n35278 & n35279;
  assign n35202 = ~n35280;
  assign n35260 = n35281 & n35239;
  assign n34406 = ~n35299;
  assign n35282 = n35325 ^ n33098;
  assign n35326 = ~n35325;
  assign n35017 = n35026 & n35027;
  assign n34984 = n35027 ^ n35028;
  assign n35018 = n35051 ^ n35052;
  assign n35059 = n31330 & n35067;
  assign n35053 = ~n35051;
  assign n35054 = ~n35072;
  assign n31373 = ~n31330;
  assign n35133 = ~n35152;
  assign n35094 = ~n35153;
  assign n35141 = n35056 & n32444;
  assign n35154 = n35195 ^ n35196;
  assign n35197 = ~n35195;
  assign n35156 = ~n35219;
  assign n35199 = n35238 ^ n35239;
  assign n35240 = ~n35238;
  assign n35241 = ~n35260;
  assign n31868 = n35282 ^ n35283;
  assign n35300 = n35326 & n35327;
  assign n34945 = n46 ^ n34984;
  assign n34985 = ~n35017;
  assign n34949 = n35018 ^ n35019;
  assign n35033 = n35053 & n35054;
  assign n33706 = ~n35059;
  assign n33666 = n31373 ^ n32468;
  assign n35068 = n31373 & n33687;
  assign n35092 = n35133 & n35134;
  assign n35058 = ~n35141;
  assign n35112 = n465 ^ n35154;
  assign n35181 = n35197 & n35198;
  assign n35115 = n35199 ^ n35200;
  assign n35220 = n35240 & n35241;
  assign n35160 = n35242 ^ n31868;
  assign n35243 = n31868 & n34350;
  assign n31983 = ~n31868;
  assign n35284 = ~n35300;
  assign n33613 = n34944 ^ n34945;
  assign n34946 = ~n34945;
  assign n34948 = n34985 & n34986;
  assign n34975 = n34949 & n45;
  assign n34974 = ~n34949;
  assign n35020 = ~n35033;
  assign n34938 = n33666 ^ n33623;
  assign n33690 = ~n35068;
  assign n35055 = n35092 ^ n32423;
  assign n35093 = ~n35092;
  assign n34981 = n35111 ^ n35112;
  assign n35113 = ~n35112;
  assign n35158 = n35115 & n464;
  assign n35155 = ~n35181;
  assign n35157 = ~n35115;
  assign n35203 = n35160 & n35213;
  assign n35201 = ~n35220;
  assign n35204 = ~n35160;
  assign n34352 = ~n35243;
  assign n35221 = n31983 & n35244;
  assign n35245 = n35284 & n35285;
  assign n34906 = ~n33613;
  assign n34866 = n34946 & n34947;
  assign n34908 = n34948 ^ n34949;
  assign n34936 = ~n34948;
  assign n34955 = n34974 & n11976;
  assign n34898 = ~n34975;
  assign n34976 = n35020 & n35021;
  assign n34996 = n34938 & n34977;
  assign n34997 = ~n34938;
  assign n31289 = n35055 ^ n35056;
  assign n35073 = n35093 & n35094;
  assign n35034 = n35113 & n35111;
  assign n35114 = n35155 & n35156;
  assign n35142 = n35157 & n17666;
  assign n35076 = ~n35158;
  assign n35159 = n35201 & n35202;
  assign n35162 = ~n35203;
  assign n35182 = n35204 & n35119;
  assign n34372 = ~n35221;
  assign n35205 = n35245 ^ n35246;
  assign n35247 = ~n35245;
  assign n34867 = n45 ^ n34908;
  assign n34869 = ~n34866;
  assign n34935 = ~n34955;
  assign n34937 = n34976 ^ n34977;
  assign n34978 = ~n34976;
  assign n34979 = ~n34996;
  assign n34987 = n34997 & n34998;
  assign n34994 = n31289 & n33651;
  assign n33629 = n32444 ^ n31289;
  assign n31322 = ~n31289;
  assign n35057 = ~n35073;
  assign n35074 = n35114 ^ n35115;
  assign n35116 = ~n35114;
  assign n35117 = ~n35142;
  assign n35118 = n35159 ^ n35160;
  assign n35161 = ~n35159;
  assign n35121 = ~n35182;
  assign n31800 = n35205 ^ n33047;
  assign n35222 = n35247 & n35248;
  assign n33575 = n34866 ^ n34867;
  assign n34868 = ~n34867;
  assign n34918 = n34935 & n34936;
  assign n34854 = n34937 ^ n34938;
  assign n34956 = n34978 & n34979;
  assign n34858 = n33629 ^ n33621;
  assign n34940 = ~n34987;
  assign n33653 = ~n34994;
  assign n34983 = n31322 & n34995;
  assign n35022 = n35057 & n35058;
  assign n35035 = n464 ^ n35074;
  assign n35100 = n35116 & n35117;
  assign n35002 = n35118 ^ n35119;
  assign n35143 = n35161 & n35162;
  assign n35080 = n35163 ^ n31800;
  assign n35165 = n31800 & n34335;
  assign n31942 = ~n31800;
  assign n35206 = ~n35222;
  assign n34826 = ~n33575;
  assign n34773 = n34868 & n34869;
  assign n34899 = n34854 & n11934;
  assign n34897 = ~n34918;
  assign n34900 = ~n34854;
  assign n34942 = n34858 & n34950;
  assign n34939 = ~n34956;
  assign n34941 = ~n34858;
  assign n33669 = ~n34983;
  assign n34980 = n35022 ^ n32391;
  assign n35025 = n35022 & n32391;
  assign n35023 = ~n35022;
  assign n35024 = n35034 ^ n35035;
  assign n34957 = n35035 & n35034;
  assign n35078 = n35002 & n479;
  assign n35075 = ~n35100;
  assign n35077 = ~n35002;
  assign n35123 = n35080 & n35135;
  assign n35120 = ~n35143;
  assign n35122 = ~n35080;
  assign n35144 = n31942 & n35164;
  assign n34317 = ~n35165;
  assign n35166 = n35206 & n35207;
  assign n34776 = ~n34773;
  assign n34853 = n34897 & n34898;
  assign n34855 = ~n34899;
  assign n34877 = n34900 & n44;
  assign n34901 = n34939 & n34940;
  assign n34919 = n34941 & n34902;
  assign n34860 = ~n34942;
  assign n31292 = n34980 ^ n34981;
  assign n34999 = n35023 & n32420;
  assign n35000 = n35024 & n32374;
  assign n34988 = ~n35025;
  assign n34870 = ~n35024;
  assign n35036 = n35075 & n35076;
  assign n35063 = n35077 & n17570;
  assign n35004 = ~n35078;
  assign n35079 = n35120 & n35121;
  assign n35101 = n35122 & n35040;
  assign n35082 = ~n35123;
  assign n34337 = ~n35144;
  assign n35125 = n35166 ^ n33069;
  assign n35167 = ~n35166;
  assign n34814 = n34853 ^ n34854;
  assign n34856 = ~n34853;
  assign n34816 = ~n34877;
  assign n34857 = n34901 ^ n34902;
  assign n34896 = n31292 & n34906;
  assign n34903 = ~n34901;
  assign n34904 = ~n34919;
  assign n33591 = n32420 ^ n31292;
  assign n31248 = ~n31292;
  assign n34982 = n34988 & n34981;
  assign n34952 = ~n34999;
  assign n34911 = ~n35000;
  assign n34989 = n34870 & n32355;
  assign n35001 = n479 ^ n35036;
  assign n35037 = ~n35036;
  assign n35038 = ~n35063;
  assign n35039 = n35079 ^ n35080;
  assign n35081 = ~n35079;
  assign n35042 = ~n35101;
  assign n31728 = n35124 ^ n35125;
  assign n35145 = n35167 & n35168;
  assign n34774 = n44 ^ n34814;
  assign n34836 = n34855 & n34856;
  assign n34778 = n34857 ^ n34858;
  assign n33615 = ~n34896;
  assign n34878 = n34903 & n34904;
  assign n34782 = n33591 ^ n33547;
  assign n34907 = n31248 & n33613;
  assign n34951 = ~n34982;
  assign n34873 = ~n34989;
  assign n34958 = n35001 ^ n35002;
  assign n35029 = n35037 & n35038;
  assign n34960 = n35039 ^ n35040;
  assign n35064 = n35081 & n35082;
  assign n35008 = n35083 ^ n31728;
  assign n35084 = n31728 & n35095;
  assign n31816 = ~n31728;
  assign n35126 = ~n35145;
  assign n33537 = n34773 ^ n34774;
  assign n34775 = ~n34774;
  assign n34818 = n34778 & n43;
  assign n34815 = ~n34836;
  assign n34817 = ~n34778;
  assign n34861 = n34782 & n34820;
  assign n34859 = ~n34878;
  assign n34862 = ~n34782;
  assign n33633 = ~n34907;
  assign n34909 = n34951 & n34952;
  assign n34943 = n34957 ^ n34958;
  assign n34879 = n34958 & n34957;
  assign n35006 = n34960 & n478;
  assign n35003 = ~n35029;
  assign n35005 = ~n34960;
  assign n35043 = n35008 & n34964;
  assign n35041 = ~n35064;
  assign n35044 = ~n35008;
  assign n34276 = ~n35084;
  assign n35065 = n31816 & n34273;
  assign n35085 = n35126 & n35127;
  assign n34737 = ~n33537;
  assign n34703 = n34775 & n34776;
  assign n34777 = n34815 & n34816;
  assign n34794 = n34817 & n11895;
  assign n34741 = ~n34818;
  assign n34819 = n34859 & n34860;
  assign n34822 = ~n34861;
  assign n34837 = n34862 & n34863;
  assign n34871 = n34909 ^ n32355;
  assign n34910 = ~n34909;
  assign n34920 = n34943 & n32317;
  assign n34787 = ~n34943;
  assign n34882 = ~n34879;
  assign n34959 = n35003 & n35004;
  assign n34990 = n35005 & n17477;
  assign n34923 = ~n35006;
  assign n35007 = n35041 & n35042;
  assign n35010 = ~n35043;
  assign n35030 = n35044 & n35045;
  assign n34299 = ~n35065;
  assign n35047 = n35085 ^ n32974;
  assign n35086 = ~n35085;
  assign n34706 = ~n34703;
  assign n34739 = n34777 ^ n34778;
  assign n34780 = ~n34777;
  assign n34779 = ~n34794;
  assign n34781 = n34819 ^ n34820;
  assign n34821 = ~n34819;
  assign n34784 = ~n34837;
  assign n31203 = n34870 ^ n34871;
  assign n34905 = n34910 & n34911;
  assign n34829 = ~n34920;
  assign n34912 = n34787 & n32342;
  assign n34921 = n34959 ^ n34960;
  assign n34961 = ~n34959;
  assign n34962 = ~n34990;
  assign n34963 = n35007 ^ n35008;
  assign n35009 = ~n35007;
  assign n34966 = ~n35030;
  assign n31747 = n35046 ^ n35047;
  assign n35066 = n35086 & n35087;
  assign n34704 = n43 ^ n34739;
  assign n34761 = n34779 & n34780;
  assign n34708 = n34781 ^ n34782;
  assign n34795 = n34821 & n34822;
  assign n34812 = n31203 & n34826;
  assign n33553 = n31203 ^ n32355;
  assign n31251 = ~n31203;
  assign n34872 = ~n34905;
  assign n34789 = ~n34912;
  assign n34880 = n478 ^ n34921;
  assign n34953 = n34961 & n34962;
  assign n34884 = n34963 ^ n34964;
  assign n34991 = n35009 & n35010;
  assign n34888 = n35011 ^ n31747;
  assign n35012 = n31747 & n34242;
  assign n31698 = ~n31747;
  assign n35048 = ~n35066;
  assign n34679 = n34703 ^ n34704;
  assign n34705 = ~n34704;
  assign n34742 = n34708 & n11867;
  assign n34740 = ~n34761;
  assign n34743 = ~n34708;
  assign n34696 = n33553 ^ n33507;
  assign n34783 = ~n34795;
  assign n33595 = ~n34812;
  assign n34813 = n31251 & n33575;
  assign n34827 = n34872 & n34873;
  assign n34864 = n34879 ^ n34880;
  assign n34881 = ~n34880;
  assign n34924 = n34884 & n17431;
  assign n34922 = ~n34953;
  assign n34925 = ~n34884;
  assign n34969 = n34888 & n34927;
  assign n34965 = ~n34991;
  assign n34967 = ~n34888;
  assign n34244 = ~n35012;
  assign n34992 = n31698 & n35013;
  assign n35014 = n35048 & n35049;
  assign n34670 = ~n34679;
  assign n34635 = n34705 & n34706;
  assign n34707 = n34740 & n34741;
  assign n34710 = ~n34742;
  assign n34723 = n34743 & n42;
  assign n34747 = n34696 & n34724;
  assign n34762 = n34783 & n34784;
  assign n34748 = ~n34696;
  assign n33578 = ~n34813;
  assign n34786 = n34827 ^ n32317;
  assign n34828 = ~n34827;
  assign n34839 = n34864 & n32262;
  assign n34838 = ~n34864;
  assign n34796 = n34881 & n34882;
  assign n34883 = n34922 & n34923;
  assign n34886 = ~n34924;
  assign n34913 = n34925 & n477;
  assign n34926 = n34965 & n34966;
  assign n34954 = n34967 & n34968;
  assign n34890 = ~n34969;
  assign n34260 = ~n34992;
  assign n34970 = n35014 ^ n32918;
  assign n35015 = ~n35014;
  assign n34638 = ~n34635;
  assign n34672 = n34707 ^ n34708;
  assign n34709 = ~n34707;
  assign n34674 = ~n34723;
  assign n34681 = ~n34747;
  assign n34744 = n34748 & n34749;
  assign n34713 = ~n34762;
  assign n31193 = n34786 ^ n34787;
  assign n34823 = n34828 & n34829;
  assign n34830 = n34838 & n32328;
  assign n34715 = ~n34839;
  assign n34799 = ~n34796;
  assign n34840 = n34883 ^ n34884;
  assign n34885 = ~n34883;
  assign n34842 = ~n34913;
  assign n34887 = n34926 ^ n34927;
  assign n34928 = ~n34926;
  assign n34929 = ~n34954;
  assign n31628 = n34970 ^ n34971;
  assign n34993 = n35015 & n35016;
  assign n34636 = n42 ^ n34672;
  assign n34694 = n34709 & n34710;
  assign n34695 = n34713 ^ n34724;
  assign n34722 = n31193 & n34737;
  assign n34712 = ~n34744;
  assign n33514 = n32342 ^ n31193;
  assign n31153 = ~n31193;
  assign n34788 = ~n34823;
  assign n34753 = ~n34830;
  assign n34797 = n477 ^ n34840;
  assign n34874 = n34885 & n34886;
  assign n34801 = n34887 ^ n34888;
  assign n34914 = n34928 & n34929;
  assign n34930 = n31628 & n34224;
  assign n31667 = ~n31628;
  assign n34972 = ~n34993;
  assign n33473 = n34635 ^ n34636;
  assign n34637 = ~n34636;
  assign n34673 = ~n34694;
  assign n34640 = n34695 ^ n34696;
  assign n34711 = n34712 & n34713;
  assign n34614 = n33514 ^ n33505;
  assign n33540 = ~n34722;
  assign n34738 = n31153 & n33537;
  assign n34751 = n34788 & n34789;
  assign n34750 = n34753 & n34715;
  assign n34685 = n34796 ^ n34797;
  assign n34798 = ~n34797;
  assign n34843 = n34801 & n17352;
  assign n34841 = ~n34874;
  assign n34844 = ~n34801;
  assign n34889 = ~n34914;
  assign n34805 = n34915 ^ n31667;
  assign n34226 = ~n34930;
  assign n34916 = n31667 & n34931;
  assign n34932 = n34972 & n34973;
  assign n34607 = ~n33473;
  assign n34581 = n34637 & n34638;
  assign n34639 = n34673 & n34674;
  assign n34662 = n34640 & n41;
  assign n34661 = ~n34640;
  assign n34683 = n34614 & n34697;
  assign n34680 = ~n34711;
  assign n34682 = ~n34614;
  assign n33557 = ~n34738;
  assign n31077 = n34750 ^ n34751;
  assign n34752 = ~n34751;
  assign n34764 = n34685 & n32311;
  assign n34763 = ~n34685;
  assign n34725 = n34798 & n34799;
  assign n34800 = n34841 & n34842;
  assign n34803 = ~n34843;
  assign n34831 = n34844 & n476;
  assign n34845 = n34889 & n34890;
  assign n34875 = n34805 & n34891;
  assign n34876 = ~n34805;
  assign n34205 = ~n34916;
  assign n34892 = n34932 ^ n32905;
  assign n34933 = ~n34932;
  assign n34609 = n34639 ^ n34640;
  assign n34631 = ~n34639;
  assign n34645 = n34661 & n11822;
  assign n34603 = ~n34662;
  assign n34660 = n31077 & n34670;
  assign n34646 = n34680 & n34681;
  assign n34675 = n34682 & n34647;
  assign n34617 = ~n34683;
  assign n33495 = n31077 ^ n32262;
  assign n31169 = ~n31077;
  assign n34745 = n34752 & n34753;
  assign n34754 = n34763 & n32222;
  assign n34687 = ~n34764;
  assign n34765 = n34800 ^ n34801;
  assign n34802 = ~n34800;
  assign n34767 = ~n34831;
  assign n34804 = n34845 ^ n34846;
  assign n34832 = ~n34845;
  assign n34792 = ~n34875;
  assign n34865 = n34876 & n34846;
  assign n31599 = n34892 ^ n34893;
  assign n34917 = n34933 & n34934;
  assign n34582 = n41 ^ n34609;
  assign n34632 = ~n34645;
  assign n34613 = n34646 ^ n34647;
  assign n33520 = ~n34660;
  assign n34648 = ~n34646;
  assign n34649 = ~n34675;
  assign n34671 = n31169 & n34679;
  assign n34568 = n33495 ^ n33488;
  assign n34714 = ~n34745;
  assign n34653 = ~n34754;
  assign n34726 = n476 ^ n34765;
  assign n34790 = n34802 & n34803;
  assign n34729 = n34804 ^ n34805;
  assign n34718 = n34847 ^ n31599;
  assign n34833 = ~n34865;
  assign n34849 = n31599 & n34161;
  assign n31563 = ~n31599;
  assign n34894 = ~n34917;
  assign n33421 = n34581 ^ n34582;
  assign n34534 = n34582 & n34581;
  assign n34576 = n34613 ^ n34614;
  assign n34615 = n34631 & n34632;
  assign n34641 = n34648 & n34649;
  assign n34650 = n34568 & n34663;
  assign n33499 = ~n34671;
  assign n34651 = ~n34568;
  assign n34684 = n34714 & n34715;
  assign n34592 = n34725 ^ n34726;
  assign n34727 = ~n34726;
  assign n34769 = n34729 & n475;
  assign n34766 = ~n34790;
  assign n34768 = ~n34729;
  assign n34807 = n34718 & n34824;
  assign n34825 = n34832 & n34833;
  assign n34806 = ~n34718;
  assign n34834 = n31563 & n34848;
  assign n34163 = ~n34849;
  assign n34850 = n34894 & n34895;
  assign n34562 = ~n33421;
  assign n34587 = n34576 & n40;
  assign n34586 = ~n34576;
  assign n34602 = ~n34615;
  assign n34630 = n33520 & n33499;
  assign n34616 = ~n34641;
  assign n34570 = ~n34650;
  assign n34642 = n34651 & n34589;
  assign n33436 = n34684 ^ n34685;
  assign n34686 = ~n34684;
  assign n34664 = n34727 & n34725;
  assign n34728 = n34766 & n34767;
  assign n34755 = n34768 & n17233;
  assign n34700 = ~n34769;
  assign n34793 = n34806 & n34757;
  assign n34720 = ~n34807;
  assign n34791 = ~n34825;
  assign n34188 = ~n34834;
  assign n34809 = n34850 ^ n32855;
  assign n34851 = ~n34850;
  assign n34583 = n34586 & n11752;
  assign n34544 = ~n34587;
  assign n34575 = n34602 & n34603;
  assign n34588 = n34616 & n34617;
  assign n33518 = ~n34630;
  assign n34591 = ~n34642;
  assign n34548 = n33436 ^ n33371;
  assign n31011 = n33436 ^ n32222;
  assign n34676 = n34686 & n34687;
  assign n34698 = n34728 ^ n34729;
  assign n34730 = ~n34728;
  assign n34731 = ~n34755;
  assign n34756 = n34791 & n34792;
  assign n34759 = ~n34793;
  assign n31496 = n34808 ^ n34809;
  assign n34835 = n34851 & n34852;
  assign n34558 = n34575 ^ n34576;
  assign n34565 = ~n34583;
  assign n34566 = ~n34575;
  assign n34567 = n34588 ^ n34589;
  assign n34601 = n31011 & n34607;
  assign n34590 = ~n34588;
  assign n34620 = n34548 & n34525;
  assign n34618 = ~n34548;
  assign n31111 = ~n31011;
  assign n34652 = ~n34676;
  assign n34665 = n475 ^ n34698;
  assign n34716 = n34730 & n34731;
  assign n34717 = n34756 ^ n34757;
  assign n34657 = n34770 ^ n31496;
  assign n34758 = ~n34756;
  assign n34771 = n31496 & n34785;
  assign n31538 = ~n31496;
  assign n34810 = ~n34835;
  assign n34535 = n40 ^ n34558;
  assign n34564 = n34565 & n34566;
  assign n34502 = n34567 ^ n34568;
  assign n34584 = n34590 & n34591;
  assign n33456 = ~n34601;
  assign n34608 = n31111 & n33473;
  assign n34610 = n34618 & n34619;
  assign n34527 = ~n34620;
  assign n34621 = n34652 & n34653;
  assign n34643 = n34664 ^ n34665;
  assign n34605 = n34665 & n34664;
  assign n34699 = ~n34716;
  assign n34667 = n34717 ^ n34718;
  assign n34734 = n34657 & n34691;
  assign n34746 = n34758 & n34759;
  assign n34732 = ~n34657;
  assign n34129 = ~n34771;
  assign n34760 = n31538 & n34143;
  assign n34772 = n34810 & n34811;
  assign n33379 = n34534 ^ n34535;
  assign n34480 = n34535 & n34534;
  assign n34546 = n34502 & n55;
  assign n34543 = ~n34564;
  assign n34545 = ~n34502;
  assign n34569 = ~n34584;
  assign n33475 = ~n34608;
  assign n34550 = ~n34610;
  assign n34593 = n34621 ^ n32237;
  assign n34623 = n34621 & n32237;
  assign n34622 = ~n34621;
  assign n34633 = n34643 & n32172;
  assign n34538 = ~n34643;
  assign n34666 = n34699 & n34700;
  assign n34689 = n34667 & n474;
  assign n34688 = ~n34667;
  assign n34721 = n34732 & n34733;
  assign n34659 = ~n34734;
  assign n34719 = ~n34746;
  assign n34145 = ~n34760;
  assign n34736 = n34772 ^ n34074;
  assign n34514 = ~n33379;
  assign n34483 = ~n34480;
  assign n34521 = n34543 & n34544;
  assign n34541 = n34545 & n11714;
  assign n34504 = ~n34546;
  assign n34547 = n34569 & n34570;
  assign n30937 = n34592 ^ n34593;
  assign n34611 = n34622 & n32186;
  assign n34604 = ~n34623;
  assign n34624 = n34538 & n32194;
  assign n34561 = ~n34633;
  assign n34634 = n34666 ^ n34667;
  assign n34654 = ~n34666;
  assign n34677 = n34688 & n17168;
  assign n34626 = ~n34689;
  assign n34690 = n34719 & n34720;
  assign n34693 = ~n34721;
  assign n31503 = n34735 ^ n34736;
  assign n34501 = n55 ^ n34521;
  assign n34522 = ~n34521;
  assign n34523 = ~n34541;
  assign n34524 = n34547 ^ n34548;
  assign n34557 = n30937 & n34562;
  assign n34549 = ~n34547;
  assign n33396 = n30937 ^ n32186;
  assign n31048 = ~n30937;
  assign n34594 = n34604 & n34592;
  assign n34578 = ~n34611;
  assign n34540 = ~n34624;
  assign n34606 = n474 ^ n34634;
  assign n34655 = ~n34677;
  assign n34656 = n34690 ^ n34691;
  assign n34600 = n34701 ^ n31503;
  assign n34668 = n34702 ^ n31503;
  assign n34692 = ~n34690;
  assign n34090 = ~n31503;
  assign n34481 = n34501 ^ n34502;
  assign n34518 = n34522 & n34523;
  assign n34485 = n34524 ^ n34525;
  assign n34542 = n34549 & n34550;
  assign n34508 = n33396 ^ n33388;
  assign n33423 = ~n34557;
  assign n34563 = n31048 & n33421;
  assign n34577 = ~n34594;
  assign n34493 = n34605 ^ n34606;
  assign n34552 = n34606 & n34605;
  assign n34644 = n34654 & n34655;
  assign n34596 = n34656 ^ n34657;
  assign n34112 = n34668 ^ n34669;
  assign n34678 = n34692 & n34693;
  assign n33341 = n34480 ^ n34481;
  assign n34482 = ~n34481;
  assign n34505 = n34485 & n11658;
  assign n34503 = ~n34518;
  assign n34506 = ~n34485;
  assign n34529 = n34508 & n34536;
  assign n34526 = ~n34542;
  assign n34528 = ~n34508;
  assign n33441 = ~n34563;
  assign n34559 = n34577 & n34578;
  assign n34580 = n34493 & n32129;
  assign n34579 = ~n34493;
  assign n34627 = n34596 & n17141;
  assign n34625 = ~n34644;
  assign n34628 = ~n34596;
  assign n34658 = ~n34678;
  assign n34463 = ~n33341;
  assign n34445 = n34482 & n34483;
  assign n34484 = n34503 & n34504;
  assign n34487 = ~n34505;
  assign n34496 = n34506 & n54;
  assign n34507 = n34526 & n34527;
  assign n34519 = n34528 & n34489;
  assign n34509 = ~n34529;
  assign n34537 = n34559 ^ n32172;
  assign n34560 = ~n34559;
  assign n34571 = n34579 & n32162;
  assign n34517 = ~n34580;
  assign n34595 = n34625 & n34626;
  assign n34598 = ~n34627;
  assign n34612 = n34628 & n473;
  assign n34629 = n34658 & n34659;
  assign n34448 = ~n34445;
  assign n34465 = n34484 ^ n34485;
  assign n34486 = ~n34484;
  assign n34467 = ~n34496;
  assign n34488 = n34507 ^ n34508;
  assign n34510 = ~n34507;
  assign n34491 = ~n34519;
  assign n30979 = n34537 ^ n34538;
  assign n34551 = n34560 & n34561;
  assign n34495 = ~n34571;
  assign n34572 = n34595 ^ n34596;
  assign n34597 = ~n34595;
  assign n34574 = ~n34612;
  assign n34599 = n472 ^ n34629;
  assign n34446 = n54 ^ n34465;
  assign n34478 = n34486 & n34487;
  assign n34450 = n34488 ^ n34489;
  assign n34497 = n34509 & n34510;
  assign n34499 = n30979 & n34514;
  assign n33359 = n30979 ^ n32194;
  assign n30908 = ~n30979;
  assign n34539 = ~n34551;
  assign n34553 = n473 ^ n34572;
  assign n34585 = n34597 & n34598;
  assign n34556 = n34599 ^ n34600;
  assign n34436 = n34445 ^ n34446;
  assign n34447 = ~n34446;
  assign n34469 = n34450 & n53;
  assign n34466 = ~n34478;
  assign n34468 = ~n34450;
  assign n34443 = n33359 ^ n33351;
  assign n34490 = ~n34497;
  assign n33382 = ~n34499;
  assign n34500 = n30908 & n33379;
  assign n34515 = n34539 & n34540;
  assign n34456 = n34552 ^ n34553;
  assign n34554 = ~n34553;
  assign n34573 = ~n34585;
  assign n33303 = ~n34436;
  assign n34411 = n34447 & n34448;
  assign n34449 = n34466 & n34467;
  assign n34461 = n34468 & n11582;
  assign n34431 = ~n34469;
  assign n34472 = n34443 & n34462;
  assign n34479 = n34490 & n34491;
  assign n34473 = ~n34443;
  assign n33400 = ~n34500;
  assign n34492 = n34515 ^ n32129;
  assign n34516 = ~n34515;
  assign n34531 = n34456 & n32111;
  assign n34530 = ~n34456;
  assign n34532 = n34554 & n34552;
  assign n34555 = n34573 & n34574;
  assign n34429 = n34449 ^ n34450;
  assign n34451 = ~n34449;
  assign n34452 = ~n34461;
  assign n34438 = ~n34472;
  assign n34470 = n34473 & n34474;
  assign n34455 = ~n34479;
  assign n30839 = n34492 ^ n34493;
  assign n34511 = n34516 & n34517;
  assign n34520 = n34530 & n32082;
  assign n34459 = ~n34531;
  assign n34533 = n34555 ^ n34556;
  assign n34412 = n53 ^ n34429;
  assign n34442 = n34451 & n34452;
  assign n34444 = n34455 ^ n34462;
  assign n34460 = n30839 & n34463;
  assign n34454 = ~n34470;
  assign n30898 = ~n30839;
  assign n34494 = ~n34511;
  assign n34477 = ~n34520;
  assign n34421 = n34532 ^ n34533;
  assign n34398 = n34411 ^ n34412;
  assign n34375 = n34412 & n34411;
  assign n34430 = ~n34442;
  assign n34414 = n34443 ^ n34444;
  assign n34453 = n34454 & n34455;
  assign n33364 = ~n34460;
  assign n33318 = n30898 ^ n32162;
  assign n34464 = n30898 & n33341;
  assign n34475 = n34494 & n34495;
  assign n34513 = n34421 & n32069;
  assign n34512 = ~n34421;
  assign n33262 = ~n34398;
  assign n34413 = n34430 & n34431;
  assign n34426 = n34414 & n52;
  assign n34425 = ~n34414;
  assign n34437 = ~n34453;
  assign n34400 = n33318 ^ n33272;
  assign n33344 = ~n34464;
  assign n34457 = n34475 ^ n32082;
  assign n34476 = ~n34475;
  assign n34498 = n34512 & n32027;
  assign n34423 = ~n34513;
  assign n34393 = n34413 ^ n34414;
  assign n34408 = ~n34413;
  assign n34417 = n34425 & n11500;
  assign n34391 = ~n34426;
  assign n34418 = n34437 & n34438;
  assign n34432 = n34400 & n34419;
  assign n34433 = ~n34400;
  assign n30793 = n34456 ^ n34457;
  assign n34471 = n34476 & n34477;
  assign n34441 = ~n34498;
  assign n34376 = n52 ^ n34393;
  assign n34407 = ~n34417;
  assign n34399 = n34418 ^ n34419;
  assign n34424 = n30793 & n33303;
  assign n34416 = ~n34418;
  assign n34395 = ~n34432;
  assign n34427 = n34433 & n34434;
  assign n33278 = n30793 ^ n32111;
  assign n30768 = ~n30793;
  assign n34458 = ~n34471;
  assign n33224 = n34375 ^ n34376;
  assign n34329 = n34376 & n34375;
  assign n34366 = n34399 ^ n34400;
  assign n34401 = n34407 & n34408;
  assign n34359 = n33278 ^ n33270;
  assign n33305 = ~n34424;
  assign n34415 = ~n34427;
  assign n34428 = n30768 & n34436;
  assign n34439 = n34458 & n34459;
  assign n34356 = ~n33224;
  assign n34382 = n34366 & n11429;
  assign n34383 = ~n34366;
  assign n34390 = ~n34401;
  assign n34402 = n34359 & n34409;
  assign n34410 = n34415 & n34416;
  assign n34403 = ~n34359;
  assign n33322 = ~n34428;
  assign n34420 = n34439 ^ n32027;
  assign n34440 = ~n34439;
  assign n34373 = ~n34382;
  assign n34377 = n34383 & n51;
  assign n34384 = n34390 & n34391;
  assign n34361 = ~n34402;
  assign n34396 = n34403 & n34379;
  assign n34394 = ~n34410;
  assign n30743 = n34420 ^ n34421;
  assign n34435 = n34440 & n34441;
  assign n34355 = ~n34377;
  assign n34365 = ~n34384;
  assign n34389 = n30743 & n33262;
  assign n34378 = n34394 & n34395;
  assign n34381 = ~n34396;
  assign n33237 = n30743 ^ n32069;
  assign n30671 = ~n30743;
  assign n34422 = ~n34435;
  assign n34348 = n34365 ^ n34366;
  assign n34364 = n34373 & n34365;
  assign n34358 = n34378 ^ n34379;
  assign n34323 = n33237 ^ n33221;
  assign n33264 = ~n34389;
  assign n34380 = ~n34378;
  assign n34392 = n30671 & n34398;
  assign n34404 = n34422 & n34423;
  assign n34330 = n51 ^ n34348;
  assign n34339 = n34358 ^ n34359;
  assign n34354 = ~n34364;
  assign n34369 = n34323 & n34345;
  assign n34374 = n34380 & n34381;
  assign n34367 = ~n34323;
  assign n33283 = ~n34392;
  assign n34385 = n34404 ^ n32007;
  assign n34405 = ~n34404;
  assign n34318 = n34329 ^ n34330;
  assign n34300 = n34330 & n34329;
  assign n34343 = n34339 & n50;
  assign n34338 = n34354 & n34355;
  assign n34342 = ~n34339;
  assign n34362 = n34367 & n34368;
  assign n34326 = ~n34369;
  assign n34360 = ~n34374;
  assign n30660 = n34385 ^ n34386;
  assign n34397 = n34405 & n34406;
  assign n34315 = ~n34318;
  assign n34319 = n34338 ^ n34339;
  assign n34340 = n34342 & n11352;
  assign n34307 = ~n34343;
  assign n34322 = ~n34338;
  assign n34353 = n30660 & n34356;
  assign n34344 = n34360 & n34361;
  assign n34347 = ~n34362;
  assign n33201 = n30660 ^ n31968;
  assign n30597 = ~n30660;
  assign n34387 = ~n34397;
  assign n34301 = n50 ^ n34319;
  assign n34321 = ~n34340;
  assign n34324 = n34344 ^ n34345;
  assign n34286 = n33201 ^ n33192;
  assign n33227 = ~n34353;
  assign n34346 = ~n34344;
  assign n34357 = n30597 & n33224;
  assign n34370 = n34387 & n34388;
  assign n33145 = n34300 ^ n34301;
  assign n34246 = n34301 & n34300;
  assign n34320 = n34321 & n34322;
  assign n34282 = n34323 ^ n34324;
  assign n34331 = n34286 & n34311;
  assign n34341 = n34346 & n34347;
  assign n34332 = ~n34286;
  assign n33244 = ~n34357;
  assign n34349 = n34370 ^ n31983;
  assign n34371 = ~n34370;
  assign n34277 = ~n33145;
  assign n34257 = ~n34246;
  assign n34308 = n34282 & n11263;
  assign n34306 = ~n34320;
  assign n34309 = ~n34282;
  assign n34288 = ~n34331;
  assign n34327 = n34332 & n34333;
  assign n34325 = ~n34341;
  assign n30483 = n34349 ^ n34350;
  assign n34363 = n34371 & n34372;
  assign n34281 = n34306 & n34307;
  assign n34283 = ~n34308;
  assign n34302 = n34309 & n49;
  assign n34305 = n30483 & n34315;
  assign n34310 = n34325 & n34326;
  assign n34312 = ~n34327;
  assign n33177 = n31868 ^ n30483;
  assign n30595 = ~n30483;
  assign n34351 = ~n34363;
  assign n34263 = n34281 ^ n34282;
  assign n34284 = ~n34281;
  assign n34265 = ~n34302;
  assign n33186 = ~n34305;
  assign n34285 = n34310 ^ n34311;
  assign n34269 = n33163 ^ n33177;
  assign n34314 = n30595 & n34318;
  assign n34313 = ~n34310;
  assign n34334 = n34351 & n34352;
  assign n34247 = n49 ^ n34263;
  assign n34279 = n34283 & n34284;
  assign n34249 = n34285 ^ n34286;
  assign n34293 = n34269 & n34303;
  assign n34304 = n34312 & n34313;
  assign n34292 = ~n34269;
  assign n33207 = ~n34314;
  assign n33124 = n34334 ^ n34335;
  assign n34336 = ~n34334;
  assign n33127 = n34246 ^ n34247;
  assign n34208 = n34247 & n34257;
  assign n34266 = n34249 & n11173;
  assign n34264 = ~n34279;
  assign n34267 = ~n34249;
  assign n34280 = n33186 & n33207;
  assign n34289 = n34292 & n34253;
  assign n34271 = ~n34293;
  assign n34287 = ~n34304;
  assign n34238 = n33124 ^ n33047;
  assign n30411 = n33124 ^ n31942;
  assign n34328 = n34336 & n34337;
  assign n34231 = ~n33127;
  assign n34211 = ~n34208;
  assign n34248 = n34264 & n34265;
  assign n34250 = ~n34266;
  assign n34261 = n34267 & n48;
  assign n34272 = n30411 & n34277;
  assign n33205 = ~n34280;
  assign n34268 = n34287 & n34288;
  assign n34255 = ~n34289;
  assign n34294 = n34238 & n34216;
  assign n34295 = ~n34238;
  assign n30508 = ~n30411;
  assign n34316 = ~n34328;
  assign n34232 = n34248 ^ n34249;
  assign n34251 = ~n34248;
  assign n34234 = ~n34261;
  assign n34252 = n34268 ^ n34269;
  assign n33148 = ~n34272;
  assign n34270 = ~n34268;
  assign n34278 = n30508 & n33145;
  assign n34240 = ~n34294;
  assign n34290 = n34295 & n34296;
  assign n34297 = n34316 & n34317;
  assign n34209 = n48 ^ n34232;
  assign n34245 = n34250 & n34251;
  assign n34195 = n34252 ^ n34253;
  assign n34262 = n34270 & n34271;
  assign n33166 = ~n34278;
  assign n34218 = ~n34290;
  assign n34274 = n34297 ^ n31728;
  assign n34298 = ~n34297;
  assign n33058 = n34208 ^ n34209;
  assign n34210 = ~n34209;
  assign n34236 = n34195 & n63;
  assign n34233 = ~n34245;
  assign n34235 = ~n34195;
  assign n34254 = ~n34262;
  assign n30338 = n34273 ^ n34274;
  assign n34291 = n34298 & n34299;
  assign n34193 = ~n33058;
  assign n34165 = n34210 & n34211;
  assign n34227 = n30338 & n34231;
  assign n34212 = n34233 & n34234;
  assign n34228 = n34235 & n11134;
  assign n34197 = ~n34236;
  assign n34237 = n34254 & n34255;
  assign n30433 = ~n30338;
  assign n34275 = ~n34291;
  assign n34168 = ~n34165;
  assign n34194 = n63 ^ n34212;
  assign n33109 = ~n34227;
  assign n34213 = ~n34212;
  assign n34214 = ~n34228;
  assign n34215 = n34237 ^ n34238;
  assign n34230 = n30433 & n33127;
  assign n34239 = ~n34237;
  assign n33080 = n30433 ^ n31728;
  assign n34258 = n34275 & n34276;
  assign n34166 = n34194 ^ n34195;
  assign n34206 = n34213 & n34214;
  assign n34170 = n34215 ^ n34216;
  assign n33129 = ~n34230;
  assign n34229 = n34239 & n34240;
  assign n34201 = n33080 ^ n33069;
  assign n34241 = n34258 ^ n31698;
  assign n34259 = ~n34258;
  assign n33011 = n34165 ^ n34166;
  assign n34167 = ~n34166;
  assign n34198 = n34170 & n10999;
  assign n34196 = ~n34206;
  assign n34199 = ~n34170;
  assign n34219 = n34201 & n34174;
  assign n34217 = ~n34229;
  assign n34220 = ~n34201;
  assign n30373 = n34241 ^ n34242;
  assign n34256 = n34259 & n34260;
  assign n34149 = ~n33011;
  assign n34131 = n34167 & n34168;
  assign n34189 = n30373 & n34193;
  assign n34169 = n34196 & n34197;
  assign n34172 = ~n34198;
  assign n34190 = n34199 & n62;
  assign n34200 = n34217 & n34218;
  assign n34176 = ~n34219;
  assign n34207 = n34220 & n34221;
  assign n33034 = n31747 ^ n30373;
  assign n30302 = ~n30373;
  assign n34243 = ~n34256;
  assign n34151 = n34169 ^ n34170;
  assign n33060 = ~n34189;
  assign n34171 = ~n34169;
  assign n34153 = ~n34190;
  assign n34173 = n34200 ^ n34201;
  assign n34192 = n30302 & n33058;
  assign n34138 = n33034 ^ n32974;
  assign n34202 = ~n34200;
  assign n34203 = ~n34207;
  assign n34223 = n34243 & n34244;
  assign n34132 = n62 ^ n34151;
  assign n34164 = n34171 & n34172;
  assign n34134 = n34173 ^ n34174;
  assign n34182 = n34138 & n34157;
  assign n33084 = ~n34192;
  assign n34191 = n34202 & n34203;
  assign n34180 = ~n34138;
  assign n32984 = n34223 ^ n34224;
  assign n34225 = ~n34223;
  assign n32962 = n34131 ^ n34132;
  assign n34092 = n34132 & n34131;
  assign n34154 = n34134 & n10917;
  assign n34152 = ~n34164;
  assign n34155 = ~n34134;
  assign n34177 = n34180 & n34181;
  assign n34159 = ~n34182;
  assign n34175 = ~n34191;
  assign n34101 = n32984 ^ n32972;
  assign n30217 = n31628 ^ n32984;
  assign n34222 = n34225 & n34226;
  assign n34118 = ~n32962;
  assign n34095 = ~n34092;
  assign n34146 = n30217 & n34149;
  assign n34133 = n34152 & n34153;
  assign n34136 = ~n34154;
  assign n34147 = n34155 & n61;
  assign n34156 = n34175 & n34176;
  assign n34140 = ~n34177;
  assign n34183 = n34101 & n34125;
  assign n34184 = ~n34101;
  assign n30300 = ~n30217;
  assign n34204 = ~n34222;
  assign n34119 = n34133 ^ n34134;
  assign n33038 = ~n34146;
  assign n34135 = ~n34133;
  assign n34121 = ~n34147;
  assign n34137 = n34156 ^ n34157;
  assign n34150 = n30300 & n33011;
  assign n34158 = ~n34156;
  assign n34103 = ~n34183;
  assign n34178 = n34184 & n34185;
  assign n34186 = n34204 & n34205;
  assign n34093 = n61 ^ n34119;
  assign n34130 = n34135 & n34136;
  assign n34097 = n34137 ^ n34138;
  assign n33014 = ~n34150;
  assign n34148 = n34158 & n34159;
  assign n34127 = ~n34178;
  assign n34160 = n34186 ^ n31563;
  assign n34187 = ~n34186;
  assign n32907 = n34092 ^ n34093;
  assign n34094 = ~n34093;
  assign n34122 = n34097 & n10873;
  assign n34120 = ~n34130;
  assign n34123 = ~n34097;
  assign n34139 = ~n34148;
  assign n30215 = n34160 ^ n34161;
  assign n34179 = n34187 & n34188;
  assign n34079 = ~n32907;
  assign n34080 = n34094 & n34095;
  assign n34096 = n34120 & n34121;
  assign n34099 = ~n34122;
  assign n34114 = n34123 & n60;
  assign n34117 = n30215 & n32962;
  assign n34124 = n34139 & n34140;
  assign n32930 = n31599 ^ n30215;
  assign n30146 = ~n30215;
  assign n34162 = ~n34179;
  assign n34072 = ~n34080;
  assign n34081 = n34096 ^ n34097;
  assign n34098 = ~n34096;
  assign n34083 = ~n34114;
  assign n32964 = ~n34117;
  assign n34113 = n30146 & n34118;
  assign n34100 = n34124 ^ n34125;
  assign n34069 = n32930 ^ n32905;
  assign n34126 = ~n34124;
  assign n34142 = n34162 & n34163;
  assign n34063 = n60 ^ n34081;
  assign n34091 = n34098 & n34099;
  assign n34065 = n34100 ^ n34101;
  assign n32989 = ~n34113;
  assign n34108 = n34069 & n34087;
  assign n34115 = n34126 & n34127;
  assign n34106 = ~n34069;
  assign n32871 = n34142 ^ n34143;
  assign n34144 = ~n34142;
  assign n34039 = n34063 & n34072;
  assign n34084 = n34065 & n10788;
  assign n34082 = ~n34091;
  assign n34085 = ~n34065;
  assign n34104 = n34106 & n34107;
  assign n34089 = ~n34108;
  assign n34102 = ~n34115;
  assign n34046 = n32871 ^ n32855;
  assign n30129 = n32871 ^ n31496;
  assign n34141 = n34144 & n34145;
  assign n34075 = n30129 & n34079;
  assign n34064 = n34082 & n34083;
  assign n34067 = ~n34084;
  assign n34076 = n34085 & n59;
  assign n34086 = n34102 & n34103;
  assign n34071 = ~n34104;
  assign n34110 = n34046 & n34116;
  assign n34109 = ~n34046;
  assign n30078 = ~n30129;
  assign n34128 = ~n34141;
  assign n34051 = n34064 ^ n34065;
  assign n32949 = ~n34075;
  assign n34066 = ~n34064;
  assign n34053 = ~n34076;
  assign n34068 = n34086 ^ n34087;
  assign n34078 = n30078 & n32907;
  assign n34088 = ~n34086;
  assign n34105 = n34109 & n34057;
  assign n34048 = ~n34110;
  assign n34111 = n34128 & n34129;
  assign n34040 = n59 ^ n34051;
  assign n34061 = n34066 & n34067;
  assign n34042 = n34068 ^ n34069;
  assign n32922 = ~n34078;
  assign n34077 = n34088 & n34089;
  assign n34059 = ~n34105;
  assign n31540 = n34111 ^ n34112;
  assign n32164 = n34039 ^ n34040;
  assign n34019 = n34040 & n34039;
  assign n34054 = n34042 & n10703;
  assign n34052 = ~n34061;
  assign n34055 = ~n34042;
  assign n34070 = ~n34077;
  assign n34062 = n34080 ^ n31540;
  assign n34073 = n34090 ^ n31540;
  assign n33085 = n32164 ^ n33088;
  assign n34018 = n32164 ^ n34031;
  assign n33995 = n32164 & n32155;
  assign n34022 = ~n34019;
  assign n34041 = n34052 & n34053;
  assign n34043 = ~n34054;
  assign n34049 = n34055 & n58;
  assign n32891 = n34062 ^ n34063;
  assign n34056 = n34070 & n34071;
  assign n32860 = n34073 ^ n34074;
  assign n31268 = n33085 ^ n33110;
  assign n32525 = n135 ^ n34018;
  assign n33958 = n33085 & n34029;
  assign n33919 = n34018 & n135;
  assign n34032 = n34041 ^ n34042;
  assign n34044 = ~n34041;
  assign n34034 = ~n34049;
  assign n34045 = n34056 ^ n34057;
  assign n34028 = n32860 ^ n34060;
  assign n34058 = ~n34056;
  assign n32547 = ~n32525;
  assign n34020 = n58 ^ n34032;
  assign n34038 = n34043 & n34044;
  assign n34024 = n34045 ^ n34046;
  assign n34050 = n34058 & n34059;
  assign n34016 = n34019 ^ n34020;
  assign n34021 = ~n34020;
  assign n34036 = n34024 & n57;
  assign n34033 = ~n34038;
  assign n34035 = ~n34024;
  assign n34047 = ~n34050;
  assign n34012 = n34016 & n32133;
  assign n34011 = ~n34016;
  assign n34004 = n34021 & n34022;
  assign n34023 = n34033 & n34034;
  assign n34030 = n34035 & n10623;
  assign n34015 = ~n34036;
  assign n34037 = n34047 & n34048;
  assign n34010 = n34011 & n31985;
  assign n34003 = ~n34012;
  assign n34007 = ~n34004;
  assign n34013 = n34023 ^ n34024;
  assign n34025 = ~n34023;
  assign n34026 = ~n34030;
  assign n34027 = n56 ^ n34037;
  assign n34002 = n34003 & n33995;
  assign n34001 = ~n34010;
  assign n34005 = n57 ^ n34013;
  assign n34017 = n34025 & n34026;
  assign n34009 = n34027 ^ n34028;
  assign n34000 = ~n34002;
  assign n33994 = n34001 & n34003;
  assign n33984 = n34004 ^ n34005;
  assign n34006 = ~n34005;
  assign n34014 = ~n34017;
  assign n31086 = n33994 ^ n33995;
  assign n33992 = n34000 & n34001;
  assign n33996 = n33984 & n31956;
  assign n33997 = ~n33984;
  assign n33998 = n34006 & n34007;
  assign n34008 = n34014 & n34015;
  assign n33981 = n33987 ^ n31086;
  assign n33983 = n33992 ^ n31975;
  assign n31242 = ~n31086;
  assign n33988 = ~n33992;
  assign n33980 = ~n33996;
  assign n33993 = n33997 & n31975;
  assign n33999 = n34008 ^ n34009;
  assign n33976 = n33981 & n33982;
  assign n31060 = n33983 ^ n33984;
  assign n33977 = ~n33981;
  assign n33989 = ~n33993;
  assign n33962 = n33998 ^ n33999;
  assign n33945 = n33974 ^ n31060;
  assign n33960 = ~n33976;
  assign n33975 = n33977 & n33978;
  assign n31080 = ~n31060;
  assign n33985 = n33988 & n33989;
  assign n33991 = n33962 & n31910;
  assign n33990 = ~n33962;
  assign n33965 = n33945 & n33929;
  assign n33966 = ~n33945;
  assign n33970 = ~n33975;
  assign n33979 = ~n33985;
  assign n33986 = n33990 & n31874;
  assign n33964 = ~n33991;
  assign n33933 = ~n33965;
  assign n33956 = n33966 & n33967;
  assign n33968 = n33970 & n33958;
  assign n33957 = n33970 & n33960;
  assign n33971 = n33979 & n33980;
  assign n33973 = ~n33986;
  assign n33947 = ~n33956;
  assign n33954 = n33957 ^ n33958;
  assign n33959 = ~n33968;
  assign n33961 = n33971 ^ n31874;
  assign n33972 = ~n33971;
  assign n33949 = n33954 & n134;
  assign n33948 = ~n33954;
  assign n33955 = n33959 & n33960;
  assign n31017 = n33961 ^ n33962;
  assign n33969 = n33972 & n33973;
  assign n33943 = n33948 & n6633;
  assign n33923 = ~n33949;
  assign n33898 = n33950 ^ n31017;
  assign n33944 = ~n33955;
  assign n30981 = ~n31017;
  assign n33963 = ~n33969;
  assign n33935 = n33898 & n33941;
  assign n33934 = ~n33943;
  assign n33936 = ~n33898;
  assign n33928 = n33944 ^ n33945;
  assign n33942 = n33947 & n33944;
  assign n33951 = n33963 & n33964;
  assign n33896 = n33928 ^ n33929;
  assign n33930 = n33934 & n33919;
  assign n33918 = n33934 & n33923;
  assign n33902 = ~n33935;
  assign n33931 = n33936 & n33917;
  assign n33932 = ~n33942;
  assign n33937 = n33951 ^ n31784;
  assign n33952 = ~n33951;
  assign n33912 = n33896 & n133;
  assign n33900 = n33918 ^ n33919;
  assign n33911 = ~n33896;
  assign n33922 = ~n33930;
  assign n33921 = ~n33931;
  assign n33916 = n33932 & n33933;
  assign n30914 = n33937 ^ n33938;
  assign n33946 = n33952 & n33953;
  assign n32493 = n33900 ^ n32547;
  assign n33861 = n33900 & n32525;
  assign n33909 = n33911 & n6535;
  assign n33880 = ~n33912;
  assign n33899 = n33916 ^ n33917;
  assign n33914 = n33922 & n33923;
  assign n33867 = n33924 ^ n30914;
  assign n33920 = ~n33916;
  assign n30889 = ~n30914;
  assign n33939 = ~n33946;
  assign n33644 = ~n32493;
  assign n33858 = n33898 ^ n33899;
  assign n33894 = ~n33909;
  assign n33904 = n33867 & n33910;
  assign n33895 = ~n33914;
  assign n33903 = ~n33867;
  assign n33913 = n33920 & n33921;
  assign n33925 = n33939 & n33940;
  assign n33884 = n33858 & n132;
  assign n33883 = ~n33858;
  assign n33892 = n33894 & n33895;
  assign n33878 = n33895 ^ n33896;
  assign n33897 = n33903 & n33886;
  assign n33869 = ~n33904;
  assign n33901 = ~n33913;
  assign n33905 = n33925 ^ n31703;
  assign n33926 = ~n33925;
  assign n33862 = n133 ^ n33878;
  assign n33877 = n33883 & n6467;
  assign n33845 = ~n33884;
  assign n33879 = ~n33892;
  assign n33888 = ~n33897;
  assign n33885 = n33901 & n33902;
  assign n30860 = n33905 ^ n33906;
  assign n33915 = n33926 & n33927;
  assign n32460 = n33861 ^ n33862;
  assign n33821 = n33862 & n33861;
  assign n33863 = ~n33877;
  assign n33875 = n33879 & n33880;
  assign n33866 = n33885 ^ n33886;
  assign n33836 = n33889 ^ n30860;
  assign n33887 = ~n33885;
  assign n30797 = ~n30860;
  assign n33907 = ~n33915;
  assign n33606 = ~n32460;
  assign n33824 = ~n33821;
  assign n33831 = n33866 ^ n33867;
  assign n33857 = ~n33875;
  assign n33872 = n33836 & n33853;
  assign n33870 = ~n33836;
  assign n33881 = n33887 & n33888;
  assign n33893 = n33907 & n33908;
  assign n33851 = n33831 & n131;
  assign n33840 = n33857 ^ n33858;
  assign n33856 = n33863 & n33857;
  assign n33850 = ~n33831;
  assign n33864 = n33870 & n33871;
  assign n33838 = ~n33872;
  assign n33868 = ~n33881;
  assign n33891 = n33893 & n31605;
  assign n33890 = ~n33893;
  assign n33822 = n132 ^ n33840;
  assign n33846 = n33850 & n6372;
  assign n33812 = ~n33851;
  assign n33844 = ~n33856;
  assign n33855 = ~n33864;
  assign n33852 = n33868 & n33869;
  assign n33882 = n33890 & n31706;
  assign n33874 = ~n33891;
  assign n32428 = n33821 ^ n33822;
  assign n33823 = ~n33822;
  assign n33830 = n33844 & n33845;
  assign n33832 = ~n33846;
  assign n33835 = n33852 ^ n33853;
  assign n33854 = ~n33852;
  assign n33873 = n33874 & n33876;
  assign n33860 = ~n33882;
  assign n33568 = ~n32428;
  assign n33791 = n33823 & n33824;
  assign n33810 = n33830 ^ n33831;
  assign n33796 = n33835 ^ n33836;
  assign n33833 = ~n33830;
  assign n33847 = n33854 & n33855;
  assign n33859 = ~n33873;
  assign n33865 = n33860 & n33874;
  assign n33792 = n131 ^ n33810;
  assign n33794 = ~n33791;
  assign n33817 = n33796 & n6286;
  assign n33825 = n33832 & n33833;
  assign n33818 = ~n33796;
  assign n33837 = ~n33847;
  assign n33841 = n33859 & n33860;
  assign n33849 = ~n33865;
  assign n32396 = n33791 ^ n33792;
  assign n33793 = ~n33792;
  assign n33798 = ~n33817;
  assign n33813 = n33818 & n130;
  assign n33811 = ~n33825;
  assign n33819 = n33837 & n33838;
  assign n33826 = n33841 ^ n31542;
  assign n30778 = n33848 ^ n33849;
  assign n33842 = ~n33841;
  assign n33516 = ~n32396;
  assign n33757 = n33793 & n33794;
  assign n33795 = n33811 & n33812;
  assign n33776 = ~n33813;
  assign n33802 = n33819 ^ n33816;
  assign n30711 = n33826 ^ n33827;
  assign n33801 = ~n33819;
  assign n33803 = n33834 ^ n30778;
  assign n33839 = n33842 & n33843;
  assign n30727 = ~n30778;
  assign n33760 = ~n33757;
  assign n33774 = n33795 ^ n33796;
  assign n33762 = n33802 ^ n33803;
  assign n33797 = ~n33795;
  assign n33738 = n33805 ^ n30711;
  assign n33814 = n33803 & n33820;
  assign n30656 = ~n30711;
  assign n33815 = ~n33803;
  assign n33828 = ~n33839;
  assign n33758 = n130 ^ n33774;
  assign n33781 = n33762 & n129;
  assign n33783 = n33797 & n33798;
  assign n33780 = ~n33762;
  assign n33785 = n33738 & n33799;
  assign n33784 = ~n33738;
  assign n33779 = ~n33814;
  assign n33806 = n33815 & n33816;
  assign n33807 = n33828 & n33829;
  assign n33497 = n33757 ^ n33758;
  assign n33759 = ~n33758;
  assign n33777 = n33780 & n6214;
  assign n33744 = ~n33781;
  assign n33775 = ~n33783;
  assign n33782 = n33784 & n33754;
  assign n33766 = ~n33785;
  assign n33800 = ~n33806;
  assign n33786 = n33807 ^ n31473;
  assign n33808 = ~n33807;
  assign n33510 = ~n33497;
  assign n33726 = n33759 & n33760;
  assign n33761 = n33775 & n33776;
  assign n33764 = ~n33777;
  assign n33746 = ~n33782;
  assign n30568 = n33786 ^ n33787;
  assign n33788 = n33800 & n33801;
  assign n33804 = n33808 & n33809;
  assign n33729 = ~n33726;
  assign n33742 = n33761 ^ n33762;
  assign n33763 = ~n33761;
  assign n33708 = n33768 ^ n30568;
  assign n30604 = ~n30568;
  assign n33778 = ~n33788;
  assign n33789 = ~n33804;
  assign n33727 = n129 ^ n33742;
  assign n33748 = n33763 & n33764;
  assign n33750 = n33708 & n33765;
  assign n33749 = ~n33708;
  assign n33769 = n33778 & n33779;
  assign n33770 = n33789 & n33790;
  assign n32344 = n33726 ^ n33727;
  assign n33728 = ~n33727;
  assign n33743 = ~n33748;
  assign n33747 = n33749 & n33732;
  assign n33712 = ~n33750;
  assign n33753 = ~n33769;
  assign n33752 = n33770 ^ n33771;
  assign n33772 = ~n33770;
  assign n33438 = ~n32344;
  assign n33679 = n33728 & n33729;
  assign n33715 = n33743 & n33744;
  assign n33734 = ~n33747;
  assign n30549 = n33752 ^ n31418;
  assign n33737 = n33753 ^ n33754;
  assign n33751 = n33766 & n33753;
  assign n33767 = n33772 & n33773;
  assign n33682 = ~n33679;
  assign n33709 = ~n33715;
  assign n33673 = n33736 ^ n30549;
  assign n33716 = n33737 ^ n33738;
  assign n30490 = ~n30549;
  assign n33745 = ~n33751;
  assign n33755 = ~n33767;
  assign n33701 = n33715 ^ n33716;
  assign n33717 = n33716 & n6136;
  assign n33718 = n33673 & n33730;
  assign n33719 = ~n33673;
  assign n33720 = ~n33716;
  assign n33731 = n33745 & n33746;
  assign n33739 = n33755 & n33756;
  assign n33680 = n128 ^ n33701;
  assign n33710 = ~n33717;
  assign n33677 = ~n33718;
  assign n33713 = n33719 & n33697;
  assign n33714 = n33720 & n128;
  assign n33707 = n33731 ^ n33732;
  assign n33733 = ~n33731;
  assign n33723 = n33739 ^ n31427;
  assign n33740 = ~n33739;
  assign n33413 = n33679 ^ n33680;
  assign n33681 = ~n33680;
  assign n33675 = n33707 ^ n33708;
  assign n33702 = n33709 & n33710;
  assign n33699 = ~n33713;
  assign n33694 = ~n33714;
  assign n30458 = n33722 ^ n33723;
  assign n33721 = n33733 & n33734;
  assign n33735 = n33740 & n33741;
  assign n32283 = ~n33413;
  assign n33634 = n33681 & n33682;
  assign n33692 = n33675 & n143;
  assign n33691 = ~n33675;
  assign n33693 = ~n33702;
  assign n33641 = n33703 ^ n30458;
  assign n30421 = ~n30458;
  assign n33711 = ~n33721;
  assign n33724 = ~n33735;
  assign n33683 = n33691 & n6045;
  assign n33656 = ~n33692;
  assign n33674 = n33693 & n33694;
  assign n33684 = n33641 & n33695;
  assign n33685 = ~n33641;
  assign n33696 = n33711 & n33712;
  assign n33704 = n33724 & n33725;
  assign n33654 = n33674 ^ n33675;
  assign n33670 = ~n33683;
  assign n33671 = ~n33674;
  assign n33643 = ~n33684;
  assign n33678 = n33685 & n33661;
  assign n33672 = n33696 ^ n33697;
  assign n33698 = ~n33696;
  assign n33688 = n33704 ^ n31330;
  assign n33705 = ~n33704;
  assign n33635 = n143 ^ n33654;
  assign n33665 = n33670 & n33671;
  assign n33637 = n33672 ^ n33673;
  assign n33663 = ~n33678;
  assign n30388 = n33687 ^ n33688;
  assign n33686 = n33698 & n33699;
  assign n33700 = n33705 & n33706;
  assign n33360 = n33634 ^ n33635;
  assign n33596 = n33635 & n33634;
  assign n33658 = n33637 & n142;
  assign n33655 = ~n33665;
  assign n33657 = ~n33637;
  assign n33603 = n33666 ^ n30388;
  assign n30326 = ~n30388;
  assign n33676 = ~n33686;
  assign n33689 = ~n33700;
  assign n32249 = ~n33360;
  assign n33636 = n33655 & n33656;
  assign n33646 = n33657 & n5959;
  assign n33618 = ~n33658;
  assign n33647 = n33603 & n33659;
  assign n33648 = ~n33603;
  assign n33660 = n33676 & n33677;
  assign n33667 = n33689 & n33690;
  assign n33616 = n33636 ^ n33637;
  assign n33639 = ~n33636;
  assign n33638 = ~n33646;
  assign n33605 = ~n33647;
  assign n33645 = n33648 & n33623;
  assign n33640 = n33660 ^ n33661;
  assign n33662 = ~n33660;
  assign n33650 = n33667 ^ n31322;
  assign n33668 = ~n33667;
  assign n33597 = n142 ^ n33616;
  assign n33628 = n33638 & n33639;
  assign n33599 = n33640 ^ n33641;
  assign n33625 = ~n33645;
  assign n30233 = n33650 ^ n33651;
  assign n33649 = n33662 & n33663;
  assign n33664 = n33668 & n33669;
  assign n32214 = n33596 ^ n33597;
  assign n33558 = n33597 & n33596;
  assign n33620 = n33599 & n141;
  assign n33617 = ~n33628;
  assign n33619 = ~n33599;
  assign n33565 = n33629 ^ n30233;
  assign n33630 = n30233 & n33644;
  assign n30269 = ~n30233;
  assign n33642 = ~n33649;
  assign n33652 = ~n33664;
  assign n33335 = ~n32214;
  assign n33598 = n33617 & n33618;
  assign n33608 = n33619 & n5852;
  assign n33581 = ~n33620;
  assign n33609 = n33565 & n33621;
  assign n33610 = ~n33565;
  assign n33626 = n30269 & n32493;
  assign n32495 = ~n33630;
  assign n33622 = n33642 & n33643;
  assign n33631 = n33652 & n33653;
  assign n33579 = n33598 ^ n33599;
  assign n33600 = ~n33598;
  assign n33601 = ~n33608;
  assign n33567 = ~n33609;
  assign n33607 = n33610 & n33585;
  assign n33602 = n33622 ^ n33623;
  assign n32512 = ~n33626;
  assign n33624 = ~n33622;
  assign n33612 = n33631 ^ n31248;
  assign n33632 = ~n33631;
  assign n33559 = n141 ^ n33579;
  assign n33590 = n33600 & n33601;
  assign n33561 = n33602 ^ n33603;
  assign n33587 = ~n33607;
  assign n30160 = n33612 ^ n33613;
  assign n33611 = n33624 & n33625;
  assign n33627 = n33632 & n33633;
  assign n33279 = n33558 ^ n33559;
  assign n33521 = n33559 & n33558;
  assign n33583 = n33561 & n140;
  assign n33580 = ~n33590;
  assign n33582 = ~n33561;
  assign n33528 = n33591 ^ n30160;
  assign n33592 = n30160 & n33606;
  assign n30197 = ~n30160;
  assign n33604 = ~n33611;
  assign n33614 = ~n33627;
  assign n32175 = ~n33279;
  assign n33560 = n33580 & n33581;
  assign n33570 = n33582 & n5747;
  assign n33543 = ~n33583;
  assign n33573 = n33528 & n33547;
  assign n33571 = ~n33528;
  assign n32478 = ~n33592;
  assign n33588 = n30197 & n32460;
  assign n33584 = n33604 & n33605;
  assign n33593 = n33614 & n33615;
  assign n33541 = n33560 ^ n33561;
  assign n33562 = ~n33560;
  assign n33563 = ~n33570;
  assign n33569 = n33571 & n33572;
  assign n33549 = ~n33573;
  assign n33564 = n33584 ^ n33585;
  assign n32463 = ~n33588;
  assign n33586 = ~n33584;
  assign n33576 = n33593 ^ n31203;
  assign n33594 = ~n33593;
  assign n33522 = n140 ^ n33541;
  assign n33552 = n33562 & n33563;
  assign n33524 = n33564 ^ n33565;
  assign n33530 = ~n33569;
  assign n30134 = n33575 ^ n33576;
  assign n33574 = n33586 & n33587;
  assign n33589 = n33594 & n33595;
  assign n32136 = n33521 ^ n33522;
  assign n33476 = n33522 & n33521;
  assign n33545 = n33524 & n139;
  assign n33542 = ~n33552;
  assign n33544 = ~n33524;
  assign n33485 = n30134 ^ n33553;
  assign n33554 = n30134 & n33568;
  assign n30091 = ~n30134;
  assign n33566 = ~n33574;
  assign n33577 = ~n33589;
  assign n33255 = ~n32136;
  assign n33479 = ~n33476;
  assign n33523 = n33542 & n33543;
  assign n33532 = n33544 & n5694;
  assign n33502 = ~n33545;
  assign n33535 = n33485 & n33507;
  assign n33533 = ~n33485;
  assign n32430 = ~n33554;
  assign n33550 = n30091 & n32428;
  assign n33546 = n33566 & n33567;
  assign n33555 = n33577 & n33578;
  assign n33500 = n33523 ^ n33524;
  assign n33525 = ~n33523;
  assign n33526 = ~n33532;
  assign n33531 = n33533 & n33534;
  assign n33509 = ~n33535;
  assign n33527 = n33546 ^ n33547;
  assign n32447 = ~n33550;
  assign n33548 = ~n33546;
  assign n33538 = n33555 ^ n31193;
  assign n33556 = ~n33555;
  assign n33477 = n139 ^ n33500;
  assign n33513 = n33525 & n33526;
  assign n33481 = n33527 ^ n33528;
  assign n33487 = ~n33531;
  assign n30032 = n33537 ^ n33538;
  assign n33536 = n33548 & n33549;
  assign n33551 = n33556 & n33557;
  assign n32087 = n33476 ^ n33477;
  assign n33478 = ~n33477;
  assign n33503 = n33481 & n5626;
  assign n33501 = ~n33513;
  assign n33504 = ~n33481;
  assign n33449 = n33514 ^ n30032;
  assign n33515 = n30032 & n32396;
  assign n30040 = ~n30032;
  assign n33529 = ~n33536;
  assign n33539 = ~n33551;
  assign n33203 = ~n32087;
  assign n33442 = n33478 & n33479;
  assign n33480 = n33501 & n33502;
  assign n33483 = ~n33503;
  assign n33491 = n33504 & n138;
  assign n33492 = n33449 & n33505;
  assign n33493 = ~n33449;
  assign n32398 = ~n33515;
  assign n33511 = n30040 & n33516;
  assign n33506 = n33529 & n33530;
  assign n33517 = n33539 & n33540;
  assign n33457 = n33480 ^ n33481;
  assign n33482 = ~n33480;
  assign n33459 = ~n33491;
  assign n33451 = ~n33492;
  assign n33489 = n33493 & n33463;
  assign n33484 = n33506 ^ n33507;
  assign n32413 = ~n33511;
  assign n33508 = ~n33506;
  assign n29983 = n33517 ^ n33518;
  assign n33519 = ~n33517;
  assign n33443 = n138 ^ n33457;
  assign n33469 = n33482 & n33483;
  assign n33445 = n33484 ^ n33485;
  assign n33465 = ~n33489;
  assign n33430 = n29983 ^ n33495;
  assign n33494 = n33508 & n33509;
  assign n33496 = n29983 & n33510;
  assign n29934 = ~n29983;
  assign n33512 = n33519 & n33520;
  assign n33197 = n33442 ^ n33443;
  assign n33401 = n33443 & n33442;
  assign n33460 = n33445 & n5602;
  assign n33458 = ~n33469;
  assign n33461 = ~n33445;
  assign n33471 = n33430 & n33488;
  assign n33470 = ~n33430;
  assign n33486 = ~n33494;
  assign n32363 = ~n33496;
  assign n33490 = n29934 & n33497;
  assign n33498 = ~n33512;
  assign n33183 = ~n33197;
  assign n33404 = ~n33401;
  assign n33444 = n33458 & n33459;
  assign n33447 = ~n33460;
  assign n33452 = n33461 & n137;
  assign n33466 = n33470 & n33410;
  assign n33432 = ~n33471;
  assign n33462 = n33486 & n33487;
  assign n32382 = ~n33490;
  assign n33472 = n33498 & n33499;
  assign n33424 = n33444 ^ n33445;
  assign n33446 = ~n33444;
  assign n33426 = ~n33452;
  assign n33448 = n33462 ^ n33463;
  assign n33412 = ~n33466;
  assign n33464 = ~n33462;
  assign n33467 = n32382 & n32363;
  assign n33454 = n33472 ^ n33473;
  assign n33474 = ~n33472;
  assign n33402 = n137 ^ n33424;
  assign n33435 = n33446 & n33447;
  assign n33406 = n33448 ^ n33449;
  assign n29891 = n31011 ^ n33454;
  assign n33453 = n33464 & n33465;
  assign n32380 = ~n33467;
  assign n33468 = n33474 & n33475;
  assign n32009 = n33401 ^ n33402;
  assign n33403 = ~n33402;
  assign n33428 = n33406 & n136;
  assign n33425 = ~n33435;
  assign n33427 = ~n33406;
  assign n33390 = n33436 ^ n29891;
  assign n33437 = n29891 & n32344;
  assign n29926 = ~n29891;
  assign n33450 = ~n33453;
  assign n33455 = ~n33468;
  assign n33142 = ~n32009;
  assign n33365 = n33403 & n33404;
  assign n33405 = n33425 & n33426;
  assign n33415 = n33427 & n5544;
  assign n33385 = ~n33428;
  assign n33416 = n33390 & n33371;
  assign n33417 = ~n33390;
  assign n32324 = ~n33437;
  assign n33433 = n29926 & n33438;
  assign n33429 = n33450 & n33451;
  assign n33439 = n33455 & n33456;
  assign n33383 = n33405 ^ n33406;
  assign n33407 = ~n33405;
  assign n33408 = ~n33415;
  assign n33373 = ~n33416;
  assign n33414 = n33417 & n33418;
  assign n33409 = n33429 ^ n33430;
  assign n32346 = ~n33433;
  assign n33431 = ~n33429;
  assign n33420 = n33439 ^ n31048;
  assign n33440 = ~n33439;
  assign n33366 = n136 ^ n33383;
  assign n33395 = n33407 & n33408;
  assign n33346 = n33409 ^ n33410;
  assign n33392 = ~n33414;
  assign n29876 = n33420 ^ n33421;
  assign n33419 = n33431 & n33432;
  assign n33434 = n33440 & n33441;
  assign n31911 = n33365 ^ n33366;
  assign n33323 = n33366 & n33365;
  assign n33387 = n33346 & n151;
  assign n33384 = ~n33395;
  assign n33386 = ~n33346;
  assign n33353 = n33396 ^ n29876;
  assign n33397 = n29876 & n33413;
  assign n29841 = ~n29876;
  assign n33411 = ~n33419;
  assign n33422 = ~n33434;
  assign n33101 = ~n31911;
  assign n33326 = ~n33323;
  assign n33367 = n33384 & n33385;
  assign n33375 = n33386 & n5509;
  assign n33348 = ~n33387;
  assign n33377 = n33353 & n33388;
  assign n33376 = ~n33353;
  assign n33393 = n29841 & n32283;
  assign n32307 = ~n33397;
  assign n33389 = n33411 & n33412;
  assign n33398 = n33422 & n33423;
  assign n33345 = n151 ^ n33367;
  assign n33368 = ~n33367;
  assign n33369 = ~n33375;
  assign n33374 = n33376 & n33332;
  assign n33355 = ~n33377;
  assign n33370 = n33389 ^ n33390;
  assign n32286 = ~n33393;
  assign n33391 = ~n33389;
  assign n33380 = n33398 ^ n30979;
  assign n33399 = ~n33398;
  assign n33324 = n33345 ^ n33346;
  assign n33358 = n33368 & n33369;
  assign n33328 = n33370 ^ n33371;
  assign n33334 = ~n33374;
  assign n29823 = n33379 ^ n33380;
  assign n33378 = n33391 & n33392;
  assign n33394 = n33399 & n33400;
  assign n31841 = n33323 ^ n33324;
  assign n33325 = ~n33324;
  assign n33349 = n33328 & n5464;
  assign n33347 = ~n33358;
  assign n33350 = ~n33328;
  assign n33293 = n33359 ^ n29823;
  assign n33361 = n29823 & n32249;
  assign n29862 = ~n29823;
  assign n33372 = ~n33378;
  assign n33381 = ~n33394;
  assign n33050 = ~n31841;
  assign n33284 = n33325 & n33326;
  assign n33327 = n33347 & n33348;
  assign n33330 = ~n33349;
  assign n33337 = n33350 & n150;
  assign n33338 = n33293 & n33351;
  assign n33339 = ~n33293;
  assign n33356 = n29862 & n33360;
  assign n32251 = ~n33361;
  assign n33352 = n33372 & n33373;
  assign n33362 = n33381 & n33382;
  assign n33287 = ~n33284;
  assign n33306 = n33327 ^ n33328;
  assign n33329 = ~n33327;
  assign n33308 = ~n33337;
  assign n33295 = ~n33338;
  assign n33336 = n33339 & n33312;
  assign n33331 = n33352 ^ n33353;
  assign n32270 = ~n33356;
  assign n33354 = ~n33352;
  assign n33342 = n33362 ^ n30839;
  assign n33363 = ~n33362;
  assign n33285 = n150 ^ n33306;
  assign n33317 = n33329 & n33330;
  assign n33289 = n33331 ^ n33332;
  assign n33314 = ~n33336;
  assign n29835 = n33341 ^ n33342;
  assign n33340 = n33354 & n33355;
  assign n33357 = n33363 & n33364;
  assign n32986 = n33284 ^ n33285;
  assign n33286 = ~n33285;
  assign n33310 = n33289 & n149;
  assign n33307 = ~n33317;
  assign n33309 = ~n33289;
  assign n33251 = n33318 ^ n29835;
  assign n33319 = n29835 & n33335;
  assign n29789 = ~n29835;
  assign n33333 = ~n33340;
  assign n33343 = ~n33357;
  assign n31774 = ~n32986;
  assign n33245 = n33286 & n33287;
  assign n33288 = n33307 & n33308;
  assign n33297 = n33309 & n5423;
  assign n33267 = ~n33310;
  assign n33298 = n33251 & n33272;
  assign n33299 = ~n33251;
  assign n32216 = ~n33319;
  assign n33315 = n29789 & n32214;
  assign n33311 = n33333 & n33334;
  assign n33320 = n33343 & n33344;
  assign n33265 = n33288 ^ n33289;
  assign n33290 = ~n33288;
  assign n33291 = ~n33297;
  assign n33254 = ~n33298;
  assign n33296 = n33299 & n33300;
  assign n33292 = n33311 ^ n33312;
  assign n32235 = ~n33315;
  assign n33313 = ~n33311;
  assign n33302 = n33320 ^ n30768;
  assign n33321 = ~n33320;
  assign n33246 = n149 ^ n33265;
  assign n33277 = n33290 & n33291;
  assign n33248 = n33292 ^ n33293;
  assign n33274 = ~n33296;
  assign n29798 = n33302 ^ n33303;
  assign n33301 = n33313 & n33314;
  assign n33316 = n33321 & n33322;
  assign n31709 = n33245 ^ n33246;
  assign n33208 = n33246 & n33245;
  assign n33269 = n33248 & n148;
  assign n33266 = ~n33277;
  assign n33268 = ~n33248;
  assign n33215 = n33278 ^ n29798;
  assign n33280 = n29798 & n32175;
  assign n29750 = ~n29798;
  assign n33294 = ~n33301;
  assign n33304 = ~n33316;
  assign n32948 = ~n31709;
  assign n33247 = n33266 & n33267;
  assign n33257 = n33268 & n5391;
  assign n33230 = ~n33269;
  assign n33259 = n33215 & n33270;
  assign n33258 = ~n33215;
  assign n33275 = n29750 & n33279;
  assign n32178 = ~n33280;
  assign n33271 = n33294 & n33295;
  assign n33281 = n33304 & n33305;
  assign n33228 = n33247 ^ n33248;
  assign n33249 = ~n33247;
  assign n33250 = ~n33257;
  assign n33256 = n33258 & n33234;
  assign n33217 = ~n33259;
  assign n33252 = n33271 ^ n33272;
  assign n32199 = ~n33275;
  assign n33273 = ~n33271;
  assign n33261 = n33281 ^ n30671;
  assign n33282 = ~n33281;
  assign n33209 = n148 ^ n33228;
  assign n33240 = n33249 & n33250;
  assign n33211 = n33251 ^ n33252;
  assign n33236 = ~n33256;
  assign n29713 = n33261 ^ n33262;
  assign n33260 = n33273 & n33274;
  assign n33276 = n33282 & n33283;
  assign n31632 = n33208 ^ n33209;
  assign n32827 = n33209 & n33208;
  assign n33231 = n33211 & n5352;
  assign n33229 = ~n33240;
  assign n33232 = ~n33211;
  assign n33241 = n29713 & n33255;
  assign n29760 = ~n29713;
  assign n33253 = ~n33260;
  assign n33263 = ~n33276;
  assign n32889 = ~n31632;
  assign n33210 = n33229 & n33230;
  assign n33213 = ~n33231;
  assign n33222 = n33232 & n147;
  assign n33173 = n33237 ^ n29760;
  assign n32139 = ~n33241;
  assign n33238 = n29760 & n32136;
  assign n33233 = n33253 & n33254;
  assign n33242 = n33263 & n33264;
  assign n33187 = n33210 ^ n33211;
  assign n33212 = ~n33210;
  assign n33189 = ~n33222;
  assign n33219 = n33173 & n33194;
  assign n33214 = n33233 ^ n33234;
  assign n33220 = ~n33173;
  assign n32160 = ~n33238;
  assign n33235 = ~n33233;
  assign n33225 = n33242 ^ n30660;
  assign n33243 = ~n33242;
  assign n32861 = n147 ^ n33187;
  assign n33200 = n33212 & n33213;
  assign n33169 = n33214 ^ n33215;
  assign n33196 = ~n33219;
  assign n33218 = n33220 & n33221;
  assign n29673 = n33224 ^ n33225;
  assign n33223 = n33235 & n33236;
  assign n33239 = n33243 & n33244;
  assign n33167 = ~n32861;
  assign n33191 = n33169 & n146;
  assign n33188 = ~n33200;
  assign n33190 = ~n33169;
  assign n33139 = n33201 ^ n29673;
  assign n33175 = ~n33218;
  assign n33202 = n29673 & n32087;
  assign n29722 = ~n29673;
  assign n33216 = ~n33223;
  assign n33226 = ~n33239;
  assign n33130 = n33167 & n32827;
  assign n33168 = n33188 & n33189;
  assign n33179 = n33190 & n5311;
  assign n33151 = ~n33191;
  assign n33181 = n33139 & n33192;
  assign n33180 = ~n33139;
  assign n32090 = ~n33202;
  assign n33198 = n29722 & n33203;
  assign n33193 = n33216 & n33217;
  assign n33204 = n33226 & n33227;
  assign n33133 = ~n33130;
  assign n33149 = n33168 ^ n33169;
  assign n33170 = ~n33168;
  assign n33171 = ~n33179;
  assign n33176 = n33180 & n33155;
  assign n33141 = ~n33181;
  assign n33172 = n33193 ^ n33194;
  assign n32115 = ~n33198;
  assign n33195 = ~n33193;
  assign n29620 = n33204 ^ n33205;
  assign n33206 = ~n33204;
  assign n33131 = n146 ^ n33149;
  assign n33162 = n33170 & n33171;
  assign n33135 = n33172 ^ n33173;
  assign n33157 = ~n33176;
  assign n33182 = n33195 & n33196;
  assign n33184 = n29620 & n33197;
  assign n29692 = ~n29620;
  assign n33199 = n33206 & n33207;
  assign n31274 = n33130 ^ n33131;
  assign n33132 = ~n33131;
  assign n33152 = n33135 & n5261;
  assign n33150 = ~n33162;
  assign n33153 = ~n33135;
  assign n33118 = n33177 ^ n29692;
  assign n33174 = ~n33182;
  assign n33178 = n29692 & n33183;
  assign n32037 = ~n33184;
  assign n33185 = ~n33199;
  assign n33086 = n31274 ^ n33110;
  assign n33016 = n31274 & n31268;
  assign n33089 = n33132 & n33133;
  assign n33134 = n33150 & n33151;
  assign n33137 = ~n33152;
  assign n33143 = n33153 & n145;
  assign n33160 = n33118 & n33163;
  assign n33154 = n33174 & n33175;
  assign n33159 = ~n33118;
  assign n32066 = ~n33178;
  assign n33164 = n33185 & n33186;
  assign n29400 = n33085 ^ n33086;
  assign n32366 = n231 ^ n33086;
  assign n32835 = n33086 & n231;
  assign n33087 = ~n33086;
  assign n33092 = ~n33089;
  assign n33111 = n33134 ^ n33135;
  assign n33136 = ~n33134;
  assign n33113 = ~n33143;
  assign n33138 = n33154 ^ n33155;
  assign n33158 = n33159 & n33098;
  assign n33120 = ~n33160;
  assign n33156 = ~n33154;
  assign n32063 = n32037 & n32066;
  assign n33146 = n33164 ^ n30411;
  assign n33165 = ~n33164;
  assign n33075 = n32835 & n230;
  assign n32360 = ~n32366;
  assign n32867 = n33087 & n33088;
  assign n33074 = ~n32835;
  assign n33090 = n145 ^ n33111;
  assign n33123 = n33136 & n33137;
  assign n33094 = n33138 ^ n33139;
  assign n29685 = n33145 ^ n33146;
  assign n33144 = n33156 & n33157;
  assign n33100 = ~n33158;
  assign n33161 = n33165 & n33166;
  assign n33061 = n33074 & n19809;
  assign n32807 = ~n33075;
  assign n33076 = n33089 ^ n33090;
  assign n33091 = ~n33090;
  assign n33115 = n33094 & n144;
  assign n33112 = ~n33123;
  assign n33114 = ~n33094;
  assign n33071 = n33124 ^ n29685;
  assign n33125 = n29685 & n33142;
  assign n29587 = ~n29685;
  assign n33140 = ~n33144;
  assign n33147 = ~n33161;
  assign n32839 = ~n33061;
  assign n33062 = n33076 & n31242;
  assign n33063 = ~n33076;
  assign n33041 = n33091 & n33092;
  assign n33093 = n33112 & n33113;
  assign n33103 = n33114 & n5208;
  assign n33066 = ~n33115;
  assign n33104 = n33071 & n33116;
  assign n33105 = ~n33071;
  assign n31980 = ~n33125;
  assign n33121 = n29587 & n32009;
  assign n33117 = n33140 & n33141;
  assign n33126 = n33147 & n33148;
  assign n33040 = ~n33062;
  assign n33052 = n33063 & n31086;
  assign n33064 = n33093 ^ n33094;
  assign n33095 = ~n33093;
  assign n33096 = ~n33103;
  assign n33073 = ~n33104;
  assign n33102 = n33105 & n33047;
  assign n33097 = n33117 ^ n33118;
  assign n32011 = ~n33121;
  assign n33119 = ~n33117;
  assign n33107 = n33126 ^ n33127;
  assign n33128 = ~n33126;
  assign n33039 = n33040 & n33016;
  assign n33029 = ~n33052;
  assign n33042 = n144 ^ n33064;
  assign n33079 = n33095 & n33096;
  assign n33019 = n33097 ^ n33098;
  assign n33049 = ~n33102;
  assign n29645 = n33107 ^ n30338;
  assign n33106 = n33119 & n33120;
  assign n33122 = n33128 & n33129;
  assign n33028 = ~n33039;
  assign n33015 = n33040 & n33029;
  assign n33030 = n33041 ^ n33042;
  assign n32991 = n33042 & n33041;
  assign n33068 = n33019 & n159;
  assign n33065 = ~n33079;
  assign n33067 = ~n33019;
  assign n33025 = n33080 ^ n29645;
  assign n33081 = n29645 & n33101;
  assign n29549 = ~n29645;
  assign n33099 = ~n33106;
  assign n33108 = ~n33122;
  assign n29335 = n33015 ^ n33016;
  assign n33001 = n33028 & n33029;
  assign n33017 = n33030 & n31080;
  assign n32978 = ~n33030;
  assign n33043 = n33065 & n33066;
  assign n33053 = n33067 & n5179;
  assign n33021 = ~n33068;
  assign n33054 = n33025 & n33069;
  assign n33055 = ~n33025;
  assign n31914 = ~n33081;
  assign n33077 = n29549 & n31911;
  assign n33070 = n33099 & n33100;
  assign n33082 = n33108 & n33109;
  assign n32041 = n31086 ^ n29335;
  assign n32977 = n33001 ^ n31080;
  assign n29384 = ~n29335;
  assign n33003 = ~n33001;
  assign n33002 = ~n33017;
  assign n33005 = n32978 & n31060;
  assign n33018 = n159 ^ n33043;
  assign n33044 = ~n33043;
  assign n33045 = ~n33053;
  assign n33027 = ~n33054;
  assign n33051 = n33055 & n32998;
  assign n33046 = n33070 ^ n33071;
  assign n31947 = ~n33077;
  assign n33072 = ~n33070;
  assign n33057 = n33082 ^ n30302;
  assign n33083 = ~n33082;
  assign n32950 = n32041 ^ n31985;
  assign n29324 = n32977 ^ n32978;
  assign n32990 = n33002 & n33003;
  assign n32980 = ~n33005;
  assign n32992 = n33018 ^ n33019;
  assign n33033 = n33044 & n33045;
  assign n32994 = n33046 ^ n33047;
  assign n33000 = ~n33051;
  assign n29530 = n33057 ^ n33058;
  assign n33056 = n33072 & n33073;
  assign n33078 = n33083 & n33084;
  assign n32936 = n32950 & n32951;
  assign n32002 = n29324 ^ n31060;
  assign n32934 = ~n32950;
  assign n29332 = ~n29324;
  assign n32979 = ~n32990;
  assign n32924 = n32991 ^ n32992;
  assign n32938 = n32992 & n32991;
  assign n33023 = n32994 & n158;
  assign n33020 = ~n33033;
  assign n33022 = ~n32994;
  assign n32945 = n33034 ^ n29530;
  assign n33035 = n29530 & n33050;
  assign n29554 = ~n29530;
  assign n33048 = ~n33056;
  assign n33059 = ~n33078;
  assign n32805 = n32002 ^ n31956;
  assign n32928 = n32934 & n32935;
  assign n32875 = ~n32936;
  assign n32952 = n32979 & n32980;
  assign n32966 = n32924 & n30981;
  assign n32965 = ~n32924;
  assign n32993 = n33020 & n33021;
  assign n33006 = n33022 & n5130;
  assign n32969 = ~n33023;
  assign n33009 = n32945 & n32974;
  assign n33007 = ~n32945;
  assign n33031 = n29554 & n31841;
  assign n31878 = ~n33035;
  assign n33024 = n33048 & n33049;
  assign n33036 = n33059 & n33060;
  assign n32894 = n32805 & n32841;
  assign n32892 = ~n32805;
  assign n32909 = ~n32928;
  assign n32923 = n32952 ^ n30981;
  assign n32953 = ~n32952;
  assign n32956 = n32965 & n31017;
  assign n32954 = ~n32966;
  assign n32967 = n32993 ^ n32994;
  assign n32995 = ~n32993;
  assign n32996 = ~n33006;
  assign n33004 = n33007 & n33008;
  assign n32976 = ~n33009;
  assign n32997 = n33024 ^ n33025;
  assign n31844 = ~n33031;
  assign n33026 = ~n33024;
  assign n33012 = n33036 ^ n30217;
  assign n33037 = ~n33036;
  assign n32873 = n32892 & n32893;
  assign n32812 = ~n32894;
  assign n32899 = n32909 & n32867;
  assign n32900 = n32909 & n32875;
  assign n29290 = n32923 ^ n32924;
  assign n32937 = n32953 & n32954;
  assign n32926 = ~n32956;
  assign n32939 = n158 ^ n32967;
  assign n32983 = n32995 & n32996;
  assign n32941 = n32997 ^ n32998;
  assign n32947 = ~n33004;
  assign n29518 = n33011 ^ n33012;
  assign n33010 = n33026 & n33027;
  assign n33032 = n33037 & n33038;
  assign n32847 = ~n32873;
  assign n32874 = ~n32899;
  assign n32868 = ~n32900;
  assign n29300 = ~n29290;
  assign n32925 = ~n32937;
  assign n32862 = n32938 ^ n32939;
  assign n32877 = n32939 & n32938;
  assign n32971 = n32941 & n157;
  assign n32968 = ~n32983;
  assign n32970 = ~n32941;
  assign n32886 = n32984 ^ n29518;
  assign n32985 = n29518 & n31774;
  assign n29493 = ~n29518;
  assign n32999 = ~n33010;
  assign n33013 = ~n33032;
  assign n32836 = n32867 ^ n32868;
  assign n32869 = n32874 & n32875;
  assign n31922 = n31017 ^ n29300;
  assign n32895 = n32925 & n32926;
  assign n32911 = n32862 & n30889;
  assign n32910 = ~n32862;
  assign n32880 = ~n32877;
  assign n32940 = n32968 & n32969;
  assign n32957 = n32970 & n5088;
  assign n32914 = ~n32971;
  assign n32959 = n32886 & n32972;
  assign n32958 = ~n32886;
  assign n31776 = ~n32985;
  assign n32981 = n29493 & n32986;
  assign n32973 = n32999 & n33000;
  assign n32987 = n33013 & n33014;
  assign n32803 = n32835 ^ n32836;
  assign n32753 = n31922 ^ n31910;
  assign n32838 = ~n32836;
  assign n32840 = ~n32869;
  assign n32863 = n32895 ^ n30914;
  assign n32897 = ~n32895;
  assign n32901 = n32910 & n30914;
  assign n32896 = ~n32911;
  assign n32912 = n32940 ^ n32941;
  assign n32942 = ~n32940;
  assign n32943 = ~n32957;
  assign n32955 = n32958 & n32918;
  assign n32888 = ~n32959;
  assign n32944 = n32973 ^ n32974;
  assign n31813 = ~n32981;
  assign n32975 = ~n32973;
  assign n32961 = n32987 ^ n30146;
  assign n32988 = ~n32987;
  assign n31171 = n230 ^ n32803;
  assign n32813 = n32753 & n32831;
  assign n32832 = n32838 & n32839;
  assign n32814 = ~n32753;
  assign n32804 = n32840 ^ n32841;
  assign n32837 = n32847 & n32840;
  assign n29272 = n32862 ^ n32863;
  assign n32876 = n32896 & n32897;
  assign n32865 = ~n32901;
  assign n32878 = n157 ^ n32912;
  assign n32929 = n32942 & n32943;
  assign n32882 = n32944 ^ n32945;
  assign n32920 = ~n32955;
  assign n29458 = n32961 ^ n32962;
  assign n32960 = n32975 & n32976;
  assign n32982 = n32988 & n32989;
  assign n32304 = ~n31171;
  assign n32777 = n32804 ^ n32805;
  assign n32755 = ~n32813;
  assign n32808 = n32814 & n32785;
  assign n32806 = ~n32832;
  assign n31855 = n29272 ^ n30914;
  assign n32811 = ~n32837;
  assign n29256 = ~n29272;
  assign n32864 = ~n32876;
  assign n32802 = n32877 ^ n32878;
  assign n32879 = ~n32878;
  assign n32915 = n32882 & n5043;
  assign n32913 = ~n32929;
  assign n32916 = ~n32882;
  assign n32826 = n32930 ^ n29458;
  assign n32931 = n29458 & n32948;
  assign n29482 = ~n29458;
  assign n32946 = ~n32960;
  assign n32963 = ~n32982;
  assign n32779 = n32777 & n229;
  assign n32703 = n31855 ^ n31786;
  assign n32778 = ~n32777;
  assign n32776 = n32806 & n32807;
  assign n32786 = ~n32808;
  assign n32784 = n32811 & n32812;
  assign n32833 = n32864 & n32865;
  assign n32848 = n32802 & n30860;
  assign n32849 = ~n32802;
  assign n32817 = n32879 & n32880;
  assign n32881 = n32913 & n32914;
  assign n32884 = ~n32915;
  assign n32902 = n32916 & n156;
  assign n32903 = n32826 & n32857;
  assign n32904 = ~n32826;
  assign n32927 = n29482 & n31709;
  assign n31711 = ~n32931;
  assign n32917 = n32946 & n32947;
  assign n32932 = n32963 & n32964;
  assign n32747 = n32776 ^ n32777;
  assign n32772 = n32778 & n19742;
  assign n32773 = n32703 & n32731;
  assign n32724 = ~n32779;
  assign n32752 = n32784 ^ n32785;
  assign n32774 = ~n32703;
  assign n32749 = ~n32776;
  assign n32787 = ~n32784;
  assign n32801 = n32833 ^ n30797;
  assign n32815 = ~n32833;
  assign n32789 = ~n32848;
  assign n32842 = n32849 & n30797;
  assign n32820 = ~n32817;
  assign n32850 = n32881 ^ n32882;
  assign n32883 = ~n32881;
  assign n32852 = ~n32902;
  assign n32830 = ~n32903;
  assign n32898 = n32904 & n32905;
  assign n32885 = n32917 ^ n32918;
  assign n31744 = ~n32927;
  assign n32919 = ~n32917;
  assign n32908 = n32932 ^ n30129;
  assign n32933 = n32932 & n32949;
  assign n31127 = n229 ^ n32747;
  assign n32698 = n32752 ^ n32753;
  assign n32748 = ~n32772;
  assign n32705 = ~n32773;
  assign n32756 = n32774 & n32775;
  assign n32780 = n32786 & n32787;
  assign n29224 = n32801 ^ n32802;
  assign n32816 = ~n32842;
  assign n32818 = n156 ^ n32850;
  assign n32870 = n32883 & n32884;
  assign n32822 = n32885 ^ n32886;
  assign n32859 = ~n32898;
  assign n29496 = n32907 ^ n32908;
  assign n32906 = n32919 & n32920;
  assign n32921 = ~n32933;
  assign n32729 = n32698 & n228;
  assign n32273 = ~n31127;
  assign n32728 = ~n32698;
  assign n32746 = n32748 & n32749;
  assign n32732 = ~n32756;
  assign n31788 = n30860 ^ n29224;
  assign n32754 = ~n32780;
  assign n29215 = ~n29224;
  assign n32809 = n32815 & n32816;
  assign n32734 = n32817 ^ n32818;
  assign n32819 = ~n32818;
  assign n32854 = n32822 & n155;
  assign n32851 = ~n32870;
  assign n32853 = ~n32822;
  assign n32769 = n32871 ^ n29496;
  assign n32872 = n29496 & n32889;
  assign n29430 = ~n29496;
  assign n32887 = ~n32906;
  assign n32890 = n32921 & n32922;
  assign n32722 = n32728 & n19716;
  assign n32677 = ~n32729;
  assign n32723 = ~n32746;
  assign n32663 = n31788 ^ n31705;
  assign n32730 = n32754 & n32755;
  assign n32790 = n32734 & n30727;
  assign n32788 = ~n32809;
  assign n32791 = ~n32734;
  assign n32760 = n32819 & n32820;
  assign n32821 = n32851 & n32852;
  assign n32843 = n32853 & n5010;
  assign n32794 = ~n32854;
  assign n32844 = n32769 & n32855;
  assign n32845 = ~n32769;
  assign n31635 = ~n32872;
  assign n32866 = n29430 & n31632;
  assign n32856 = n32887 & n32888;
  assign n29446 = n32890 ^ n32891;
  assign n32699 = ~n32722;
  assign n32718 = n32723 & n32724;
  assign n32719 = n32663 & n32684;
  assign n32702 = n32730 ^ n32731;
  assign n32720 = ~n32663;
  assign n32733 = ~n32730;
  assign n32757 = n32788 & n32789;
  assign n32758 = ~n32790;
  assign n32781 = n32791 & n30778;
  assign n32763 = ~n32760;
  assign n32792 = n32821 ^ n32822;
  assign n32823 = ~n32821;
  assign n32824 = ~n32843;
  assign n32771 = ~n32844;
  assign n32834 = n32845 & n32798;
  assign n32825 = n32856 ^ n32857;
  assign n32717 = n32860 ^ n29446;
  assign n32828 = n32861 ^ n29446;
  assign n31672 = ~n32866;
  assign n32858 = ~n32856;
  assign n32657 = n32702 ^ n32703;
  assign n32697 = ~n32718;
  assign n32665 = ~n32719;
  assign n32706 = n32720 & n32721;
  assign n32725 = n32732 & n32733;
  assign n32735 = n32757 ^ n30778;
  assign n32759 = ~n32757;
  assign n32737 = ~n32781;
  assign n32761 = n155 ^ n32792;
  assign n32810 = n32823 & n32824;
  assign n32765 = n32825 ^ n32826;
  assign n31602 = n32827 ^ n32828;
  assign n32800 = ~n32834;
  assign n32846 = n32858 & n32859;
  assign n32681 = n32657 & n19695;
  assign n32674 = n32697 ^ n32698;
  assign n32696 = n32699 & n32697;
  assign n32682 = ~n32657;
  assign n32685 = ~n32706;
  assign n32704 = ~n32725;
  assign n29165 = n32734 ^ n32735;
  assign n32750 = n32758 & n32759;
  assign n32687 = n32760 ^ n32761;
  assign n32762 = ~n32761;
  assign n32795 = n32765 & n4987;
  assign n32793 = ~n32810;
  assign n32796 = ~n32765;
  assign n32829 = ~n32846;
  assign n31037 = n228 ^ n32674;
  assign n32658 = ~n32681;
  assign n32678 = n32682 & n227;
  assign n32676 = ~n32696;
  assign n32683 = n32704 & n32705;
  assign n31715 = n29165 ^ n30778;
  assign n29193 = ~n29165;
  assign n32739 = n32687 & n30711;
  assign n32736 = ~n32750;
  assign n32738 = ~n32687;
  assign n32710 = n32762 & n32763;
  assign n32764 = n32793 & n32794;
  assign n32767 = ~n32795;
  assign n32782 = n32796 & n154;
  assign n32797 = n32829 & n32830;
  assign n32232 = ~n31037;
  assign n32656 = n32676 & n32677;
  assign n32637 = ~n32678;
  assign n32662 = n32683 ^ n32684;
  assign n32624 = n31715 ^ n31706;
  assign n32686 = ~n32683;
  assign n32707 = n32736 & n32737;
  assign n32726 = n32738 & n30656;
  assign n32690 = ~n32739;
  assign n32740 = n32764 ^ n32765;
  assign n32766 = ~n32764;
  assign n32742 = ~n32782;
  assign n32768 = n32797 ^ n32798;
  assign n32799 = ~n32797;
  assign n32635 = n32656 ^ n32657;
  assign n32618 = n32662 ^ n32663;
  assign n32659 = ~n32656;
  assign n32668 = n32624 & n32644;
  assign n32666 = ~n32624;
  assign n32679 = n32685 & n32686;
  assign n32688 = n32707 ^ n30711;
  assign n32708 = ~n32707;
  assign n32709 = ~n32726;
  assign n32711 = n154 ^ n32740;
  assign n32751 = n32766 & n32767;
  assign n32713 = n32768 ^ n32769;
  assign n32783 = n32799 & n32800;
  assign n30964 = n227 ^ n32635;
  assign n32641 = n32618 & n19641;
  assign n32653 = n32658 & n32659;
  assign n32642 = ~n32618;
  assign n32660 = n32666 & n32667;
  assign n32626 = ~n32668;
  assign n32664 = ~n32679;
  assign n29141 = n32687 ^ n32688;
  assign n32700 = n32708 & n32709;
  assign n32648 = n32710 ^ n32711;
  assign n32672 = n32711 & n32710;
  assign n32744 = n32713 & n153;
  assign n32741 = ~n32751;
  assign n32743 = ~n32713;
  assign n32770 = ~n32783;
  assign n32202 = ~n30964;
  assign n32619 = ~n32641;
  assign n32638 = n32642 & n226;
  assign n32636 = ~n32653;
  assign n32646 = ~n32660;
  assign n32643 = n32664 & n32665;
  assign n31643 = n29141 ^ n30711;
  assign n29169 = ~n29141;
  assign n32691 = n32648 & n30568;
  assign n32689 = ~n32700;
  assign n32692 = ~n32648;
  assign n32675 = ~n32672;
  assign n32712 = n32741 & n32742;
  assign n32727 = n32743 & n4946;
  assign n32695 = ~n32744;
  assign n32745 = n32770 & n32771;
  assign n32617 = n32636 & n32637;
  assign n32599 = ~n32638;
  assign n32623 = n32643 ^ n32644;
  assign n32590 = n31643 ^ n31542;
  assign n32645 = ~n32643;
  assign n32669 = n32689 & n32690;
  assign n32650 = ~n32691;
  assign n32680 = n32692 & n30604;
  assign n32693 = n32712 ^ n32713;
  assign n32714 = ~n32712;
  assign n32715 = ~n32727;
  assign n32716 = n152 ^ n32745;
  assign n32597 = n32617 ^ n32618;
  assign n32583 = n32623 ^ n32624;
  assign n32620 = ~n32617;
  assign n32627 = n32590 & n32632;
  assign n32628 = ~n32590;
  assign n32639 = n32645 & n32646;
  assign n32647 = n32669 ^ n30604;
  assign n32670 = ~n32669;
  assign n32671 = ~n32680;
  assign n32673 = n153 ^ n32693;
  assign n32701 = n32714 & n32715;
  assign n32634 = n32716 ^ n32717;
  assign n30855 = n226 ^ n32597;
  assign n32603 = n32583 & n19596;
  assign n32614 = n32619 & n32620;
  assign n32604 = ~n32583;
  assign n32592 = ~n32627;
  assign n32621 = n32628 & n32606;
  assign n32625 = ~n32639;
  assign n29139 = n32647 ^ n32648;
  assign n32661 = n32670 & n32671;
  assign n32610 = n32672 ^ n32673;
  assign n32655 = n32673 & n32675;
  assign n32694 = ~n32701;
  assign n30911 = ~n30855;
  assign n32584 = ~n32603;
  assign n32600 = n32604 & n225;
  assign n32598 = ~n32614;
  assign n32608 = ~n32621;
  assign n32605 = n32625 & n32626;
  assign n31579 = n29139 ^ n30604;
  assign n29110 = ~n29139;
  assign n32652 = n32610 & n30549;
  assign n32649 = ~n32661;
  assign n32651 = ~n32610;
  assign n32654 = n32694 & n32695;
  assign n32582 = n32598 & n32599;
  assign n32568 = ~n32600;
  assign n32589 = n32605 ^ n32606;
  assign n32557 = n31579 ^ n31552;
  assign n32607 = ~n32605;
  assign n32629 = n32649 & n32650;
  assign n32640 = n32651 & n30490;
  assign n32613 = ~n32652;
  assign n32633 = n32654 ^ n32655;
  assign n32566 = n32582 ^ n32583;
  assign n32551 = n32589 ^ n32590;
  assign n32585 = ~n32582;
  assign n32595 = n32557 & n32576;
  assign n32593 = ~n32557;
  assign n32601 = n32607 & n32608;
  assign n32609 = n32629 ^ n30490;
  assign n32571 = n32633 ^ n32634;
  assign n32630 = ~n32629;
  assign n32631 = ~n32640;
  assign n32548 = n225 ^ n32566;
  assign n32574 = n32551 & n224;
  assign n32581 = n32584 & n32585;
  assign n32573 = ~n32551;
  assign n32586 = n32593 & n32594;
  assign n32578 = ~n32595;
  assign n32591 = ~n32601;
  assign n29108 = n32609 ^ n32610;
  assign n32616 = n32571 & n30421;
  assign n32615 = ~n32571;
  assign n32622 = n32630 & n32631;
  assign n30805 = n32548 ^ n30855;
  assign n32549 = ~n32548;
  assign n32569 = n32573 & n19565;
  assign n32534 = ~n32574;
  assign n32567 = ~n32581;
  assign n32559 = ~n32586;
  assign n32575 = n32591 & n32592;
  assign n31514 = n29108 ^ n30549;
  assign n29076 = ~n29108;
  assign n32611 = n32615 & n30458;
  assign n32596 = ~n32616;
  assign n32612 = ~n32622;
  assign n32119 = ~n30805;
  assign n32513 = n32549 & n30911;
  assign n32550 = n32567 & n32568;
  assign n32553 = ~n32569;
  assign n32556 = n32575 ^ n32576;
  assign n32527 = n31514 ^ n31418;
  assign n32577 = ~n32575;
  assign n32580 = ~n32611;
  assign n32602 = n32612 & n32613;
  assign n32516 = ~n32513;
  assign n32532 = n32550 ^ n32551;
  assign n32518 = n32556 ^ n32557;
  assign n32552 = ~n32550;
  assign n32561 = n32527 & n32564;
  assign n32560 = ~n32527;
  assign n32570 = n32577 & n32578;
  assign n32588 = ~n32602;
  assign n32514 = n224 ^ n32532;
  assign n32538 = n32518 & n19533;
  assign n32546 = n32552 & n32553;
  assign n32539 = ~n32518;
  assign n32554 = n32560 & n32541;
  assign n32529 = ~n32561;
  assign n32558 = ~n32570;
  assign n32572 = n32588 ^ n30458;
  assign n32587 = n32588 & n32596;
  assign n30735 = n32513 ^ n32514;
  assign n32515 = ~n32514;
  assign n32520 = ~n32538;
  assign n32535 = n32539 & n239;
  assign n32533 = ~n32546;
  assign n32543 = ~n32554;
  assign n32540 = n32558 & n32559;
  assign n29038 = n32571 ^ n32572;
  assign n32579 = ~n32587;
  assign n32071 = ~n30735;
  assign n32479 = n32515 & n32516;
  assign n32517 = n32533 & n32534;
  assign n32498 = ~n32535;
  assign n32526 = n32540 ^ n32541;
  assign n32542 = ~n32540;
  assign n31451 = n29038 ^ n30458;
  assign n29074 = ~n29038;
  assign n32565 = n32579 & n32580;
  assign n32482 = ~n32479;
  assign n32496 = n32517 ^ n32518;
  assign n32484 = n32526 ^ n32527;
  assign n32519 = ~n32517;
  assign n32489 = n31451 ^ n31427;
  assign n32536 = n32542 & n32543;
  assign n32563 = n32565 & n30326;
  assign n32562 = ~n32565;
  assign n32480 = n239 ^ n32496;
  assign n32502 = n32484 & n238;
  assign n32508 = n32519 & n32520;
  assign n32501 = ~n32484;
  assign n32521 = n32489 & n32504;
  assign n32522 = ~n32489;
  assign n32528 = ~n32536;
  assign n32555 = n32562 & n30388;
  assign n32545 = ~n32563;
  assign n32040 = n32479 ^ n32480;
  assign n32481 = ~n32480;
  assign n32499 = n32501 & n19483;
  assign n32466 = ~n32502;
  assign n32497 = ~n32508;
  assign n32506 = ~n32521;
  assign n32509 = n32522 & n32523;
  assign n32503 = n32528 & n32529;
  assign n32544 = n32545 & n32547;
  assign n32531 = ~n32555;
  assign n30663 = ~n32040;
  assign n32448 = n32481 & n32482;
  assign n32483 = n32497 & n32498;
  assign n32486 = ~n32499;
  assign n32488 = n32503 ^ n32504;
  assign n32491 = ~n32509;
  assign n32505 = ~n32503;
  assign n32530 = ~n32544;
  assign n32537 = n32531 & n32545;
  assign n32464 = n32483 ^ n32484;
  assign n32451 = n32488 ^ n32489;
  assign n32485 = ~n32483;
  assign n32500 = n32505 & n32506;
  assign n32510 = n32530 & n32531;
  assign n32524 = ~n32537;
  assign n32449 = n238 ^ n32464;
  assign n32471 = n32451 & n19432;
  assign n32475 = n32485 & n32486;
  assign n32472 = ~n32451;
  assign n32490 = ~n32500;
  assign n32492 = n32510 ^ n30269;
  assign n29036 = n32524 ^ n32525;
  assign n32511 = ~n32510;
  assign n30627 = n32448 ^ n32449;
  assign n32414 = n32449 & n32448;
  assign n32452 = ~n32471;
  assign n32467 = n32472 & n237;
  assign n32465 = ~n32475;
  assign n32487 = n32490 & n32491;
  assign n28965 = n32492 ^ n32493;
  assign n31387 = n29036 ^ n30388;
  assign n32507 = n32511 & n32512;
  assign n29003 = ~n29036;
  assign n31952 = ~n30627;
  assign n32424 = ~n32414;
  assign n32450 = n32465 & n32466;
  assign n32433 = ~n32467;
  assign n32458 = ~n32487;
  assign n32455 = n31387 ^ n31330;
  assign n28994 = ~n28965;
  assign n32494 = ~n32507;
  assign n32431 = n32450 ^ n32451;
  assign n32453 = ~n32450;
  assign n32454 = n32458 ^ n32468;
  assign n32470 = n32455 & n32473;
  assign n31344 = n28994 ^ n30233;
  assign n32469 = ~n32455;
  assign n32476 = n32494 & n32495;
  assign n32415 = n237 ^ n32431;
  assign n32443 = n32452 & n32453;
  assign n32417 = n32454 ^ n32455;
  assign n32403 = n31344 ^ n31289;
  assign n32459 = n32469 & n32468;
  assign n32457 = ~n32470;
  assign n32461 = n32476 ^ n30160;
  assign n32477 = ~n32476;
  assign n30554 = n32414 ^ n32415;
  assign n32383 = n32415 & n32424;
  assign n32434 = n32417 & n19414;
  assign n32432 = ~n32443;
  assign n32438 = n32403 & n32444;
  assign n32435 = ~n32417;
  assign n32439 = ~n32403;
  assign n32456 = n32457 & n32458;
  assign n32441 = ~n32459;
  assign n28927 = n32460 ^ n32461;
  assign n32474 = n32477 & n32478;
  assign n31884 = ~n30554;
  assign n32386 = ~n32383;
  assign n32416 = n32432 & n32433;
  assign n32419 = ~n32434;
  assign n32426 = n32435 & n236;
  assign n32405 = ~n32438;
  assign n32436 = n32439 & n32423;
  assign n31304 = n28927 ^ n30197;
  assign n32440 = ~n32456;
  assign n28956 = ~n28927;
  assign n32462 = ~n32474;
  assign n32399 = n32416 ^ n32417;
  assign n32418 = ~n32416;
  assign n32401 = ~n32426;
  assign n32368 = n31304 ^ n31292;
  assign n32425 = ~n32436;
  assign n32437 = n32440 & n32441;
  assign n32445 = n32462 & n32463;
  assign n32384 = n236 ^ n32399;
  assign n32408 = n32418 & n32419;
  assign n32410 = n32368 & n32420;
  assign n32409 = ~n32368;
  assign n32422 = ~n32437;
  assign n32427 = n32445 ^ n30091;
  assign n32446 = ~n32445;
  assign n30435 = n32383 ^ n32384;
  assign n32385 = ~n32384;
  assign n32400 = ~n32408;
  assign n32406 = n32409 & n32391;
  assign n32372 = ~n32410;
  assign n32402 = n32422 ^ n32423;
  assign n32421 = n32425 & n32422;
  assign n28885 = n32427 ^ n32428;
  assign n32442 = n32446 & n32447;
  assign n31818 = ~n30435;
  assign n32336 = n32385 & n32386;
  assign n32394 = n32400 & n32401;
  assign n32377 = n32402 ^ n32403;
  assign n32393 = ~n32406;
  assign n32404 = ~n32421;
  assign n28917 = ~n28885;
  assign n32429 = ~n32442;
  assign n32339 = ~n32336;
  assign n32387 = n32377 & n19360;
  assign n32370 = ~n32394;
  assign n32388 = ~n32377;
  assign n32390 = n32404 & n32405;
  assign n31263 = n30134 ^ n28917;
  assign n32411 = n32429 & n32430;
  assign n32359 = n32370 ^ n32377;
  assign n32369 = ~n32387;
  assign n32378 = n32388 & n235;
  assign n32367 = n32390 ^ n32391;
  assign n32330 = n31263 ^ n31251;
  assign n32392 = ~n32390;
  assign n32395 = n32411 ^ n30040;
  assign n32412 = ~n32411;
  assign n32337 = n235 ^ n32359;
  assign n32327 = n32367 ^ n32368;
  assign n32364 = n32369 & n32370;
  assign n32375 = n32330 & n32355;
  assign n32353 = ~n32378;
  assign n32373 = ~n32330;
  assign n32389 = n32392 & n32393;
  assign n28875 = n32395 ^ n32396;
  assign n32407 = n32412 & n32413;
  assign n30357 = n32336 ^ n32337;
  assign n32338 = ~n32337;
  assign n32351 = n32327 & n234;
  assign n32350 = ~n32327;
  assign n32352 = ~n32364;
  assign n32365 = n32373 & n32374;
  assign n32333 = ~n32375;
  assign n31216 = n28875 ^ n30040;
  assign n32371 = ~n32389;
  assign n28843 = ~n28875;
  assign n32397 = ~n32407;
  assign n31740 = ~n30357;
  assign n32287 = n32338 & n32339;
  assign n32347 = n32350 & n19316;
  assign n32313 = ~n32351;
  assign n32348 = n32352 & n32353;
  assign n32295 = n31216 ^ n31193;
  assign n32357 = ~n32365;
  assign n32354 = n32371 & n32372;
  assign n32379 = n32397 & n32398;
  assign n32329 = ~n32347;
  assign n32326 = ~n32348;
  assign n32340 = n32295 & n32317;
  assign n32331 = n32354 ^ n32355;
  assign n32341 = ~n32295;
  assign n32356 = ~n32354;
  assign n28789 = n32379 ^ n32380;
  assign n32381 = ~n32379;
  assign n32308 = n32326 ^ n32327;
  assign n32325 = n32329 & n32326;
  assign n32291 = n32330 ^ n32331;
  assign n32319 = ~n32340;
  assign n32334 = n32341 & n32342;
  assign n32349 = n32356 & n32357;
  assign n31194 = n29983 ^ n28789;
  assign n32361 = n28789 & n32366;
  assign n28858 = ~n28789;
  assign n32376 = n32381 & n32382;
  assign n32288 = n234 ^ n32308;
  assign n32314 = n32291 & n19279;
  assign n32312 = ~n32325;
  assign n32315 = ~n32291;
  assign n32297 = ~n32334;
  assign n32280 = n31194 ^ n31077;
  assign n32332 = ~n32349;
  assign n32358 = n28858 & n32360;
  assign n31196 = ~n32361;
  assign n32362 = ~n32376;
  assign n30280 = n32287 ^ n32288;
  assign n32253 = n32288 & n32287;
  assign n32290 = n32312 & n32313;
  assign n32292 = ~n32314;
  assign n32309 = n32315 & n233;
  assign n32322 = n32280 & n32328;
  assign n32316 = n32332 & n32333;
  assign n32321 = ~n32280;
  assign n31220 = ~n32358;
  assign n32343 = n32362 & n32363;
  assign n31680 = ~n30280;
  assign n32256 = ~n32253;
  assign n32274 = n32290 ^ n32291;
  assign n32293 = ~n32290;
  assign n32276 = ~n32309;
  assign n32294 = n32316 ^ n32317;
  assign n32320 = n32321 & n32262;
  assign n32282 = ~n32322;
  assign n32318 = ~n32316;
  assign n31217 = n31220 & n31196;
  assign n31125 = n32343 ^ n32344;
  assign n32345 = ~n32343;
  assign n32254 = n233 ^ n32274;
  assign n32289 = n32292 & n32293;
  assign n32258 = n32294 ^ n32295;
  assign n32310 = n32318 & n32319;
  assign n32264 = ~n32320;
  assign n32245 = n31125 ^ n31011;
  assign n28750 = n31125 ^ n29891;
  assign n32335 = n32345 & n32346;
  assign n30204 = n32253 ^ n32254;
  assign n32255 = ~n32254;
  assign n32277 = n32258 & n19255;
  assign n32275 = ~n32289;
  assign n32278 = ~n32258;
  assign n32296 = ~n32310;
  assign n32302 = n32245 & n32311;
  assign n32303 = n28750 & n31171;
  assign n32301 = ~n32245;
  assign n28798 = ~n28750;
  assign n32323 = ~n32335;
  assign n31612 = ~n30204;
  assign n31566 = n32255 & n32256;
  assign n32257 = n32275 & n32276;
  assign n32259 = ~n32277;
  assign n32271 = n32278 & n232;
  assign n32279 = n32296 & n32297;
  assign n32298 = n32301 & n32222;
  assign n32247 = ~n32302;
  assign n31173 = ~n32303;
  assign n32299 = n28798 & n32304;
  assign n32305 = n32323 & n32324;
  assign n32228 = ~n31566;
  assign n32239 = n32257 ^ n32258;
  assign n32260 = ~n32257;
  assign n32241 = ~n32271;
  assign n32261 = n32279 ^ n32280;
  assign n32281 = ~n32279;
  assign n32224 = ~n32298;
  assign n31145 = ~n32299;
  assign n32284 = n32305 ^ n29876;
  assign n32306 = ~n32305;
  assign n31532 = n232 ^ n32239;
  assign n32252 = n32259 & n32260;
  assign n32204 = n32261 ^ n32262;
  assign n32272 = n32281 & n32282;
  assign n28711 = n32283 ^ n32284;
  assign n32300 = n32306 & n32307;
  assign n32180 = n31532 & n32228;
  assign n32243 = n32204 & n247;
  assign n32240 = ~n32252;
  assign n32242 = ~n32204;
  assign n31069 = n29876 ^ n28711;
  assign n32263 = ~n32272;
  assign n32267 = n28711 & n32273;
  assign n28759 = ~n28711;
  assign n32285 = ~n32300;
  assign n32192 = ~n32180;
  assign n32218 = n32240 & n32241;
  assign n32236 = n32242 & n19197;
  assign n32206 = ~n32243;
  assign n32210 = n31069 ^ n30937;
  assign n32244 = n32263 & n32264;
  assign n31099 = ~n32267;
  assign n32265 = n28759 & n31127;
  assign n32268 = n32285 & n32286;
  assign n32203 = n247 ^ n32218;
  assign n32220 = ~n32218;
  assign n32219 = ~n32236;
  assign n32230 = n32210 & n32237;
  assign n32221 = n32244 ^ n32245;
  assign n32229 = ~n32210;
  assign n32246 = ~n32244;
  assign n31129 = ~n32265;
  assign n32248 = n32268 ^ n29862;
  assign n32269 = ~n32268;
  assign n32181 = n32203 ^ n32204;
  assign n32217 = n32219 & n32220;
  assign n32166 = n32221 ^ n32222;
  assign n32225 = n32229 & n32186;
  assign n32212 = ~n32230;
  assign n32238 = n32246 & n32247;
  assign n28722 = n32248 ^ n32249;
  assign n32266 = n32269 & n32270;
  assign n29402 = n32180 ^ n32181;
  assign n32142 = n32181 & n32192;
  assign n32208 = n32166 & n246;
  assign n32205 = ~n32217;
  assign n32207 = ~n32166;
  assign n32188 = ~n32225;
  assign n31004 = n28722 ^ n29823;
  assign n32223 = ~n32238;
  assign n32231 = n28722 & n31037;
  assign n28690 = ~n28722;
  assign n32250 = ~n32266;
  assign n32154 = n31268 ^ n29402;
  assign n32141 = n32164 ^ n29402;
  assign n28460 = n29400 ^ n29402;
  assign n32073 = n29402 & n29400;
  assign n32182 = n32205 & n32206;
  assign n32200 = n32207 & n19179;
  assign n32168 = ~n32208;
  assign n32149 = n31004 ^ n30908;
  assign n32209 = n32223 & n32224;
  assign n31039 = ~n32231;
  assign n32226 = n28690 & n32232;
  assign n32233 = n32250 & n32251;
  assign n29777 = n327 ^ n32141;
  assign n32015 = n32154 & n32155;
  assign n31886 = n32141 & n327;
  assign n32165 = n246 ^ n32182;
  assign n32183 = ~n32182;
  assign n32184 = ~n32200;
  assign n32195 = n32149 & n32172;
  assign n32185 = n32209 ^ n32210;
  assign n32193 = ~n32149;
  assign n32211 = ~n32209;
  assign n31072 = ~n32226;
  assign n32213 = n32233 ^ n29789;
  assign n32234 = ~n32233;
  assign n32134 = n32015 & n31985;
  assign n30700 = ~n29777;
  assign n32132 = ~n32015;
  assign n32143 = n32165 ^ n32166;
  assign n32179 = n32183 & n32184;
  assign n32145 = n32185 ^ n32186;
  assign n32189 = n32193 & n32194;
  assign n32174 = ~n32195;
  assign n32201 = n32211 & n32212;
  assign n28651 = n32213 ^ n32214;
  assign n32227 = n32234 & n32235;
  assign n32120 = n32132 & n32133;
  assign n32004 = ~n32134;
  assign n32135 = n32142 ^ n32143;
  assign n32095 = n32143 & n32142;
  assign n32170 = n32145 & n245;
  assign n32167 = ~n32179;
  assign n32169 = ~n32145;
  assign n32151 = ~n32189;
  assign n30931 = n29835 ^ n28651;
  assign n32187 = ~n32201;
  assign n32196 = n28651 & n32202;
  assign n28688 = ~n28651;
  assign n32215 = ~n32227;
  assign n32031 = ~n32120;
  assign n32122 = n32135 & n29384;
  assign n32121 = ~n32135;
  assign n32098 = ~n32095;
  assign n32144 = n32167 & n32168;
  assign n32161 = n32169 & n19125;
  assign n32125 = ~n32170;
  assign n32104 = n30931 ^ n30839;
  assign n32171 = n32187 & n32188;
  assign n31007 = ~n32196;
  assign n32190 = n28688 & n30964;
  assign n32197 = n32215 & n32216;
  assign n32116 = n32121 & n29335;
  assign n32094 = ~n32122;
  assign n32123 = n32144 ^ n32145;
  assign n32146 = ~n32144;
  assign n32147 = ~n32161;
  assign n32156 = n32104 & n32162;
  assign n32148 = n32171 ^ n32172;
  assign n32157 = ~n32104;
  assign n32173 = ~n32171;
  assign n30967 = ~n32190;
  assign n32176 = n32197 ^ n29798;
  assign n32198 = ~n32197;
  assign n32093 = n32094 & n32073;
  assign n32086 = ~n32116;
  assign n32096 = n245 ^ n32123;
  assign n32140 = n32146 & n32147;
  assign n32100 = n32148 ^ n32149;
  assign n32106 = ~n32156;
  assign n32152 = n32157 & n32129;
  assign n32163 = n32173 & n32174;
  assign n28613 = n32175 ^ n32176;
  assign n32191 = n32198 & n32199;
  assign n32085 = ~n32093;
  assign n32072 = n32086 & n32094;
  assign n32033 = n32095 ^ n32096;
  assign n32097 = ~n32096;
  assign n32126 = n32100 & n19082;
  assign n32124 = ~n32140;
  assign n32127 = ~n32100;
  assign n32131 = ~n32152;
  assign n32150 = ~n32163;
  assign n28649 = ~n28613;
  assign n32177 = ~n32191;
  assign n28327 = n32072 ^ n32073;
  assign n32059 = n32085 & n32086;
  assign n32074 = n32033 & n29324;
  assign n32075 = ~n32033;
  assign n32044 = n32097 & n32098;
  assign n32099 = n32124 & n32125;
  assign n32102 = ~n32126;
  assign n32117 = n32127 & n244;
  assign n32128 = n32150 & n32151;
  assign n30815 = n28649 ^ n29798;
  assign n32158 = n32177 & n32178;
  assign n32016 = n28327 ^ n32041;
  assign n32032 = n32059 ^ n29332;
  assign n28307 = ~n28327;
  assign n32042 = ~n32059;
  assign n32019 = ~n32074;
  assign n32067 = n32075 & n29332;
  assign n32047 = ~n32044;
  assign n32076 = n32099 ^ n32100;
  assign n32101 = ~n32099;
  assign n32078 = ~n32117;
  assign n32103 = n32128 ^ n32129;
  assign n32053 = n30815 ^ n30793;
  assign n32130 = ~n32128;
  assign n32137 = n32158 ^ n29713;
  assign n32159 = ~n32158;
  assign n31984 = n32015 ^ n32016;
  assign n32017 = n32016 & n32031;
  assign n28213 = n32032 ^ n32033;
  assign n32043 = ~n32067;
  assign n32045 = n244 ^ n32076;
  assign n32091 = n32101 & n32102;
  assign n32049 = n32103 ^ n32104;
  assign n32108 = n32053 & n32111;
  assign n32107 = ~n32053;
  assign n32118 = n32130 & n32131;
  assign n28611 = n32136 ^ n32137;
  assign n32153 = n32159 & n32160;
  assign n31972 = n31984 ^ n31985;
  assign n31920 = n32002 ^ n28213;
  assign n32003 = ~n32017;
  assign n28249 = ~n28213;
  assign n32038 = n32042 & n32043;
  assign n32034 = n32044 ^ n32045;
  assign n32046 = ~n32045;
  assign n32080 = n32049 & n243;
  assign n32077 = ~n32091;
  assign n32079 = ~n32049;
  assign n32092 = n32107 & n32082;
  assign n32055 = ~n32108;
  assign n30769 = n29713 ^ n28611;
  assign n32105 = ~n32118;
  assign n32112 = n28611 & n32119;
  assign n28573 = ~n28611;
  assign n32138 = ~n32153;
  assign n31954 = n31972 & n326;
  assign n31973 = n31920 & n31956;
  assign n31953 = ~n31972;
  assign n31974 = ~n31920;
  assign n31986 = n32003 & n32004;
  assign n32020 = n32034 & n29290;
  assign n32018 = ~n32038;
  assign n31957 = ~n32034;
  assign n31990 = n32046 & n32047;
  assign n32048 = n32077 & n32078;
  assign n32068 = n32079 & n19042;
  assign n32023 = ~n32080;
  assign n31997 = n30769 ^ n30743;
  assign n32084 = ~n32092;
  assign n32081 = n32105 & n32106;
  assign n32109 = n28573 & n30805;
  assign n30807 = ~n32112;
  assign n32113 = n32138 & n32139;
  assign n31948 = n31953 & n13593;
  assign n31888 = ~n31954;
  assign n31909 = ~n31973;
  assign n31955 = n31974 & n31975;
  assign n31940 = ~n31986;
  assign n31987 = n32018 & n32019;
  assign n32012 = n31957 & n29300;
  assign n31989 = ~n32020;
  assign n32021 = n32048 ^ n32049;
  assign n32050 = ~n32048;
  assign n32051 = ~n32068;
  assign n32061 = n31997 & n32069;
  assign n32052 = n32081 ^ n32082;
  assign n32060 = ~n31997;
  assign n32083 = ~n32081;
  assign n30844 = ~n32109;
  assign n32088 = n32113 ^ n29673;
  assign n32114 = ~n32113;
  assign n31918 = ~n31948;
  assign n31939 = ~n31955;
  assign n31919 = n31940 ^ n31956;
  assign n31958 = n31987 ^ n29290;
  assign n31988 = ~n31987;
  assign n31960 = ~n32012;
  assign n31991 = n243 ^ n32021;
  assign n32039 = n32050 & n32051;
  assign n31993 = n32052 ^ n32053;
  assign n32056 = n32060 & n32027;
  assign n31999 = ~n32061;
  assign n32070 = n32083 & n32084;
  assign n28530 = n32087 ^ n32088;
  assign n32110 = n32114 & n32115;
  assign n31915 = n31918 & n31886;
  assign n31885 = n31918 & n31888;
  assign n31850 = n31919 ^ n31920;
  assign n31921 = n31939 & n31940;
  assign n28158 = n31957 ^ n31958;
  assign n31981 = n31988 & n31989;
  assign n31976 = n31990 ^ n31991;
  assign n31926 = n31991 & n31990;
  assign n32025 = n31993 & n242;
  assign n32022 = ~n32039;
  assign n32024 = ~n31993;
  assign n32029 = ~n32056;
  assign n30698 = n28530 ^ n29673;
  assign n32054 = ~n32070;
  assign n32062 = n28530 & n32071;
  assign n28564 = ~n28530;
  assign n32089 = ~n32110;
  assign n29742 = n31885 ^ n31886;
  assign n31890 = n31850 & n325;
  assign n31887 = ~n31915;
  assign n31889 = ~n31850;
  assign n31908 = ~n31921;
  assign n31840 = n31922 ^ n28158;
  assign n28192 = ~n28158;
  assign n31961 = n31976 & n29256;
  assign n31959 = ~n31981;
  assign n31894 = ~n31976;
  assign n31992 = n32022 & n32023;
  assign n32013 = n32024 & n19000;
  assign n31964 = ~n32025;
  assign n31932 = n30698 ^ n30597;
  assign n32026 = n32054 & n32055;
  assign n30773 = ~n32062;
  assign n32057 = n28564 & n30735;
  assign n32064 = n32089 & n32090;
  assign n30624 = ~n29742;
  assign n31849 = n31887 & n31888;
  assign n31879 = n31889 & n13543;
  assign n31821 = ~n31890;
  assign n31873 = n31908 & n31909;
  assign n31892 = n31840 & n31910;
  assign n31891 = ~n31840;
  assign n31923 = n31959 & n31960;
  assign n31924 = ~n31961;
  assign n31949 = n31894 & n29272;
  assign n31962 = n31992 ^ n31993;
  assign n31994 = ~n31992;
  assign n31995 = ~n32013;
  assign n32005 = n31932 & n31968;
  assign n31996 = n32026 ^ n32027;
  assign n32006 = ~n31932;
  assign n32028 = ~n32026;
  assign n30738 = ~n32057;
  assign n28546 = n32063 ^ n32064;
  assign n32065 = ~n32064;
  assign n31819 = n31849 ^ n31850;
  assign n31839 = n31873 ^ n31874;
  assign n31851 = ~n31849;
  assign n31852 = ~n31879;
  assign n31853 = ~n31873;
  assign n31880 = n31891 & n31874;
  assign n31823 = ~n31892;
  assign n31893 = n31923 ^ n29256;
  assign n31925 = ~n31923;
  assign n31896 = ~n31949;
  assign n31927 = n242 ^ n31962;
  assign n31982 = n31994 & n31995;
  assign n31929 = n31996 ^ n31997;
  assign n31935 = ~n32005;
  assign n32000 = n32006 & n32007;
  assign n32014 = n32028 & n32029;
  assign n30623 = n29620 ^ n28546;
  assign n32035 = n28546 & n32040;
  assign n28476 = ~n28546;
  assign n32058 = n32065 & n32066;
  assign n29725 = n325 ^ n31819;
  assign n31781 = n31839 ^ n31840;
  assign n31845 = n31851 & n31852;
  assign n31854 = ~n31880;
  assign n28135 = n31893 ^ n31894;
  assign n31916 = n31924 & n31925;
  assign n31824 = n31926 ^ n31927;
  assign n31859 = n31927 & n31926;
  assign n31966 = n31929 & n241;
  assign n31963 = ~n31982;
  assign n31965 = ~n31929;
  assign n31970 = ~n32000;
  assign n31905 = n30623 ^ n30483;
  assign n31998 = ~n32014;
  assign n30703 = ~n32035;
  assign n32030 = n28476 & n30663;
  assign n32036 = ~n32058;
  assign n31807 = n31781 & n324;
  assign n30564 = ~n29725;
  assign n31806 = ~n31781;
  assign n31820 = ~n31845;
  assign n31846 = n31853 & n31854;
  assign n31752 = n28135 ^ n31855;
  assign n28105 = ~n28135;
  assign n31897 = n31824 & n29215;
  assign n31895 = ~n31916;
  assign n31898 = ~n31824;
  assign n31862 = ~n31859;
  assign n31928 = n31963 & n31964;
  assign n31950 = n31965 & n18956;
  assign n31901 = ~n31966;
  assign n31978 = n31905 & n31983;
  assign n31967 = n31998 & n31999;
  assign n31977 = ~n31905;
  assign n30666 = ~n32030;
  assign n32008 = n32036 & n32037;
  assign n31782 = n31806 & n13481;
  assign n31735 = ~n31807;
  assign n31780 = n31820 & n31821;
  assign n31822 = ~n31846;
  assign n31856 = n31895 & n31896;
  assign n31857 = ~n31897;
  assign n31881 = n31898 & n29224;
  assign n31899 = n31928 ^ n31929;
  assign n31930 = ~n31928;
  assign n31931 = ~n31950;
  assign n31933 = n31967 ^ n31968;
  assign n31971 = n31977 & n31868;
  assign n31907 = ~n31978;
  assign n31969 = ~n31967;
  assign n30551 = n32008 ^ n32009;
  assign n32010 = ~n32008;
  assign n31749 = n31780 ^ n31781;
  assign n31770 = ~n31782;
  assign n31771 = ~n31780;
  assign n31783 = n31822 & n31823;
  assign n31825 = n31856 ^ n29224;
  assign n31858 = ~n31856;
  assign n31827 = ~n31881;
  assign n31860 = n241 ^ n31899;
  assign n31917 = n31930 & n31931;
  assign n31864 = n31932 ^ n31933;
  assign n31951 = n31969 & n31970;
  assign n31870 = ~n31971;
  assign n31836 = n30551 ^ n30411;
  assign n28428 = n30551 ^ n29685;
  assign n32001 = n32010 & n32011;
  assign n29687 = n324 ^ n31749;
  assign n31750 = n31770 & n31771;
  assign n31751 = n31783 ^ n31784;
  assign n31787 = n31783 & n31784;
  assign n31785 = ~n31783;
  assign n28093 = n31824 ^ n31825;
  assign n31847 = n31857 & n31858;
  assign n31755 = n31859 ^ n31860;
  assign n31861 = ~n31860;
  assign n31902 = n31864 & n18899;
  assign n31900 = ~n31917;
  assign n31903 = ~n31864;
  assign n31934 = ~n31951;
  assign n31943 = n31836 & n31800;
  assign n31944 = n28428 & n31952;
  assign n31941 = ~n31836;
  assign n28487 = ~n28428;
  assign n31979 = ~n32001;
  assign n30471 = ~n29687;
  assign n31734 = ~n31750;
  assign n31674 = n31751 ^ n31752;
  assign n31777 = n31785 & n31786;
  assign n31772 = ~n31787;
  assign n31664 = n31788 ^ n28093;
  assign n28052 = ~n28093;
  assign n31829 = n31755 & n29165;
  assign n31826 = ~n31847;
  assign n31828 = ~n31755;
  assign n31792 = n31861 & n31862;
  assign n31863 = n31900 & n31901;
  assign n31866 = ~n31902;
  assign n31882 = n31903 & n240;
  assign n31904 = n31934 & n31935;
  assign n31936 = n31941 & n31942;
  assign n31802 = ~n31943;
  assign n30589 = ~n31944;
  assign n31937 = n28487 & n30627;
  assign n31945 = n31979 & n31980;
  assign n31712 = n31734 & n31735;
  assign n31753 = n31772 & n31752;
  assign n31737 = ~n31777;
  assign n31789 = n31826 & n31827;
  assign n31814 = n31828 & n29193;
  assign n31757 = ~n31829;
  assign n31795 = ~n31792;
  assign n31830 = n31863 ^ n31864;
  assign n31865 = ~n31863;
  assign n31832 = ~n31882;
  assign n31867 = n31904 ^ n31905;
  assign n31906 = ~n31904;
  assign n31838 = ~n31936;
  assign n30629 = ~n31937;
  assign n31912 = n31945 ^ n29645;
  assign n31946 = ~n31945;
  assign n31701 = n31712 & n13439;
  assign n31681 = ~n31712;
  assign n31736 = ~n31753;
  assign n31754 = n31789 ^ n29193;
  assign n31790 = ~n31789;
  assign n31791 = ~n31814;
  assign n31793 = n240 ^ n31830;
  assign n31848 = n31865 & n31866;
  assign n31761 = n31867 ^ n31868;
  assign n31883 = n31906 & n31907;
  assign n28379 = n31911 ^ n31912;
  assign n31938 = n31946 & n31947;
  assign n31642 = n31681 ^ n31674;
  assign n31682 = n31681 & n323;
  assign n31673 = ~n31701;
  assign n31702 = n31736 & n31737;
  assign n28006 = n31754 ^ n31755;
  assign n31778 = n31790 & n31791;
  assign n31687 = n31792 ^ n31793;
  assign n31794 = ~n31793;
  assign n31834 = n31761 & n255;
  assign n31831 = ~n31848;
  assign n31833 = ~n31761;
  assign n30461 = n28379 ^ n29549;
  assign n31869 = ~n31883;
  assign n31875 = n28379 & n31884;
  assign n28450 = ~n28379;
  assign n31913 = ~n31938;
  assign n29609 = n323 ^ n31642;
  assign n31662 = n31673 & n31674;
  assign n31637 = ~n31682;
  assign n31663 = n31702 ^ n31703;
  assign n31707 = n31702 & n31703;
  assign n31704 = ~n31702;
  assign n31571 = n31715 ^ n28006;
  assign n28034 = ~n28006;
  assign n31758 = n31687 & n29141;
  assign n31756 = ~n31778;
  assign n31759 = ~n31687;
  assign n31719 = n31794 & n31795;
  assign n31796 = n31831 & n31832;
  assign n31815 = n31833 & n18888;
  assign n31763 = ~n31834;
  assign n31767 = n30461 ^ n30338;
  assign n31835 = n31869 & n31870;
  assign n30513 = ~n31875;
  assign n31871 = n28450 & n30554;
  assign n31876 = n31913 & n31914;
  assign n29629 = ~n29609;
  assign n31636 = ~n31662;
  assign n31578 = n31663 ^ n31664;
  assign n31683 = n31704 & n31705;
  assign n31684 = n31571 & n31706;
  assign n31675 = ~n31707;
  assign n31685 = ~n31571;
  assign n31716 = n31756 & n31757;
  assign n31717 = ~n31758;
  assign n31745 = n31759 & n29169;
  assign n31722 = ~n31719;
  assign n31760 = n255 ^ n31796;
  assign n31797 = ~n31796;
  assign n31798 = ~n31815;
  assign n31809 = n31767 & n31816;
  assign n31799 = n31835 ^ n31836;
  assign n31808 = ~n31767;
  assign n31837 = ~n31835;
  assign n30556 = ~n31871;
  assign n31842 = n31876 ^ n29530;
  assign n31877 = ~n31876;
  assign n31613 = n31636 & n31637;
  assign n31665 = n31675 & n31664;
  assign n31639 = ~n31683;
  assign n31573 = ~n31684;
  assign n31676 = n31685 & n31605;
  assign n31686 = n31716 ^ n29169;
  assign n31718 = ~n31716;
  assign n31689 = ~n31745;
  assign n31720 = n31760 ^ n31761;
  assign n31779 = n31797 & n31798;
  assign n31724 = n31799 ^ n31800;
  assign n31803 = n31808 & n31728;
  assign n31769 = ~n31809;
  assign n31817 = n31837 & n31838;
  assign n28386 = n31841 ^ n31842;
  assign n31872 = n31877 & n31878;
  assign n31603 = n31613 & n13411;
  assign n31596 = ~n31613;
  assign n31638 = ~n31665;
  assign n31607 = ~n31676;
  assign n27968 = n31686 ^ n31687;
  assign n31713 = n31717 & n31718;
  assign n31618 = n31719 ^ n31720;
  assign n31721 = ~n31720;
  assign n31764 = n31724 & n18839;
  assign n31762 = ~n31779;
  assign n31765 = ~n31724;
  assign n31730 = ~n31803;
  assign n30395 = n28386 ^ n29554;
  assign n31801 = ~n31817;
  assign n31810 = n28386 & n31818;
  assign n28355 = ~n28386;
  assign n31843 = ~n31872;
  assign n31568 = n31596 ^ n31578;
  assign n31597 = n31596 & n322;
  assign n31577 = ~n31603;
  assign n31604 = n31638 & n31639;
  assign n31506 = n31643 ^ n27968;
  assign n27991 = ~n27968;
  assign n31690 = n31618 & n29139;
  assign n31688 = ~n31713;
  assign n31691 = ~n31618;
  assign n31647 = n31721 & n31722;
  assign n31723 = n31762 & n31763;
  assign n31726 = ~n31764;
  assign n31746 = n31765 & n254;
  assign n31656 = n30395 ^ n30373;
  assign n31766 = n31801 & n31802;
  assign n30438 = ~n31810;
  assign n31804 = n28355 & n30435;
  assign n31811 = n31843 & n31844;
  assign n31533 = n322 ^ n31568;
  assign n31569 = n31577 & n31578;
  assign n31549 = ~n31597;
  assign n31570 = n31604 ^ n31605;
  assign n31606 = ~n31604;
  assign n31614 = n31506 & n31542;
  assign n31615 = ~n31506;
  assign n31644 = n31688 & n31689;
  assign n31620 = ~n31690;
  assign n31677 = n31691 & n29110;
  assign n31650 = ~n31647;
  assign n31692 = n31723 ^ n31724;
  assign n31725 = ~n31723;
  assign n31694 = ~n31746;
  assign n31738 = n31656 & n31747;
  assign n31727 = n31766 ^ n31767;
  assign n31739 = ~n31656;
  assign n31768 = ~n31766;
  assign n30475 = ~n31804;
  assign n31773 = n31811 ^ n29493;
  assign n31812 = ~n31811;
  assign n30318 = n31533 ^ n29609;
  assign n31534 = ~n31533;
  assign n31548 = ~n31569;
  assign n31500 = n31570 ^ n31571;
  assign n31598 = n31606 & n31607;
  assign n31544 = ~n31614;
  assign n31608 = n31615 & n31616;
  assign n31617 = n31644 ^ n29110;
  assign n31645 = ~n31644;
  assign n31646 = ~n31677;
  assign n31648 = n254 ^ n31692;
  assign n31714 = n31725 & n31726;
  assign n31652 = n31727 ^ n31728;
  assign n31658 = ~n31738;
  assign n31731 = n31739 & n31698;
  assign n31748 = n31768 & n31769;
  assign n28353 = n31773 ^ n31774;
  assign n31805 = n31812 & n31813;
  assign n29575 = ~n30318;
  assign n31449 = n31534 & n29629;
  assign n31511 = n31548 & n31549;
  assign n31572 = ~n31598;
  assign n31508 = ~n31608;
  assign n27935 = n31617 ^ n31618;
  assign n31640 = n31645 & n31646;
  assign n31631 = n31647 ^ n31648;
  assign n31649 = ~n31648;
  assign n31696 = n31652 & n253;
  assign n31693 = ~n31714;
  assign n31695 = ~n31652;
  assign n31700 = ~n31731;
  assign n30317 = n28353 ^ n29518;
  assign n31729 = ~n31748;
  assign n31741 = n28353 & n30357;
  assign n28298 = ~n28353;
  assign n31775 = ~n31805;
  assign n31480 = n31511 ^ n31500;
  assign n31513 = n31511 & n13365;
  assign n31512 = ~n31511;
  assign n31541 = n31572 & n31573;
  assign n31445 = n31579 ^ n27935;
  assign n27950 = ~n27935;
  assign n31621 = n31631 & n29076;
  assign n31619 = ~n31640;
  assign n31554 = ~n31631;
  assign n31583 = n31649 & n31650;
  assign n31651 = n31693 & n31694;
  assign n31678 = n31695 & n18788;
  assign n31624 = ~n31696;
  assign n31590 = n30317 ^ n30217;
  assign n31697 = n31729 & n31730;
  assign n31732 = n28298 & n31740;
  assign n30360 = ~n31741;
  assign n31742 = n31775 & n31776;
  assign n31450 = n321 ^ n31480;
  assign n31504 = n31512 & n321;
  assign n31499 = ~n31513;
  assign n31505 = n31541 ^ n31542;
  assign n31543 = ~n31541;
  assign n31550 = n31445 & n31473;
  assign n31551 = ~n31445;
  assign n31580 = n31619 & n31620;
  assign n31582 = ~n31621;
  assign n31609 = n31554 & n29108;
  assign n31622 = n31651 ^ n31652;
  assign n31654 = ~n31651;
  assign n31653 = ~n31678;
  assign n31668 = n31590 & n31628;
  assign n31655 = n31697 ^ n31698;
  assign n31666 = ~n31590;
  assign n31699 = ~n31697;
  assign n30398 = ~n31732;
  assign n31708 = n31742 ^ n29482;
  assign n31743 = ~n31742;
  assign n29537 = n31449 ^ n31450;
  assign n31381 = n31450 & n31449;
  assign n31481 = n31499 & n31500;
  assign n31465 = ~n31504;
  assign n31437 = n31505 ^ n31506;
  assign n31535 = n31543 & n31544;
  assign n31475 = ~n31550;
  assign n31545 = n31551 & n31552;
  assign n31553 = n31580 ^ n29076;
  assign n31581 = ~n31580;
  assign n31556 = ~n31609;
  assign n31584 = n253 ^ n31622;
  assign n31641 = n31653 & n31654;
  assign n31586 = n31655 ^ n31656;
  assign n31659 = n31666 & n31667;
  assign n31630 = ~n31668;
  assign n31679 = n31699 & n31700;
  assign n28239 = n31708 ^ n31709;
  assign n31733 = n31743 & n31744;
  assign n30259 = ~n29537;
  assign n31392 = ~n31381;
  assign n31464 = ~n31481;
  assign n31470 = n31437 & n13319;
  assign n31471 = ~n31437;
  assign n31507 = ~n31535;
  assign n31447 = ~n31545;
  assign n27924 = n31553 ^ n31554;
  assign n31574 = n31581 & n31582;
  assign n31486 = n31583 ^ n31584;
  assign n31518 = n31584 & n31583;
  assign n31626 = n31586 & n252;
  assign n31623 = ~n31641;
  assign n31625 = ~n31586;
  assign n31592 = ~n31659;
  assign n31657 = ~n31679;
  assign n31669 = n28239 & n31680;
  assign n28289 = ~n28239;
  assign n31710 = ~n31733;
  assign n31436 = n31464 & n31465;
  assign n31439 = ~n31470;
  assign n31466 = n31471 & n320;
  assign n31472 = n31507 & n31508;
  assign n31393 = n31514 ^ n27924;
  assign n27897 = ~n27924;
  assign n31555 = ~n31574;
  assign n31502 = ~n31486;
  assign n31521 = ~n31518;
  assign n31585 = n31623 & n31624;
  assign n31610 = n31625 & n18712;
  assign n31559 = ~n31626;
  assign n31627 = n31657 & n31658;
  assign n30238 = n28289 ^ n29458;
  assign n30322 = ~n31669;
  assign n31660 = n28289 & n30280;
  assign n31670 = n31710 & n31711;
  assign n31406 = n31436 ^ n31437;
  assign n31438 = ~n31436;
  assign n31408 = ~n31466;
  assign n31444 = n31472 ^ n31473;
  assign n31474 = ~n31472;
  assign n31482 = n31393 & n31418;
  assign n31483 = ~n31393;
  assign n31515 = n31555 & n31556;
  assign n31557 = n31585 ^ n31586;
  assign n31588 = ~n31585;
  assign n31587 = ~n31610;
  assign n31589 = n31627 ^ n31628;
  assign n31527 = n30238 ^ n30215;
  assign n31629 = ~n31627;
  assign n30283 = ~n31660;
  assign n31633 = n31670 ^ n29496;
  assign n31671 = ~n31670;
  assign n31382 = n320 ^ n31406;
  assign n31424 = n31438 & n31439;
  assign n31384 = n31444 ^ n31445;
  assign n31467 = n31474 & n31475;
  assign n31396 = ~n31482;
  assign n31476 = n31483 & n31484;
  assign n31485 = n31515 ^ n29074;
  assign n31517 = n31515 & n29038;
  assign n31516 = ~n31515;
  assign n31519 = n252 ^ n31557;
  assign n31575 = n31587 & n31588;
  assign n31523 = n31589 ^ n31590;
  assign n31593 = n31527 & n31599;
  assign n31594 = ~n31527;
  assign n31611 = n31629 & n31630;
  assign n28230 = n31632 ^ n31633;
  assign n31661 = n31671 & n31672;
  assign n29520 = n31381 ^ n31382;
  assign n30131 = n31382 & n31392;
  assign n31407 = ~n31424;
  assign n31415 = n31384 & n13293;
  assign n31416 = ~n31384;
  assign n31446 = ~n31467;
  assign n31420 = ~n31476;
  assign n27889 = n31485 ^ n31486;
  assign n31509 = n31516 & n29074;
  assign n31501 = ~n31517;
  assign n31412 = n31518 ^ n31519;
  assign n31520 = ~n31519;
  assign n31560 = n31523 & n18693;
  assign n31558 = ~n31575;
  assign n31561 = ~n31523;
  assign n31529 = ~n31593;
  assign n31576 = n31594 & n31563;
  assign n30155 = n28230 ^ n29496;
  assign n31591 = ~n31611;
  assign n31600 = n28230 & n31612;
  assign n28179 = ~n28230;
  assign n31634 = ~n31661;
  assign n30166 = ~n29520;
  assign n31383 = n31407 & n31408;
  assign n31386 = ~n31415;
  assign n31409 = n31416 & n335;
  assign n31417 = n31446 & n31447;
  assign n31349 = n31451 ^ n27889;
  assign n27863 = ~n27889;
  assign n31487 = n31501 & n31502;
  assign n31488 = n31412 & n29036;
  assign n31469 = ~n31509;
  assign n31489 = ~n31412;
  assign n31452 = n31520 & n31521;
  assign n31522 = n31558 & n31559;
  assign n31525 = ~n31560;
  assign n31546 = n31561 & n251;
  assign n31461 = n30155 ^ n30129;
  assign n31565 = ~n31576;
  assign n31562 = n31591 & n31592;
  assign n31595 = n28179 & n30204;
  assign n30260 = ~n31600;
  assign n31601 = n31634 & n31635;
  assign n31356 = n31383 ^ n31384;
  assign n31385 = ~n31383;
  assign n31358 = ~n31409;
  assign n31394 = n31417 ^ n31418;
  assign n31419 = ~n31417;
  assign n31425 = n31349 & n31370;
  assign n31426 = ~n31349;
  assign n31468 = ~n31487;
  assign n31414 = ~n31488;
  assign n31477 = n31489 & n29003;
  assign n31455 = ~n31452;
  assign n31490 = n31522 ^ n31523;
  assign n31524 = ~n31522;
  assign n31492 = ~n31546;
  assign n31536 = n31461 & n31496;
  assign n31526 = n31562 ^ n31563;
  assign n31537 = ~n31461;
  assign n31564 = ~n31562;
  assign n30221 = ~n31595;
  assign n29462 = n31601 ^ n31602;
  assign n30097 = n335 ^ n31356;
  assign n31375 = n31385 & n31386;
  assign n31341 = n31393 ^ n31394;
  assign n31410 = n31419 & n31420;
  assign n31372 = ~n31425;
  assign n31421 = n31426 & n31427;
  assign n31440 = n31468 & n31469;
  assign n31442 = ~n31477;
  assign n31453 = n251 ^ n31490;
  assign n31510 = n31524 & n31525;
  assign n31457 = n31526 ^ n31527;
  assign n31463 = ~n31536;
  assign n31530 = n31537 & n31538;
  assign n31547 = n31564 & n31565;
  assign n31539 = n29462 ^ n29446;
  assign n31567 = ~n29462;
  assign n31298 = n30097 & n30131;
  assign n31357 = ~n31375;
  assign n31367 = n31341 & n13253;
  assign n31368 = ~n31341;
  assign n31395 = ~n31410;
  assign n31351 = ~n31421;
  assign n31411 = n31440 ^ n29003;
  assign n31441 = ~n31440;
  assign n31443 = n31452 ^ n31453;
  assign n31454 = ~n31453;
  assign n31494 = n31457 & n250;
  assign n31491 = ~n31510;
  assign n31493 = ~n31457;
  assign n31498 = ~n31530;
  assign n30149 = n31539 ^ n31540;
  assign n31528 = ~n31547;
  assign n31531 = n31566 ^ n31567;
  assign n31340 = n31357 & n31358;
  assign n31343 = ~n31367;
  assign n31359 = n31368 & n334;
  assign n31369 = n31395 & n31396;
  assign n27853 = n31411 ^ n31412;
  assign n31428 = n31441 & n31442;
  assign n31429 = n31443 & n28965;
  assign n31363 = ~n31443;
  assign n31398 = n31454 & n31455;
  assign n31456 = n31491 & n31492;
  assign n31478 = n31493 & n18624;
  assign n31432 = ~n31494;
  assign n31405 = n30149 ^ n31503;
  assign n31495 = n31528 & n31529;
  assign n30184 = n31531 ^ n31532;
  assign n31315 = n31340 ^ n31341;
  assign n31342 = ~n31340;
  assign n31317 = ~n31359;
  assign n31348 = n31369 ^ n31370;
  assign n31371 = ~n31369;
  assign n31309 = n31387 ^ n27853;
  assign n27828 = ~n27853;
  assign n31413 = ~n31428;
  assign n31390 = ~n31429;
  assign n31422 = n31363 & n28994;
  assign n31430 = n31456 ^ n31457;
  assign n31459 = ~n31456;
  assign n31458 = ~n31478;
  assign n31460 = n31495 ^ n31496;
  assign n31497 = ~n31495;
  assign n31299 = n334 ^ n31315;
  assign n31334 = n31342 & n31343;
  assign n31301 = n31348 ^ n31349;
  assign n31360 = n31371 & n31372;
  assign n31362 = n31309 & n31373;
  assign n31361 = ~n31309;
  assign n31388 = n31413 & n31414;
  assign n31366 = ~n31422;
  assign n31399 = n250 ^ n31430;
  assign n31448 = n31458 & n31459;
  assign n31401 = n31460 ^ n31461;
  assign n31479 = n31497 & n31498;
  assign n28480 = n31298 ^ n31299;
  assign n31255 = n31299 & n31298;
  assign n31316 = ~n31334;
  assign n31327 = n31301 & n13222;
  assign n31328 = ~n31301;
  assign n31350 = ~n31360;
  assign n31352 = n31361 & n31330;
  assign n31311 = ~n31362;
  assign n31364 = n31388 ^ n28965;
  assign n31389 = ~n31388;
  assign n31391 = n31398 ^ n31399;
  assign n31353 = n31399 & n31398;
  assign n31433 = n31401 & n18560;
  assign n31431 = ~n31448;
  assign n31434 = ~n31401;
  assign n31462 = ~n31479;
  assign n31254 = n31274 ^ n28480;
  assign n31267 = n29400 ^ n28480;
  assign n27490 = n28460 ^ n28480;
  assign n31184 = n28480 & n28460;
  assign n31258 = ~n31255;
  assign n31300 = n31316 & n31317;
  assign n31303 = ~n31327;
  assign n31318 = n31328 & n333;
  assign n31329 = n31350 & n31351;
  assign n31332 = ~n31352;
  assign n27796 = n31363 ^ n31364;
  assign n31376 = n31389 & n31390;
  assign n31377 = n31391 & n28956;
  assign n31324 = ~n31391;
  assign n31400 = n31431 & n31432;
  assign n31403 = ~n31433;
  assign n31423 = n31434 & n249;
  assign n31435 = n31462 & n31463;
  assign n29302 = n423 ^ n31254;
  assign n31115 = n31267 & n31268;
  assign n30990 = n31254 & n423;
  assign n31275 = n31300 ^ n31301;
  assign n31302 = ~n31300;
  assign n31277 = ~n31318;
  assign n31308 = n31329 ^ n31330;
  assign n31331 = ~n31329;
  assign n31270 = n31344 ^ n27796;
  assign n27799 = ~n27796;
  assign n31365 = ~n31376;
  assign n31374 = n31324 & n28927;
  assign n31347 = ~n31377;
  assign n31378 = n31400 ^ n31401;
  assign n31402 = ~n31400;
  assign n31380 = ~n31423;
  assign n31404 = n248 ^ n31435;
  assign n31243 = n31115 & n31086;
  assign n30996 = ~n29302;
  assign n31241 = ~n31115;
  assign n31256 = n333 ^ n31275;
  assign n31294 = n31302 & n31303;
  assign n31260 = n31308 ^ n31309;
  assign n31319 = n31331 & n31332;
  assign n31320 = n31270 & n31289;
  assign n31321 = ~n31270;
  assign n31345 = n31365 & n31366;
  assign n31326 = ~n31374;
  assign n31354 = n249 ^ n31378;
  assign n31397 = n31402 & n31403;
  assign n31314 = n31404 ^ n31405;
  assign n31227 = n31241 & n31242;
  assign n31101 = ~n31243;
  assign n31244 = n31255 ^ n31256;
  assign n31257 = ~n31256;
  assign n31276 = ~n31294;
  assign n31287 = n31260 & n332;
  assign n31286 = ~n31260;
  assign n31310 = ~n31319;
  assign n31272 = ~n31320;
  assign n31312 = n31321 & n31322;
  assign n31323 = n31345 ^ n28956;
  assign n31346 = ~n31345;
  assign n31282 = n31353 ^ n31354;
  assign n31355 = ~n31354;
  assign n31379 = ~n31397;
  assign n31130 = ~n31227;
  assign n31228 = n31244 & n28307;
  assign n31229 = ~n31244;
  assign n31210 = n31257 & n31258;
  assign n31259 = n31276 & n31277;
  assign n31278 = n31286 & n13196;
  assign n31232 = ~n31287;
  assign n31288 = n31310 & n31311;
  assign n31291 = ~n31312;
  assign n27736 = n31323 ^ n31324;
  assign n31335 = n31346 & n31347;
  assign n31337 = n31282 & n28917;
  assign n31336 = ~n31282;
  assign n31339 = n31355 & n31353;
  assign n31338 = n31379 & n31380;
  assign n31209 = ~n31228;
  assign n31225 = n31229 & n28327;
  assign n31230 = n31259 ^ n31260;
  assign n31261 = ~n31259;
  assign n31262 = ~n31278;
  assign n31269 = n31288 ^ n31289;
  assign n31290 = ~n31288;
  assign n31222 = n31304 ^ n27736;
  assign n27768 = ~n27736;
  assign n31325 = ~n31335;
  assign n31333 = n31336 & n28885;
  assign n31285 = ~n31337;
  assign n31313 = n31338 ^ n31339;
  assign n31208 = n31209 & n31184;
  assign n31198 = ~n31225;
  assign n31211 = n332 ^ n31230;
  assign n31252 = n31261 & n31262;
  assign n31213 = n31269 ^ n31270;
  assign n31279 = n31290 & n31291;
  assign n31280 = n31222 & n31292;
  assign n31281 = ~n31222;
  assign n31238 = n31313 ^ n31314;
  assign n31305 = n31325 & n31326;
  assign n31307 = ~n31333;
  assign n31197 = ~n31208;
  assign n31183 = n31209 & n31198;
  assign n31199 = n31210 ^ n31211;
  assign n31160 = n31211 & n31210;
  assign n31231 = ~n31252;
  assign n31245 = n31213 & n13171;
  assign n31246 = ~n31213;
  assign n31271 = ~n31279;
  assign n31224 = ~n31280;
  assign n31273 = n31281 & n31248;
  assign n31295 = n31238 & n28875;
  assign n31283 = n31305 ^ n28885;
  assign n31296 = ~n31238;
  assign n31306 = ~n31305;
  assign n27434 = n31183 ^ n31184;
  assign n31174 = n31197 & n31198;
  assign n31185 = n31199 & n28249;
  assign n31147 = ~n31199;
  assign n31212 = n31231 & n31232;
  assign n31215 = ~n31245;
  assign n31233 = n31246 & n331;
  assign n31247 = n31271 & n31272;
  assign n31250 = ~n31273;
  assign n27748 = n31282 ^ n31283;
  assign n31240 = ~n31295;
  assign n31293 = n31296 & n28843;
  assign n31297 = n31306 & n31307;
  assign n29353 = n28327 ^ n27434;
  assign n31146 = n31174 ^ n28249;
  assign n27416 = ~n27434;
  assign n31176 = ~n31174;
  assign n31181 = n31147 & n28213;
  assign n31175 = ~n31185;
  assign n31186 = n31212 ^ n31213;
  assign n31214 = ~n31212;
  assign n31188 = ~n31233;
  assign n31221 = n31247 ^ n31248;
  assign n31249 = ~n31247;
  assign n31178 = n31263 ^ n27748;
  assign n27714 = ~n27748;
  assign n31266 = ~n31293;
  assign n31284 = ~n31297;
  assign n31116 = n29353 ^ n29335;
  assign n27325 = n31146 ^ n31147;
  assign n31159 = n31175 & n31176;
  assign n31149 = ~n31181;
  assign n31161 = n331 ^ n31186;
  assign n31206 = n31214 & n31215;
  assign n31164 = n31221 ^ n31222;
  assign n31234 = n31249 & n31250;
  assign n31236 = n31178 & n31251;
  assign n31235 = ~n31178;
  assign n31264 = n31284 & n31285;
  assign n31085 = n31115 ^ n31116;
  assign n31117 = n31116 & n31130;
  assign n29340 = n27325 ^ n28249;
  assign n27333 = ~n27325;
  assign n31148 = ~n31159;
  assign n31102 = n31160 ^ n31161;
  assign n31162 = ~n31161;
  assign n31187 = ~n31206;
  assign n31201 = n31164 & n330;
  assign n31200 = ~n31164;
  assign n31223 = ~n31234;
  assign n31226 = n31235 & n31203;
  assign n31180 = ~n31236;
  assign n31237 = n31264 ^ n28843;
  assign n31265 = ~n31264;
  assign n31073 = n31085 ^ n31086;
  assign n31026 = n29340 ^ n29324;
  assign n31100 = ~n31117;
  assign n31131 = n31148 & n31149;
  assign n31119 = n31162 & n31160;
  assign n31163 = n31187 & n31188;
  assign n31189 = n31200 & n13098;
  assign n31140 = ~n31201;
  assign n31202 = n31223 & n31224;
  assign n31205 = ~n31226;
  assign n27697 = n31237 ^ n31238;
  assign n31253 = n31265 & n31266;
  assign n31058 = n31073 & n422;
  assign n31075 = n31026 & n31080;
  assign n31057 = ~n31073;
  assign n31074 = ~n31026;
  assign n31087 = n31100 & n31101;
  assign n31103 = n31131 ^ n28158;
  assign n31133 = n31131 & n28192;
  assign n31132 = ~n31131;
  assign n31138 = n31163 ^ n31164;
  assign n31165 = ~n31163;
  assign n31166 = ~n31189;
  assign n31177 = n31202 ^ n31203;
  assign n31204 = ~n31202;
  assign n31135 = n31216 ^ n27697;
  assign n27676 = ~n27697;
  assign n31239 = ~n31253;
  assign n31051 = n31057 & n7609;
  assign n30992 = ~n31058;
  assign n31059 = n31074 & n31060;
  assign n31049 = ~n31075;
  assign n31050 = ~n31087;
  assign n27246 = n31102 ^ n31103;
  assign n31118 = n31132 & n28158;
  assign n31112 = ~n31133;
  assign n31120 = n330 ^ n31138;
  assign n31156 = n31165 & n31166;
  assign n31122 = n31177 ^ n31178;
  assign n31190 = n31204 & n31205;
  assign n31191 = n31135 & n31153;
  assign n31192 = ~n31135;
  assign n31218 = n31239 & n31240;
  assign n31040 = n31049 & n31050;
  assign n31024 = ~n31051;
  assign n31015 = ~n31059;
  assign n31025 = n31050 ^ n31060;
  assign n29313 = n27246 ^ n28158;
  assign n27221 = ~n27246;
  assign n31104 = n31112 & n31102;
  assign n31082 = ~n31118;
  assign n31019 = n31119 ^ n31120;
  assign n31061 = n31120 & n31119;
  assign n31139 = ~n31156;
  assign n31151 = n31122 & n329;
  assign n31150 = ~n31122;
  assign n31179 = ~n31190;
  assign n31155 = ~n31191;
  assign n31182 = n31192 & n31193;
  assign n27623 = n31217 ^ n31218;
  assign n31219 = ~n31218;
  assign n31016 = n31024 & n30990;
  assign n30989 = n31024 & n30992;
  assign n30951 = n31025 ^ n31026;
  assign n31014 = ~n31040;
  assign n30942 = n29313 ^ n29290;
  assign n31081 = ~n31104;
  assign n31088 = n31019 & n28105;
  assign n31089 = ~n31019;
  assign n31064 = ~n31061;
  assign n31121 = n31139 & n31140;
  assign n31141 = n31150 & n13075;
  assign n31092 = ~n31151;
  assign n31152 = n31179 & n31180;
  assign n31137 = ~n31182;
  assign n31108 = n31194 ^ n27623;
  assign n27686 = ~n27623;
  assign n31207 = n31219 & n31220;
  assign n29246 = n30989 ^ n30990;
  assign n30993 = n30951 & n7523;
  assign n30980 = n31014 & n31015;
  assign n30991 = ~n31016;
  assign n31009 = n30942 & n31017;
  assign n30994 = ~n30951;
  assign n31008 = ~n30942;
  assign n31052 = n31081 & n31082;
  assign n31054 = ~n31088;
  assign n31083 = n31089 & n28135;
  assign n31090 = n31121 ^ n31122;
  assign n31123 = ~n31121;
  assign n31124 = ~n31141;
  assign n31134 = n31152 ^ n31153;
  assign n31154 = ~n31152;
  assign n31167 = n31108 & n31077;
  assign n31168 = ~n31108;
  assign n31195 = ~n31207;
  assign n29273 = ~n29246;
  assign n30941 = n30980 ^ n30981;
  assign n30950 = n30991 & n30992;
  assign n30953 = ~n30993;
  assign n30982 = n30994 & n421;
  assign n30969 = ~n30980;
  assign n30995 = n31008 & n30981;
  assign n30935 = ~n31009;
  assign n31018 = n31052 ^ n28105;
  assign n31053 = ~n31052;
  assign n31021 = ~n31083;
  assign n31062 = n329 ^ n31090;
  assign n31113 = n31123 & n31124;
  assign n31066 = n31134 ^ n31135;
  assign n31142 = n31154 & n31155;
  assign n31110 = ~n31167;
  assign n31157 = n31168 & n31169;
  assign n31170 = n31195 & n31196;
  assign n30888 = n30941 ^ n30942;
  assign n30920 = n30950 ^ n30951;
  assign n30952 = ~n30950;
  assign n30922 = ~n30982;
  assign n30968 = ~n30995;
  assign n27146 = n31018 ^ n31019;
  assign n31041 = n31053 & n31054;
  assign n30945 = n31061 ^ n31062;
  assign n31063 = ~n31062;
  assign n31091 = ~n31113;
  assign n31105 = n31066 & n13017;
  assign n31106 = ~n31066;
  assign n31136 = ~n31142;
  assign n31079 = ~n31157;
  assign n31143 = n31170 ^ n31171;
  assign n31172 = ~n31170;
  assign n30913 = n30888 & n420;
  assign n30885 = n421 ^ n30920;
  assign n30912 = ~n30888;
  assign n30943 = n30952 & n30953;
  assign n30954 = n30968 & n30969;
  assign n30983 = n27146 & n30996;
  assign n27192 = ~n27146;
  assign n31020 = ~n31041;
  assign n31028 = n30945 & n28093;
  assign n31027 = ~n30945;
  assign n30997 = n31063 & n31064;
  assign n31065 = n31091 & n31092;
  assign n31068 = ~n31105;
  assign n31093 = n31106 & n328;
  assign n31107 = n31136 & n31137;
  assign n27668 = n31143 ^ n28798;
  assign n31158 = n31172 & n31173;
  assign n29228 = n30885 ^ n29246;
  assign n30901 = n30912 & n7437;
  assign n30847 = ~n30913;
  assign n30886 = ~n30885;
  assign n30921 = ~n30943;
  assign n30934 = ~n30954;
  assign n29283 = n28135 ^ n27192;
  assign n29316 = ~n30983;
  assign n30970 = n27192 & n29302;
  assign n30984 = n31020 & n31021;
  assign n31022 = n31027 & n28052;
  assign n30947 = ~n31028;
  assign n31000 = ~n30997;
  assign n31029 = n31065 ^ n31066;
  assign n31067 = ~n31065;
  assign n31031 = ~n31093;
  assign n31076 = n31107 ^ n31108;
  assign n31109 = ~n31107;
  assign n31045 = n31125 ^ n27668;
  assign n27586 = ~n27668;
  assign n31144 = ~n31158;
  assign n30856 = ~n29228;
  assign n30816 = n30886 & n29273;
  assign n30877 = ~n30901;
  assign n30887 = n30921 & n30922;
  assign n30923 = n30934 & n30935;
  assign n30859 = n29283 ^ n29272;
  assign n29305 = ~n30970;
  assign n30944 = n30984 ^ n28052;
  assign n30985 = ~n30984;
  assign n30986 = ~n31022;
  assign n30998 = n328 ^ n31029;
  assign n31055 = n31067 & n31068;
  assign n30957 = n31076 ^ n31077;
  assign n31094 = n31109 & n31110;
  assign n31096 = n31045 & n31111;
  assign n31095 = ~n31045;
  assign n31126 = n31144 & n31145;
  assign n30819 = ~n30816;
  assign n30857 = n30887 ^ n30888;
  assign n30878 = ~n30887;
  assign n30903 = n30859 & n30914;
  assign n30870 = ~n30923;
  assign n30902 = ~n30859;
  assign n27115 = n30944 ^ n30945;
  assign n30971 = n30985 & n30986;
  assign n30972 = n30997 ^ n30998;
  assign n30999 = ~n30998;
  assign n31030 = ~n31055;
  assign n31042 = n30957 & n12996;
  assign n31043 = ~n30957;
  assign n31078 = ~n31094;
  assign n31084 = n31095 & n31011;
  assign n31047 = ~n31096;
  assign n31097 = n31126 ^ n31127;
  assign n31128 = ~n31126;
  assign n30817 = n420 ^ n30857;
  assign n30868 = n30877 & n30878;
  assign n30858 = n30870 ^ n30889;
  assign n30890 = n30902 & n30889;
  assign n30832 = ~n30903;
  assign n29231 = n28093 ^ n27115;
  assign n27075 = ~n27115;
  assign n30946 = ~n30971;
  assign n30955 = n30972 & n28034;
  assign n30880 = ~n30972;
  assign n30924 = n30999 & n31000;
  assign n31001 = n31030 & n31031;
  assign n31003 = ~n31042;
  assign n31032 = n31043 & n343;
  assign n31044 = n31078 & n31079;
  assign n31013 = ~n31084;
  assign n27547 = n28711 ^ n31097;
  assign n31114 = n31128 & n31129;
  assign n29195 = n30816 ^ n30817;
  assign n30818 = ~n30817;
  assign n30809 = n30858 ^ n30859;
  assign n30846 = ~n30868;
  assign n30760 = n29231 ^ n29224;
  assign n30869 = ~n30890;
  assign n30915 = n30946 & n30947;
  assign n30917 = ~n30955;
  assign n30948 = n30880 & n28006;
  assign n30956 = n343 ^ n31001;
  assign n31002 = ~n31001;
  assign n30959 = ~n31032;
  assign n31010 = n31044 ^ n31045;
  assign n31046 = ~n31044;
  assign n30976 = n31069 ^ n27547;
  assign n27595 = ~n27547;
  assign n31098 = ~n31114;
  assign n30775 = ~n29195;
  assign n30739 = n30818 & n30819;
  assign n30820 = n30809 & n7333;
  assign n30808 = n30846 & n30847;
  assign n30821 = ~n30809;
  assign n30848 = n30760 & n30860;
  assign n30861 = n30869 & n30870;
  assign n30849 = ~n30760;
  assign n30879 = n30915 ^ n28034;
  assign n30916 = ~n30915;
  assign n30882 = ~n30948;
  assign n30925 = n30956 ^ n30957;
  assign n30987 = n31002 & n31003;
  assign n30928 = n31010 ^ n31011;
  assign n31033 = n31046 & n31047;
  assign n31035 = n30976 & n31048;
  assign n31034 = ~n30976;
  assign n31070 = n31098 & n31099;
  assign n30776 = n30808 ^ n30809;
  assign n30794 = ~n30820;
  assign n30810 = n30821 & n419;
  assign n30795 = ~n30808;
  assign n30762 = ~n30848;
  assign n30833 = n30849 & n30797;
  assign n30831 = ~n30861;
  assign n27040 = n30879 ^ n30880;
  assign n30904 = n30916 & n30917;
  assign n30812 = n30924 ^ n30925;
  assign n30926 = ~n30925;
  assign n30958 = ~n30987;
  assign n30974 = n30928 & n342;
  assign n30973 = ~n30928;
  assign n31012 = ~n31033;
  assign n31023 = n31034 & n30937;
  assign n30978 = ~n31035;
  assign n31036 = n31070 ^ n28690;
  assign n31071 = ~n31070;
  assign n30740 = n419 ^ n30776;
  assign n30783 = n30794 & n30795;
  assign n30758 = ~n30810;
  assign n30796 = n30831 & n30832;
  assign n30799 = ~n30833;
  assign n29208 = n27040 ^ n28006;
  assign n30845 = n27040 & n30856;
  assign n26984 = ~n27040;
  assign n30881 = ~n30904;
  assign n30862 = n30926 & n30924;
  assign n30927 = n30958 & n30959;
  assign n30960 = n30973 & n12940;
  assign n30893 = ~n30974;
  assign n30975 = n31012 & n31013;
  assign n30939 = ~n31023;
  assign n27565 = n31036 ^ n31037;
  assign n31056 = n31071 & n31072;
  assign n29163 = n30739 ^ n30740;
  assign n30635 = n30740 & n30739;
  assign n30757 = ~n30783;
  assign n30759 = n30796 ^ n30797;
  assign n30692 = n29208 ^ n29193;
  assign n30798 = ~n30796;
  assign n29230 = ~n30845;
  assign n30830 = n26984 & n29228;
  assign n30850 = n30881 & n30882;
  assign n30891 = n30927 ^ n30928;
  assign n30929 = ~n30927;
  assign n30930 = ~n30960;
  assign n30936 = n30975 ^ n30976;
  assign n30977 = ~n30975;
  assign n30872 = n31004 ^ n27565;
  assign n27529 = ~n27565;
  assign n31038 = ~n31056;
  assign n30675 = ~n29163;
  assign n30746 = n30757 & n30758;
  assign n30709 = n30759 ^ n30760;
  assign n30779 = n30692 & n30727;
  assign n30784 = n30798 & n30799;
  assign n30777 = ~n30692;
  assign n29242 = ~n30830;
  assign n30811 = n30850 ^ n27991;
  assign n30852 = n30850 & n27991;
  assign n30851 = ~n30850;
  assign n30863 = n342 ^ n30891;
  assign n30918 = n30929 & n30930;
  assign n30865 = n30936 ^ n30937;
  assign n30961 = n30977 & n30978;
  assign n30963 = n30872 & n30979;
  assign n30962 = ~n30872;
  assign n31005 = n31038 & n31039;
  assign n30725 = n30709 & n418;
  assign n30690 = ~n30746;
  assign n30724 = ~n30709;
  assign n30763 = n30777 & n30778;
  assign n30729 = ~n30779;
  assign n30761 = ~n30784;
  assign n26912 = n30811 ^ n30812;
  assign n30834 = n30851 & n27968;
  assign n30822 = ~n30852;
  assign n30835 = n30862 ^ n30863;
  assign n30787 = n30863 & n30862;
  assign n30892 = ~n30918;
  assign n30906 = n30865 & n341;
  assign n30905 = ~n30865;
  assign n30938 = ~n30961;
  assign n30949 = n30962 & n30908;
  assign n30874 = ~n30963;
  assign n30965 = n31005 ^ n28651;
  assign n31006 = ~n31005;
  assign n30676 = n30690 ^ n30709;
  assign n30710 = n30724 & n7273;
  assign n30652 = ~n30725;
  assign n30726 = n30761 & n30762;
  assign n30694 = ~n30763;
  assign n29176 = n26912 ^ n27968;
  assign n30774 = n26912 & n29195;
  assign n26932 = ~n26912;
  assign n30813 = n30822 & n30812;
  assign n30786 = ~n30834;
  assign n30823 = n30835 & n27950;
  assign n30714 = ~n30835;
  assign n30864 = n30892 & n30893;
  assign n30894 = n30905 & n12900;
  assign n30826 = ~n30906;
  assign n30907 = n30938 & n30939;
  assign n30910 = ~n30949;
  assign n27527 = n30964 ^ n30965;
  assign n30988 = n31006 & n31007;
  assign n30636 = n418 ^ n30676;
  assign n30689 = ~n30710;
  assign n30691 = n30726 ^ n30727;
  assign n30620 = n29176 ^ n29169;
  assign n30728 = ~n30726;
  assign n29198 = ~n30774;
  assign n30756 = n26932 & n30775;
  assign n30785 = ~n30813;
  assign n30749 = ~n30823;
  assign n30814 = n30714 & n27935;
  assign n30824 = n30864 ^ n30865;
  assign n30866 = ~n30864;
  assign n30867 = ~n30894;
  assign n30871 = n30907 ^ n30908;
  assign n30909 = ~n30907;
  assign n30801 = n30931 ^ n27527;
  assign n27484 = ~n27527;
  assign n30966 = ~n30988;
  assign n29136 = n30635 ^ n30636;
  assign n30541 = n30636 & n30635;
  assign n30677 = n30689 & n30690;
  assign n30616 = n30691 ^ n30692;
  assign n30704 = n30620 & n30711;
  assign n30712 = n30728 & n30729;
  assign n30705 = ~n30620;
  assign n29212 = ~n30756;
  assign n30747 = n30785 & n30786;
  assign n30716 = ~n30814;
  assign n30788 = n341 ^ n30824;
  assign n30853 = n30866 & n30867;
  assign n30790 = n30871 ^ n30872;
  assign n30895 = n30909 & n30910;
  assign n30896 = n30801 & n30839;
  assign n30897 = ~n30801;
  assign n30940 = n30966 & n30967;
  assign n30601 = ~n29136;
  assign n30544 = ~n30541;
  assign n30653 = n30616 & n7227;
  assign n30651 = ~n30677;
  assign n30654 = ~n30616;
  assign n30622 = ~n30704;
  assign n30695 = n30705 & n30656;
  assign n30693 = ~n30712;
  assign n30713 = n30747 ^ n27950;
  assign n30748 = ~n30747;
  assign n30764 = n30787 ^ n30788;
  assign n30717 = n30788 & n30787;
  assign n30825 = ~n30853;
  assign n30837 = n30790 & n340;
  assign n30836 = ~n30790;
  assign n30873 = ~n30895;
  assign n30841 = ~n30896;
  assign n30883 = n30897 & n30898;
  assign n30933 = n30940 & n28613;
  assign n30932 = ~n30940;
  assign n30615 = n30651 & n30652;
  assign n30618 = ~n30653;
  assign n30637 = n30654 & n417;
  assign n30655 = n30693 & n30694;
  assign n30658 = ~n30695;
  assign n26877 = n30713 ^ n30714;
  assign n30741 = n30748 & n30749;
  assign n30750 = n30764 & n27897;
  assign n30640 = ~n30764;
  assign n30789 = n30825 & n30826;
  assign n30827 = n30836 & n12857;
  assign n30753 = ~n30837;
  assign n30838 = n30873 & n30874;
  assign n30803 = ~n30883;
  assign n30919 = n30932 & n28649;
  assign n30900 = ~n30933;
  assign n30578 = n30615 ^ n30616;
  assign n30617 = ~n30615;
  assign n30580 = ~n30637;
  assign n30619 = n30655 ^ n30656;
  assign n30657 = ~n30655;
  assign n29147 = n26877 ^ n27935;
  assign n30674 = n26877 & n29163;
  assign n26832 = ~n26877;
  assign n30715 = ~n30741;
  assign n30742 = n30640 & n27924;
  assign n30680 = ~n30750;
  assign n30751 = n30789 ^ n30790;
  assign n30791 = ~n30789;
  assign n30792 = ~n30827;
  assign n30800 = n30838 ^ n30839;
  assign n30840 = ~n30838;
  assign n30899 = n30900 & n30911;
  assign n30876 = ~n30919;
  assign n30542 = n417 ^ n30578;
  assign n30602 = n30617 & n30618;
  assign n30546 = n30619 ^ n30620;
  assign n30528 = n29147 ^ n29139;
  assign n30638 = n30657 & n30658;
  assign n29167 = ~n30674;
  assign n30667 = n26832 & n30675;
  assign n30678 = n30715 & n30716;
  assign n30642 = ~n30742;
  assign n30718 = n340 ^ n30751;
  assign n30780 = n30791 & n30792;
  assign n30720 = n30800 ^ n30801;
  assign n30828 = n30840 & n30841;
  assign n30875 = ~n30899;
  assign n30884 = n30876 & n30900;
  assign n30514 = n30541 ^ n30542;
  assign n30543 = ~n30542;
  assign n30582 = n30546 & n416;
  assign n30579 = ~n30602;
  assign n30581 = ~n30546;
  assign n30605 = n30528 & n30568;
  assign n30603 = ~n30528;
  assign n30621 = ~n30638;
  assign n29180 = ~n30667;
  assign n30639 = n30678 ^ n27897;
  assign n30679 = ~n30678;
  assign n30570 = n30717 ^ n30718;
  assign n30643 = n30718 & n30717;
  assign n30752 = ~n30780;
  assign n30765 = n30720 & n12818;
  assign n30766 = ~n30720;
  assign n30802 = ~n30828;
  assign n30842 = n30875 & n30876;
  assign n30854 = ~n30884;
  assign n29102 = ~n30514;
  assign n30464 = n30543 & n30544;
  assign n30545 = n30579 & n30580;
  assign n30565 = n30581 & n7122;
  assign n30504 = ~n30582;
  assign n30591 = n30603 & n30604;
  assign n30530 = ~n30605;
  assign n30606 = n30621 & n30622;
  assign n26813 = n30639 ^ n30640;
  assign n30668 = n30679 & n30680;
  assign n30682 = n30570 & n27863;
  assign n30681 = ~n30570;
  assign n30719 = n30752 & n30753;
  assign n30722 = ~n30765;
  assign n30754 = n30766 & n339;
  assign n30767 = n30802 & n30803;
  assign n30804 = n30842 ^ n28611;
  assign n27438 = n30854 ^ n30855;
  assign n30843 = ~n30842;
  assign n30502 = n30545 ^ n30546;
  assign n30547 = ~n30545;
  assign n30548 = ~n30565;
  assign n30566 = ~n30591;
  assign n30567 = ~n30606;
  assign n29118 = n26813 ^ n27924;
  assign n30600 = n26813 & n29136;
  assign n26773 = ~n26813;
  assign n30641 = ~n30668;
  assign n30669 = n30681 & n27889;
  assign n30609 = ~n30682;
  assign n30683 = n30719 ^ n30720;
  assign n30721 = ~n30719;
  assign n30685 = ~n30754;
  assign n30730 = n30767 ^ n30768;
  assign n30744 = ~n30767;
  assign n27384 = n30804 ^ n30805;
  assign n30731 = n30815 ^ n27438;
  assign n30829 = n30843 & n30844;
  assign n27473 = ~n27438;
  assign n30465 = n416 ^ n30502;
  assign n30526 = n30547 & n30548;
  assign n30557 = n30566 & n30567;
  assign n30453 = n29118 ^ n29108;
  assign n30527 = n30567 ^ n30568;
  assign n29138 = ~n30600;
  assign n30590 = n26773 & n30601;
  assign n30607 = n30641 & n30642;
  assign n30572 = ~n30669;
  assign n30644 = n339 ^ n30683;
  assign n30706 = n30721 & n30722;
  assign n30647 = n30730 ^ n30731;
  assign n30632 = n30769 ^ n27384;
  assign n30782 = n30731 & n30793;
  assign n27426 = ~n27384;
  assign n30781 = ~n30731;
  assign n30806 = ~n30829;
  assign n29068 = n30464 ^ n30465;
  assign n30384 = n30465 & n30464;
  assign n30503 = ~n30526;
  assign n30467 = n30527 ^ n30528;
  assign n30531 = n30453 & n30549;
  assign n30529 = ~n30557;
  assign n30532 = ~n30453;
  assign n29152 = ~n30590;
  assign n30569 = n30607 ^ n27863;
  assign n30608 = ~n30607;
  assign n30494 = n30643 ^ n30644;
  assign n30645 = ~n30644;
  assign n30684 = ~n30706;
  assign n30697 = n30647 & n338;
  assign n30696 = ~n30647;
  assign n30732 = n30632 & n30743;
  assign n30733 = ~n30632;
  assign n30770 = n30781 & n30768;
  assign n30708 = ~n30782;
  assign n30771 = n30806 & n30807;
  assign n30425 = ~n29068;
  assign n30387 = ~n30384;
  assign n30466 = n30503 & n30504;
  assign n30488 = n30467 & n431;
  assign n30487 = ~n30467;
  assign n30489 = n30529 & n30530;
  assign n30457 = ~n30531;
  assign n30515 = n30532 & n30490;
  assign n26722 = n30569 ^ n30570;
  assign n30592 = n30608 & n30609;
  assign n30573 = n30645 & n30643;
  assign n30646 = n30684 & n30685;
  assign n30686 = n30696 & n12767;
  assign n30612 = ~n30697;
  assign n30634 = ~n30732;
  assign n30723 = n30733 & n30671;
  assign n30745 = ~n30770;
  assign n30736 = n30771 ^ n28530;
  assign n30772 = ~n30771;
  assign n30427 = n30466 ^ n30467;
  assign n30454 = ~n30466;
  assign n30476 = n30487 & n7117;
  assign n30419 = ~n30488;
  assign n30452 = n30489 ^ n30490;
  assign n30501 = n26722 & n30514;
  assign n30492 = ~n30489;
  assign n30491 = ~n30515;
  assign n26748 = ~n26722;
  assign n30571 = ~n30592;
  assign n30610 = n30646 ^ n30647;
  assign n30648 = ~n30646;
  assign n30649 = ~n30686;
  assign n30673 = ~n30723;
  assign n27382 = n30735 ^ n30736;
  assign n30734 = n30744 & n30745;
  assign n30755 = n30772 & n30773;
  assign n30385 = n431 ^ n30427;
  assign n30363 = n30452 ^ n30453;
  assign n30455 = ~n30476;
  assign n30477 = n30491 & n30492;
  assign n30486 = n26748 & n29102;
  assign n29121 = ~n30501;
  assign n29085 = n27889 ^ n26748;
  assign n30533 = n30571 & n30572;
  assign n30574 = n338 ^ n30610;
  assign n30630 = n30648 & n30649;
  assign n30561 = n30698 ^ n27382;
  assign n30699 = n27382 & n29777;
  assign n27320 = ~n27382;
  assign n30707 = ~n30734;
  assign n30737 = ~n30755;
  assign n29030 = n30384 ^ n30385;
  assign n30386 = ~n30385;
  assign n30417 = n30363 & n430;
  assign n30416 = ~n30363;
  assign n30439 = n30454 & n30455;
  assign n30456 = ~n30477;
  assign n30380 = n29085 ^ n29074;
  assign n29105 = ~n30486;
  assign n30493 = n30533 ^ n27828;
  assign n30535 = n30533 & n27828;
  assign n30534 = ~n30533;
  assign n30391 = n30573 ^ n30574;
  assign n30496 = n30574 & n30573;
  assign n30611 = ~n30630;
  assign n30661 = n30561 & n30597;
  assign n30659 = ~n30561;
  assign n29779 = ~n30699;
  assign n30687 = n27320 & n30700;
  assign n30670 = n30707 & n30708;
  assign n30701 = n30737 & n30738;
  assign n30349 = ~n29030;
  assign n30284 = n30386 & n30387;
  assign n30399 = n30416 & n7047;
  assign n30344 = ~n30417;
  assign n30418 = ~n30439;
  assign n30420 = n30456 & n30457;
  assign n30441 = n30380 & n30458;
  assign n30440 = ~n30380;
  assign n26706 = n30493 ^ n30494;
  assign n30516 = n30534 & n27853;
  assign n30505 = ~n30535;
  assign n30537 = n30391 & n27799;
  assign n30536 = ~n30391;
  assign n30499 = ~n30496;
  assign n30575 = n30611 & n30612;
  assign n30650 = n30659 & n30660;
  assign n30599 = ~n30661;
  assign n30631 = n30670 ^ n30671;
  assign n29801 = ~n30687;
  assign n30672 = ~n30670;
  assign n30664 = n30701 ^ n28546;
  assign n30702 = ~n30701;
  assign n30287 = ~n30284;
  assign n30378 = ~n30399;
  assign n30400 = n30418 & n30419;
  assign n30379 = n30420 ^ n30421;
  assign n30415 = n26706 & n30425;
  assign n30401 = ~n30420;
  assign n30428 = n30440 & n30421;
  assign n30365 = ~n30441;
  assign n29050 = n27853 ^ n26706;
  assign n26676 = ~n26706;
  assign n30495 = n30505 & n30494;
  assign n30469 = ~n30516;
  assign n30517 = n30536 & n27796;
  assign n30431 = ~n30537;
  assign n30558 = ~n30575;
  assign n30576 = n30631 ^ n30632;
  assign n30563 = ~n30650;
  assign n27215 = n30663 ^ n30664;
  assign n30662 = n30672 & n30673;
  assign n30688 = n30702 & n30703;
  assign n30306 = n30379 ^ n30380;
  assign n30362 = ~n30400;
  assign n29071 = ~n30415;
  assign n30290 = n29050 ^ n29036;
  assign n30402 = ~n30428;
  assign n30426 = n26676 & n29068;
  assign n30468 = ~n30495;
  assign n30393 = ~n30517;
  assign n30538 = n30575 ^ n30576;
  assign n30594 = n30576 & n337;
  assign n30593 = ~n30576;
  assign n30523 = n30623 ^ n27215;
  assign n30625 = n27215 & n29742;
  assign n27355 = ~n27215;
  assign n30633 = ~n30662;
  assign n30665 = ~n30688;
  assign n30346 = n30306 & n429;
  assign n30345 = ~n30306;
  assign n30323 = n30362 ^ n30363;
  assign n30361 = n30378 & n30362;
  assign n30381 = n30290 & n30388;
  assign n30389 = n30401 & n30402;
  assign n30382 = ~n30290;
  assign n29088 = ~n30426;
  assign n30429 = n30468 & n30469;
  assign n30497 = n337 ^ n30538;
  assign n30583 = n30593 & n12734;
  assign n30519 = ~n30594;
  assign n30585 = n30523 & n30595;
  assign n30584 = ~n30523;
  assign n30613 = n27355 & n30624;
  assign n29744 = ~n30625;
  assign n30596 = n30633 & n30634;
  assign n30626 = n30665 & n30666;
  assign n30285 = n430 ^ n30323;
  assign n30324 = n30345 & n7015;
  assign n30264 = ~n30346;
  assign n30343 = ~n30361;
  assign n30292 = ~n30381;
  assign n30366 = n30382 & n30326;
  assign n30364 = ~n30389;
  assign n30390 = n30429 ^ n27799;
  assign n30430 = ~n30429;
  assign n30313 = n30496 ^ n30497;
  assign n30498 = ~n30497;
  assign n30559 = ~n30583;
  assign n30577 = n30584 & n30483;
  assign n30525 = ~n30585;
  assign n30560 = n30596 ^ n30597;
  assign n29763 = ~n30613;
  assign n30598 = ~n30596;
  assign n30587 = n30626 ^ n30627;
  assign n30628 = ~n30626;
  assign n30261 = n30284 ^ n30285;
  assign n30286 = ~n30285;
  assign n30307 = ~n30324;
  assign n30305 = n30343 & n30344;
  assign n30325 = n30364 & n30365;
  assign n30328 = ~n30366;
  assign n26635 = n30390 ^ n30391;
  assign n30422 = n30430 & n30431;
  assign n30460 = n30313 & n27736;
  assign n30459 = ~n30313;
  assign n30403 = n30498 & n30499;
  assign n30550 = n30558 & n30559;
  assign n30479 = n30560 ^ n30561;
  assign n30485 = ~n30577;
  assign n27150 = n28428 ^ n30587;
  assign n30586 = n30598 & n30599;
  assign n30614 = n30628 & n30629;
  assign n28997 = ~n30261;
  assign n30222 = n30286 & n30287;
  assign n30262 = n30305 ^ n30306;
  assign n30308 = ~n30305;
  assign n30289 = n30325 ^ n30326;
  assign n30341 = n26635 & n30349;
  assign n30327 = ~n30325;
  assign n29014 = n27796 ^ n26635;
  assign n26666 = ~n26635;
  assign n30392 = ~n30422;
  assign n30442 = n30459 & n27768;
  assign n30315 = ~n30460;
  assign n30406 = ~n30403;
  assign n30520 = n30479 & n12647;
  assign n30518 = ~n30550;
  assign n30521 = ~n30479;
  assign n30449 = n30551 ^ n27150;
  assign n30552 = n27150 & n30564;
  assign n27307 = ~n27150;
  assign n30562 = ~n30586;
  assign n30588 = ~n30614;
  assign n30223 = n429 ^ n30262;
  assign n30225 = n30289 ^ n30290;
  assign n30288 = n30307 & n30308;
  assign n30192 = n29014 ^ n28965;
  assign n30311 = n30327 & n30328;
  assign n29055 = ~n30341;
  assign n30342 = n26666 & n29030;
  assign n30350 = n30392 & n30393;
  assign n30352 = ~n30442;
  assign n30478 = n30518 & n30519;
  assign n30481 = ~n30520;
  assign n30506 = n30521 & n336;
  assign n30509 = n30449 & n30411;
  assign n30507 = ~n30449;
  assign n29704 = ~n30552;
  assign n30539 = n27307 & n29725;
  assign n30522 = n30562 & n30563;
  assign n30553 = n30588 & n30589;
  assign n30189 = n30222 ^ n30223;
  assign n30150 = n30223 & n30222;
  assign n30244 = n30225 & n428;
  assign n30243 = ~n30225;
  assign n30263 = ~n30288;
  assign n30270 = n30192 & n30233;
  assign n30268 = ~n30192;
  assign n30291 = ~n30311;
  assign n29033 = ~n30342;
  assign n30312 = n30350 ^ n27768;
  assign n30351 = ~n30350;
  assign n30443 = n30478 ^ n30479;
  assign n30480 = ~n30478;
  assign n30445 = ~n30506;
  assign n30500 = n30507 & n30508;
  assign n30413 = ~n30509;
  assign n30482 = n30522 ^ n30523;
  assign n29727 = ~n30539;
  assign n30524 = ~n30522;
  assign n30511 = n30553 ^ n30554;
  assign n30555 = ~n30553;
  assign n28958 = ~n30189;
  assign n30230 = n30243 & n6946;
  assign n30169 = ~n30244;
  assign n30224 = n30263 & n30264;
  assign n30265 = n30268 & n30269;
  assign n30194 = ~n30270;
  assign n30271 = n30291 & n30292;
  assign n26622 = n30312 ^ n30313;
  assign n30347 = n30351 & n30352;
  assign n30404 = n336 ^ n30443;
  assign n30470 = n30480 & n30481;
  assign n30368 = n30482 ^ n30483;
  assign n30451 = ~n30500;
  assign n27079 = n30511 ^ n28450;
  assign n30510 = n30524 & n30525;
  assign n30540 = n30555 & n30556;
  assign n30186 = n30224 ^ n30225;
  assign n30205 = ~n30230;
  assign n30229 = n26622 & n28997;
  assign n30206 = ~n30224;
  assign n30231 = ~n30265;
  assign n30232 = ~n30271;
  assign n28977 = n26622 ^ n27736;
  assign n26592 = ~n26622;
  assign n30314 = ~n30347;
  assign n30235 = n30403 ^ n30404;
  assign n30405 = ~n30404;
  assign n30447 = n30368 & n351;
  assign n30444 = ~n30470;
  assign n30446 = ~n30368;
  assign n30472 = n27079 & n29687;
  assign n27237 = ~n27079;
  assign n30484 = ~n30510;
  assign n30512 = ~n30540;
  assign n30151 = n428 ^ n30186;
  assign n30190 = n30205 & n30206;
  assign n28999 = ~n30229;
  assign n30226 = n30231 & n30232;
  assign n30119 = n28977 ^ n28956;
  assign n30191 = n30232 ^ n30233;
  assign n30242 = n26592 & n30261;
  assign n30272 = n30314 & n30315;
  assign n30246 = ~n30235;
  assign n30329 = n30405 & n30406;
  assign n30407 = n30444 & n30445;
  assign n30432 = n30446 & n12617;
  assign n30370 = ~n30447;
  assign n30375 = n30461 ^ n27237;
  assign n30462 = n27237 & n30471;
  assign n29689 = ~n30472;
  assign n30448 = n30484 & n30485;
  assign n30473 = n30512 & n30513;
  assign n28921 = n30150 ^ n30151;
  assign n30065 = n30151 & n30150;
  assign n30168 = ~n30190;
  assign n30133 = n30191 ^ n30192;
  assign n30195 = n30119 & n30160;
  assign n30193 = ~n30226;
  assign n30196 = ~n30119;
  assign n29017 = ~n30242;
  assign n30234 = n30272 ^ n27714;
  assign n30274 = n30272 & n27714;
  assign n30273 = ~n30272;
  assign n30332 = ~n30329;
  assign n30367 = n351 ^ n30407;
  assign n30408 = ~n30407;
  assign n30409 = ~n30432;
  assign n30424 = n30375 & n30433;
  assign n30410 = n30448 ^ n30449;
  assign n30423 = ~n30375;
  assign n29663 = ~n30462;
  assign n30450 = ~n30448;
  assign n30436 = n30473 ^ n28386;
  assign n30474 = ~n30473;
  assign n30114 = ~n28921;
  assign n30132 = n30168 & n30169;
  assign n30158 = n30133 & n427;
  assign n30157 = ~n30133;
  assign n30159 = n30193 & n30194;
  assign n30161 = ~n30195;
  assign n30187 = n30196 & n30197;
  assign n26550 = n30234 ^ n30235;
  assign n30266 = n30273 & n27748;
  assign n30245 = ~n30274;
  assign n30330 = n30367 ^ n30368;
  assign n30394 = n30408 & n30409;
  assign n30334 = n30410 ^ n30411;
  assign n30414 = n30423 & n30338;
  assign n30377 = ~n30424;
  assign n27119 = n30435 ^ n30436;
  assign n30434 = n30450 & n30451;
  assign n30463 = n30474 & n30475;
  assign n30099 = n30132 ^ n30133;
  assign n30122 = ~n30132;
  assign n30152 = n30157 & n6920;
  assign n30089 = ~n30158;
  assign n30120 = n30159 ^ n30160;
  assign n30162 = ~n30159;
  assign n30124 = ~n30187;
  assign n30185 = n26550 & n30189;
  assign n28939 = n27748 ^ n26550;
  assign n26576 = ~n26550;
  assign n30236 = n30245 & n30246;
  assign n30208 = ~n30266;
  assign n30136 = n30329 ^ n30330;
  assign n30331 = ~n30330;
  assign n30371 = n30334 & n12503;
  assign n30369 = ~n30394;
  assign n30372 = ~n30334;
  assign n30256 = n30395 ^ n27119;
  assign n30340 = ~n30414;
  assign n27047 = ~n27119;
  assign n30412 = ~n30434;
  assign n30437 = ~n30463;
  assign n30066 = n427 ^ n30099;
  assign n30056 = n30119 ^ n30120;
  assign n30121 = ~n30152;
  assign n30153 = n30161 & n30162;
  assign n30059 = n28939 ^ n28885;
  assign n28982 = ~n30185;
  assign n30167 = n26576 & n28958;
  assign n30207 = ~n30236;
  assign n30294 = n30136 & n27697;
  assign n30293 = ~n30136;
  assign n30247 = n30331 & n30332;
  assign n30333 = n30369 & n30370;
  assign n30336 = ~n30371;
  assign n30353 = n30372 & n350;
  assign n30355 = n30256 & n30373;
  assign n30354 = ~n30256;
  assign n30374 = n30412 & n30413;
  assign n30396 = n30437 & n30438;
  assign n30036 = n30065 ^ n30066;
  assign n29996 = n30066 & n30065;
  assign n30086 = n30056 & n6878;
  assign n30087 = ~n30056;
  assign n30115 = n30121 & n30122;
  assign n30125 = n30059 & n30134;
  assign n30123 = ~n30153;
  assign n30126 = ~n30059;
  assign n28961 = ~n30167;
  assign n30170 = n30207 & n30208;
  assign n30275 = n30293 & n27676;
  assign n30138 = ~n30294;
  assign n30250 = ~n30247;
  assign n30295 = n30333 ^ n30334;
  assign n30335 = ~n30333;
  assign n30297 = ~n30353;
  assign n30348 = n30354 & n30302;
  assign n30258 = ~n30355;
  assign n30337 = n30374 ^ n30375;
  assign n30376 = ~n30374;
  assign n30358 = n30396 ^ n28298;
  assign n30397 = ~n30396;
  assign n30037 = ~n30036;
  assign n30057 = ~n30086;
  assign n30081 = n30087 & n426;
  assign n30088 = ~n30115;
  assign n30090 = n30123 & n30124;
  assign n30061 = ~n30125;
  assign n30116 = n30126 & n30091;
  assign n30135 = n30170 ^ n27676;
  assign n30171 = ~n30170;
  assign n30172 = ~n30275;
  assign n30248 = n350 ^ n30295;
  assign n30316 = n30335 & n30336;
  assign n30252 = n30337 ^ n30338;
  assign n30304 = ~n30348;
  assign n26977 = n30357 ^ n30358;
  assign n30356 = n30376 & n30377;
  assign n30383 = n30397 & n30398;
  assign n30028 = ~n30081;
  assign n30082 = n30088 & n30089;
  assign n30058 = n30090 ^ n30091;
  assign n30092 = ~n30090;
  assign n30093 = ~n30116;
  assign n26497 = n30135 ^ n30136;
  assign n30163 = n30171 & n30172;
  assign n30227 = n30247 ^ n30248;
  assign n30249 = ~n30248;
  assign n30299 = n30252 & n349;
  assign n30296 = ~n30316;
  assign n30298 = ~n30252;
  assign n30180 = n30317 ^ n26977;
  assign n30319 = n26977 & n29575;
  assign n27029 = ~n26977;
  assign n30339 = ~n30356;
  assign n30359 = ~n30383;
  assign n30001 = n30058 ^ n30059;
  assign n30055 = ~n30082;
  assign n30083 = n30092 & n30093;
  assign n28890 = n27697 ^ n26497;
  assign n30098 = n26497 & n30114;
  assign n26516 = ~n26497;
  assign n30137 = ~n30163;
  assign n30209 = n30227 & n27623;
  assign n30067 = ~n30227;
  assign n30173 = n30249 & n30250;
  assign n30251 = n30296 & n30297;
  assign n30276 = n30298 & n12444;
  assign n30212 = ~n30299;
  assign n30277 = n30180 & n30300;
  assign n30278 = ~n30180;
  assign n30309 = n27029 & n30318;
  assign n29578 = ~n30319;
  assign n30301 = n30339 & n30340;
  assign n30320 = n30359 & n30360;
  assign n30030 = n30001 & n425;
  assign n30029 = ~n30001;
  assign n30022 = n30055 ^ n30056;
  assign n30054 = n30057 & n30055;
  assign n30005 = n28890 ^ n28875;
  assign n30060 = ~n30083;
  assign n28923 = ~n30098;
  assign n30085 = n26516 & n28921;
  assign n30100 = n30137 & n30138;
  assign n30198 = n30067 & n27686;
  assign n30102 = ~n30209;
  assign n30210 = n30251 ^ n30252;
  assign n30253 = ~n30251;
  assign n30254 = ~n30276;
  assign n30182 = ~n30277;
  assign n30267 = n30278 & n30217;
  assign n30255 = n30301 ^ n30302;
  assign n29596 = ~n30309;
  assign n30303 = ~n30301;
  assign n30281 = n30320 ^ n28239;
  assign n30321 = ~n30320;
  assign n29997 = n426 ^ n30022;
  assign n30023 = n30029 & n6844;
  assign n29974 = ~n30030;
  assign n30027 = ~n30054;
  assign n30038 = n30005 & n30032;
  assign n30031 = n30060 & n30061;
  assign n30039 = ~n30005;
  assign n28944 = ~n30085;
  assign n30068 = n30100 ^ n27623;
  assign n30101 = ~n30100;
  assign n30070 = ~n30198;
  assign n30174 = n349 ^ n30210;
  assign n30237 = n30253 & n30254;
  assign n30176 = n30255 ^ n30256;
  assign n30219 = ~n30267;
  assign n26975 = n30280 ^ n30281;
  assign n30279 = n30303 & n30304;
  assign n30310 = n30321 & n30322;
  assign n28860 = n29996 ^ n29997;
  assign n29947 = n29997 & n29996;
  assign n30002 = ~n30023;
  assign n30000 = n30027 & n30028;
  assign n30004 = n30031 ^ n30032;
  assign n29981 = ~n30038;
  assign n30033 = n30039 & n30040;
  assign n30010 = ~n30031;
  assign n26412 = n30067 ^ n30068;
  assign n30094 = n30101 & n30102;
  assign n30154 = n30173 ^ n30174;
  assign n30103 = n30174 & n30173;
  assign n30214 = n30176 & n348;
  assign n30211 = ~n30237;
  assign n30213 = ~n30176;
  assign n30110 = n30238 ^ n26975;
  assign n30239 = n26975 & n30259;
  assign n26908 = ~n26975;
  assign n30257 = ~n30279;
  assign n30282 = ~n30310;
  assign n29969 = ~n28860;
  assign n29972 = n30000 ^ n30001;
  assign n29950 = n30004 ^ n30005;
  assign n30003 = ~n30000;
  assign n30009 = ~n30033;
  assign n30026 = n26412 & n30037;
  assign n28877 = n27686 ^ n26412;
  assign n26468 = ~n26412;
  assign n30069 = ~n30094;
  assign n30139 = n30154 & n27586;
  assign n30011 = ~n30154;
  assign n30175 = n30211 & n30212;
  assign n30199 = n30213 & n12352;
  assign n30142 = ~n30214;
  assign n30200 = n30110 & n30215;
  assign n30201 = ~n30110;
  assign n29539 = ~n30239;
  assign n30228 = n26908 & n29537;
  assign n30216 = n30257 & n30258;
  assign n30240 = n30282 & n30283;
  assign n29948 = n425 ^ n29972;
  assign n29975 = n29950 & n6815;
  assign n29976 = ~n29950;
  assign n29998 = n30002 & n30003;
  assign n30006 = n30009 & n30010;
  assign n29957 = n28877 ^ n28858;
  assign n28881 = ~n30026;
  assign n30025 = n26468 & n30036;
  assign n30041 = n30069 & n30070;
  assign n30127 = n30011 & n27668;
  assign n30043 = ~n30139;
  assign n30140 = n30175 ^ n30176;
  assign n30177 = ~n30175;
  assign n30178 = ~n30199;
  assign n30112 = ~n30200;
  assign n30188 = n30201 & n30146;
  assign n30179 = n30216 ^ n30217;
  assign n29561 = ~n30228;
  assign n30218 = ~n30216;
  assign n30203 = n30240 ^ n28179;
  assign n30241 = n30240 & n30260;
  assign n28801 = n29947 ^ n29948;
  assign n29905 = n29948 & n29947;
  assign n29952 = ~n29975;
  assign n29971 = n29976 & n424;
  assign n29973 = ~n29998;
  assign n29984 = n29957 & n29934;
  assign n29980 = ~n30006;
  assign n29982 = ~n29957;
  assign n28906 = ~n30025;
  assign n30012 = n30041 ^ n27668;
  assign n30042 = ~n30041;
  assign n30014 = ~n30127;
  assign n30104 = n348 ^ n30140;
  assign n30164 = n30177 & n30178;
  assign n30106 = n30179 ^ n30180;
  assign n30148 = ~n30188;
  assign n26842 = n30203 ^ n30204;
  assign n30202 = n30218 & n30219;
  assign n30220 = ~n30241;
  assign n29928 = ~n28801;
  assign n29912 = ~n29905;
  assign n29931 = ~n29971;
  assign n29949 = n29973 & n29974;
  assign n29956 = n29980 & n29981;
  assign n29977 = n29982 & n29983;
  assign n29959 = ~n29984;
  assign n29999 = n28906 & n28881;
  assign n26360 = n30011 ^ n30012;
  assign n30034 = n30042 & n30043;
  assign n30084 = n30103 ^ n30104;
  assign n30044 = n30104 & n30103;
  assign n30144 = n30106 & n347;
  assign n30141 = ~n30164;
  assign n30143 = ~n30106;
  assign n30165 = n26842 & n29520;
  assign n26906 = ~n26842;
  assign n30181 = ~n30202;
  assign n30183 = n30220 & n30221;
  assign n29929 = n29949 ^ n29950;
  assign n29933 = n29956 ^ n29957;
  assign n29951 = ~n29949;
  assign n29970 = n26360 & n28860;
  assign n29958 = ~n29956;
  assign n29936 = ~n29977;
  assign n28822 = n26360 ^ n27668;
  assign n28904 = ~n29999;
  assign n26404 = ~n26360;
  assign n30013 = ~n30034;
  assign n30071 = n30084 & n27595;
  assign n29961 = ~n30084;
  assign n30105 = n30141 & n30142;
  assign n30128 = n30143 & n12313;
  assign n30074 = ~n30144;
  assign n30051 = n30155 ^ n26906;
  assign n29512 = ~n30165;
  assign n30156 = n26906 & n30166;
  assign n30145 = n30181 & n30182;
  assign n29474 = n30183 ^ n30184;
  assign n29906 = n424 ^ n29929;
  assign n29889 = n29933 ^ n29934;
  assign n29946 = n29951 & n29952;
  assign n29953 = n29958 & n29959;
  assign n29904 = n28822 ^ n28750;
  assign n29955 = n26404 & n29969;
  assign n28862 = ~n29970;
  assign n29985 = n30013 & n30014;
  assign n30062 = n29961 & n27547;
  assign n29987 = ~n30071;
  assign n30072 = n30105 ^ n30106;
  assign n30107 = ~n30105;
  assign n30108 = ~n30128;
  assign n30117 = n30051 & n30129;
  assign n30109 = n30145 ^ n30146;
  assign n30118 = ~n30051;
  assign n29995 = n29474 ^ n30149;
  assign n29533 = ~n30156;
  assign n30147 = ~n30145;
  assign n26825 = ~n29474;
  assign n28763 = n29905 ^ n29906;
  assign n29871 = n29906 & n29912;
  assign n29913 = n29889 & n6709;
  assign n29914 = ~n29889;
  assign n29930 = ~n29946;
  assign n29935 = ~n29953;
  assign n28839 = ~n29955;
  assign n29960 = n29985 ^ n27595;
  assign n29986 = ~n29985;
  assign n29963 = ~n30062;
  assign n30045 = n347 ^ n30072;
  assign n30095 = n30107 & n30108;
  assign n30047 = n30109 ^ n30110;
  assign n30053 = ~n30117;
  assign n30113 = n30118 & n30078;
  assign n30096 = n30131 ^ n26825;
  assign n30130 = n30147 & n30148;
  assign n29887 = ~n28763;
  assign n29874 = ~n29871;
  assign n29901 = ~n29913;
  assign n29908 = n29914 & n439;
  assign n29907 = n29930 & n29931;
  assign n29925 = n29935 & n29936;
  assign n26344 = n29960 ^ n29961;
  assign n29978 = n29986 & n29987;
  assign n30024 = n30044 ^ n30045;
  assign n29988 = n30045 & n30044;
  assign n30076 = n30047 & n346;
  assign n30073 = ~n30095;
  assign n30075 = ~n30047;
  assign n29498 = n30096 ^ n30097;
  assign n30080 = ~n30113;
  assign n30111 = ~n30130;
  assign n29888 = n439 ^ n29907;
  assign n29883 = ~n29908;
  assign n29902 = ~n29907;
  assign n29915 = n29925 & n29926;
  assign n29924 = n26344 & n29928;
  assign n29909 = ~n29925;
  assign n28781 = n26344 ^ n27547;
  assign n26294 = ~n26344;
  assign n29962 = ~n29978;
  assign n30015 = n30024 & n27529;
  assign n29917 = ~n30024;
  assign n30046 = n30073 & n30074;
  assign n30063 = n30075 & n12199;
  assign n30018 = ~n30076;
  assign n30077 = n30111 & n30112;
  assign n29872 = n29888 ^ n29889;
  assign n29894 = n29901 & n29902;
  assign n29890 = n29909 ^ n29904;
  assign n29910 = n29909 & n29891;
  assign n29903 = ~n29915;
  assign n29854 = n28781 ^ n28711;
  assign n28804 = ~n29924;
  assign n29927 = n26294 & n28801;
  assign n29937 = n29962 & n29963;
  assign n30007 = n29917 & n27565;
  assign n29939 = ~n30015;
  assign n30016 = n30046 ^ n30047;
  assign n30048 = ~n30046;
  assign n30049 = ~n30063;
  assign n30050 = n30077 ^ n30078;
  assign n30079 = ~n30077;
  assign n29857 = n29871 ^ n29872;
  assign n29873 = ~n29872;
  assign n29852 = n29890 ^ n29891;
  assign n29882 = ~n29894;
  assign n29895 = n29903 & n29904;
  assign n29885 = ~n29910;
  assign n28827 = ~n29927;
  assign n29916 = n29937 ^ n27529;
  assign n29938 = ~n29937;
  assign n29919 = ~n30007;
  assign n29989 = n346 ^ n30016;
  assign n30035 = n30048 & n30049;
  assign n29991 = n30050 ^ n30051;
  assign n30064 = n30079 & n30080;
  assign n28725 = ~n29857;
  assign n29833 = n29873 & n29874;
  assign n29867 = n29882 & n29883;
  assign n29884 = ~n29895;
  assign n26239 = n29916 ^ n29917;
  assign n29932 = n29938 & n29939;
  assign n29877 = n29988 ^ n29989;
  assign n29940 = n29989 & n29988;
  assign n30020 = n29991 & n345;
  assign n30017 = ~n30035;
  assign n30019 = ~n29991;
  assign n30052 = ~n30064;
  assign n29847 = n29867 ^ n29852;
  assign n29869 = n29867 & n6678;
  assign n29868 = ~n29867;
  assign n29875 = n29884 & n29885;
  assign n29881 = n26239 & n29887;
  assign n28743 = n27565 ^ n26239;
  assign n26278 = ~n26239;
  assign n29918 = ~n29932;
  assign n29964 = n29877 & n27484;
  assign n29965 = ~n29877;
  assign n29943 = ~n29940;
  assign n29990 = n30017 & n30018;
  assign n30008 = n30019 & n12147;
  assign n29968 = ~n30020;
  assign n30021 = n30052 & n30053;
  assign n29834 = n438 ^ n29847;
  assign n29858 = n29868 & n438;
  assign n29851 = ~n29869;
  assign n29870 = n29875 & n29876;
  assign n29859 = ~n29875;
  assign n29805 = n28743 ^ n28722;
  assign n28765 = ~n29881;
  assign n29886 = n26278 & n28763;
  assign n29896 = n29918 & n29919;
  assign n29898 = ~n29964;
  assign n29954 = n29965 & n27527;
  assign n29966 = n29990 ^ n29991;
  assign n29992 = ~n29990;
  assign n29993 = ~n30008;
  assign n29994 = n344 ^ n30021;
  assign n28682 = n29833 ^ n29834;
  assign n29782 = n29834 & n29833;
  assign n29848 = n29851 & n29852;
  assign n29837 = ~n29858;
  assign n29840 = n29859 ^ n29854;
  assign n29860 = n29859 & n29841;
  assign n29853 = ~n29870;
  assign n29863 = n29805 & n29823;
  assign n29861 = ~n29805;
  assign n28786 = ~n29886;
  assign n29878 = n29896 ^ n27527;
  assign n29897 = ~n29896;
  assign n29880 = ~n29954;
  assign n29941 = n345 ^ n29966;
  assign n29979 = n29992 & n29993;
  assign n29945 = n29994 ^ n29995;
  assign n29815 = ~n28682;
  assign n29785 = ~n29782;
  assign n29810 = n29840 ^ n29841;
  assign n29836 = ~n29848;
  assign n29849 = n29853 & n29854;
  assign n29839 = ~n29860;
  assign n29855 = n29861 & n29862;
  assign n29807 = ~n29863;
  assign n26227 = n29877 ^ n29878;
  assign n29892 = n29897 & n29898;
  assign n29842 = n29940 ^ n29941;
  assign n29942 = ~n29941;
  assign n29967 = ~n29979;
  assign n29819 = n29836 & n29837;
  assign n29838 = ~n29849;
  assign n29846 = n26227 & n28725;
  assign n29825 = ~n29855;
  assign n28704 = n26227 ^ n27527;
  assign n26171 = ~n26227;
  assign n29879 = ~n29892;
  assign n29921 = n29842 & n27438;
  assign n29920 = ~n29842;
  assign n29922 = n29942 & n29943;
  assign n29944 = n29967 & n29968;
  assign n29802 = n29819 ^ n29810;
  assign n29821 = n29819 & n6625;
  assign n29820 = ~n29819;
  assign n29822 = n29838 & n29839;
  assign n29769 = n28704 ^ n28688;
  assign n28727 = ~n29846;
  assign n29850 = n26171 & n29857;
  assign n29864 = n29879 & n29880;
  assign n29911 = n29920 & n27473;
  assign n29845 = ~n29921;
  assign n29923 = n29944 ^ n29945;
  assign n29783 = n437 ^ n29802;
  assign n29817 = n29820 & n437;
  assign n29809 = ~n29821;
  assign n29804 = n29822 ^ n29823;
  assign n29824 = ~n29822;
  assign n29828 = n29769 & n29835;
  assign n29829 = ~n29769;
  assign n28748 = ~n29850;
  assign n29843 = n29864 ^ n27473;
  assign n29865 = ~n29864;
  assign n29866 = ~n29911;
  assign n29812 = n29922 ^ n29923;
  assign n28644 = n29782 ^ n29783;
  assign n29784 = ~n29783;
  assign n29773 = n29804 ^ n29805;
  assign n29803 = n29809 & n29810;
  assign n29795 = ~n29817;
  assign n29818 = n29824 & n29825;
  assign n29771 = ~n29828;
  assign n29826 = n29829 & n29789;
  assign n26099 = n29842 ^ n29843;
  assign n29856 = n29865 & n29866;
  assign n29899 = n29812 & n27384;
  assign n29900 = ~n29812;
  assign n29765 = ~n28644;
  assign n29735 = n29784 & n29785;
  assign n29786 = n29773 & n6577;
  assign n29787 = ~n29773;
  assign n29794 = ~n29803;
  assign n29808 = n26099 & n29815;
  assign n29806 = ~n29818;
  assign n29791 = ~n29826;
  assign n28663 = n27438 ^ n26099;
  assign n26120 = ~n26099;
  assign n29844 = ~n29856;
  assign n29814 = ~n29899;
  assign n29893 = n29900 & n27426;
  assign n29738 = ~n29735;
  assign n29775 = ~n29786;
  assign n29780 = n29787 & n436;
  assign n29772 = n29794 & n29795;
  assign n29788 = n29806 & n29807;
  assign n28685 = ~n29808;
  assign n29732 = n28663 ^ n28613;
  assign n29816 = n26120 & n28682;
  assign n29830 = n29844 & n29845;
  assign n29832 = ~n29893;
  assign n29755 = n29772 ^ n29773;
  assign n29757 = ~n29780;
  assign n29774 = ~n29772;
  assign n29768 = n29788 ^ n29789;
  assign n29790 = ~n29788;
  assign n29796 = n29732 & n29750;
  assign n29797 = ~n29732;
  assign n28709 = ~n29816;
  assign n29811 = n29830 ^ n27426;
  assign n29831 = ~n29830;
  assign n29736 = n436 ^ n29755;
  assign n29740 = n29768 ^ n29769;
  assign n29767 = n29774 & n29775;
  assign n29781 = n29790 & n29791;
  assign n29752 = ~n29796;
  assign n29792 = n29797 & n29798;
  assign n26064 = n29811 ^ n29812;
  assign n29827 = n29831 & n29832;
  assign n28606 = n29735 ^ n29736;
  assign n29737 = ~n29736;
  assign n29748 = n29740 & n435;
  assign n29747 = ~n29740;
  assign n29756 = ~n29767;
  assign n29766 = n26064 & n28644;
  assign n29770 = ~n29781;
  assign n29734 = ~n29792;
  assign n28625 = n26064 ^ n27384;
  assign n26016 = ~n26064;
  assign n29813 = ~n29827;
  assign n29719 = ~n28606;
  assign n29701 = n29737 & n29738;
  assign n29745 = n29747 & n6508;
  assign n29709 = ~n29748;
  assign n29739 = n29756 & n29757;
  assign n29764 = n26016 & n29765;
  assign n28646 = ~n29766;
  assign n29749 = n29770 & n29771;
  assign n29698 = n28625 ^ n28611;
  assign n29799 = n29813 & n29814;
  assign n29720 = n29739 ^ n29740;
  assign n29729 = ~n29745;
  assign n29730 = ~n29739;
  assign n29731 = n29749 ^ n29750;
  assign n28667 = ~n29764;
  assign n29751 = ~n29749;
  assign n29758 = n29698 & n29713;
  assign n29759 = ~n29698;
  assign n29776 = n29799 ^ n27320;
  assign n29800 = ~n29799;
  assign n29702 = n435 ^ n29720;
  assign n29728 = n29729 & n29730;
  assign n29694 = n29731 ^ n29732;
  assign n29746 = n29751 & n29752;
  assign n29700 = ~n29758;
  assign n29753 = n29759 & n29760;
  assign n25941 = n29776 ^ n29777;
  assign n29793 = n29800 & n29801;
  assign n29690 = n29701 ^ n29702;
  assign n29651 = n29702 & n29701;
  assign n29707 = n29719 & n25941;
  assign n29710 = n29694 & n6432;
  assign n29708 = ~n29728;
  assign n29711 = ~n29694;
  assign n29733 = ~n29746;
  assign n29715 = ~n29753;
  assign n28586 = n27382 ^ n25941;
  assign n25989 = ~n25941;
  assign n29778 = ~n29793;
  assign n29679 = ~n29690;
  assign n29661 = ~n29651;
  assign n28608 = ~n29707;
  assign n29693 = n29708 & n29709;
  assign n29696 = ~n29710;
  assign n29705 = n29711 & n434;
  assign n29718 = n25989 & n28606;
  assign n29712 = n29733 & n29734;
  assign n29657 = n28586 ^ n28564;
  assign n29761 = n29778 & n29779;
  assign n29667 = n29693 ^ n29694;
  assign n29695 = ~n29693;
  assign n29669 = ~n29705;
  assign n29697 = n29712 ^ n29713;
  assign n28630 = ~n29718;
  assign n29714 = ~n29712;
  assign n29723 = n29657 & n29673;
  assign n29721 = ~n29657;
  assign n29741 = n29761 ^ n27355;
  assign n29762 = ~n29761;
  assign n29652 = n434 ^ n29667;
  assign n29691 = n29695 & n29696;
  assign n29654 = n29697 ^ n29698;
  assign n29706 = n29714 & n29715;
  assign n29716 = n29721 & n29722;
  assign n29660 = ~n29723;
  assign n25828 = n29741 ^ n29742;
  assign n29754 = n29762 & n29763;
  assign n28548 = n29651 ^ n29652;
  assign n29613 = n29652 & n29661;
  assign n29666 = n25828 & n29679;
  assign n29670 = n29654 & n6316;
  assign n29668 = ~n29691;
  assign n29671 = ~n29654;
  assign n29699 = ~n29706;
  assign n29675 = ~n29716;
  assign n28556 = n25828 ^ n27215;
  assign n25929 = ~n25828;
  assign n29743 = ~n29754;
  assign n29630 = ~n28548;
  assign n28569 = ~n29666;
  assign n29653 = n29668 & n29669;
  assign n29656 = ~n29670;
  assign n29664 = n29671 & n433;
  assign n29680 = n25929 & n29690;
  assign n29672 = n29699 & n29700;
  assign n29638 = n28556 ^ n28546;
  assign n29724 = n29743 & n29744;
  assign n29632 = n29653 ^ n29654;
  assign n29655 = ~n29653;
  assign n29634 = ~n29664;
  assign n29658 = n29672 ^ n29673;
  assign n28591 = ~n29680;
  assign n29674 = ~n29672;
  assign n29681 = n29638 & n29692;
  assign n29682 = ~n29638;
  assign n28508 = n29724 ^ n29725;
  assign n29726 = ~n29724;
  assign n29614 = n433 ^ n29632;
  assign n29648 = n29655 & n29656;
  assign n29616 = n29657 ^ n29658;
  assign n29650 = n28591 & n28569;
  assign n29665 = n29674 & n29675;
  assign n29640 = ~n29681;
  assign n29676 = n29682 & n29620;
  assign n29605 = n28508 ^ n28487;
  assign n25833 = n28508 ^ n27150;
  assign n29717 = n29726 & n29727;
  assign n28490 = n29613 ^ n29614;
  assign n29579 = n29614 & n29613;
  assign n29626 = n25833 & n29630;
  assign n29635 = n29616 & n6292;
  assign n29633 = ~n29648;
  assign n29636 = ~n29616;
  assign n28589 = ~n29650;
  assign n29659 = ~n29665;
  assign n29622 = ~n29676;
  assign n29683 = n29605 & n29587;
  assign n29684 = ~n29605;
  assign n25755 = ~n25833;
  assign n29703 = ~n29717;
  assign n29598 = ~n28490;
  assign n29582 = ~n29579;
  assign n28526 = ~n29626;
  assign n29615 = n29633 & n29634;
  assign n29618 = ~n29635;
  assign n29627 = n29636 & n432;
  assign n29631 = n25755 & n28548;
  assign n29637 = n29659 & n29660;
  assign n29607 = ~n29683;
  assign n29677 = n29684 & n29685;
  assign n29686 = n29703 & n29704;
  assign n29599 = n29615 ^ n29616;
  assign n29617 = ~n29615;
  assign n29601 = ~n29627;
  assign n28550 = ~n29631;
  assign n29619 = n29637 ^ n29638;
  assign n29639 = ~n29637;
  assign n29589 = ~n29677;
  assign n28469 = n29686 ^ n29687;
  assign n29688 = ~n29686;
  assign n29580 = n432 ^ n29599;
  assign n29610 = n29617 & n29618;
  assign n29565 = n29619 ^ n29620;
  assign n29628 = n29639 & n29640;
  assign n29571 = n28469 ^ n28450;
  assign n25675 = n28469 ^ n27079;
  assign n29678 = n29688 & n29689;
  assign n28443 = n29579 ^ n29580;
  assign n29581 = ~n29580;
  assign n29591 = n25675 & n29598;
  assign n29603 = n29565 & n447;
  assign n29600 = ~n29610;
  assign n29602 = ~n29565;
  assign n29621 = ~n29628;
  assign n29643 = n29571 & n29549;
  assign n29644 = ~n29571;
  assign n25769 = ~n25675;
  assign n29662 = ~n29678;
  assign n29563 = ~n28443;
  assign n29540 = n29581 & n29582;
  assign n28512 = ~n29591;
  assign n29583 = n29600 & n29601;
  assign n29592 = n29602 & n6169;
  assign n29567 = ~n29603;
  assign n29597 = n25769 & n28490;
  assign n29604 = n29621 & n29622;
  assign n29573 = ~n29643;
  assign n29641 = n29644 & n29645;
  assign n29649 = n29662 & n29663;
  assign n29543 = ~n29540;
  assign n29564 = n447 ^ n29583;
  assign n29584 = ~n29583;
  assign n29585 = ~n29592;
  assign n28492 = ~n29597;
  assign n29586 = n29604 ^ n29605;
  assign n29606 = ~n29604;
  assign n29551 = ~n29641;
  assign n29647 = n29649 & n27047;
  assign n29646 = ~n29649;
  assign n29541 = n29564 ^ n29565;
  assign n29574 = n29584 & n29585;
  assign n29545 = n29586 ^ n29587;
  assign n29593 = n29606 & n29607;
  assign n29642 = n29646 & n27119;
  assign n29625 = ~n29647;
  assign n28400 = n29540 ^ n29541;
  assign n29542 = ~n29541;
  assign n29568 = n29545 & n6144;
  assign n29566 = ~n29574;
  assign n29569 = ~n29545;
  assign n29588 = ~n29593;
  assign n29624 = n29625 & n29629;
  assign n29612 = ~n29642;
  assign n29522 = ~n28400;
  assign n29500 = n29542 & n29543;
  assign n29544 = n29566 & n29567;
  assign n29547 = ~n29568;
  assign n29557 = n29569 & n446;
  assign n29570 = n29588 & n29589;
  assign n29611 = ~n29624;
  assign n29623 = n29612 & n29625;
  assign n29524 = n29544 ^ n29545;
  assign n29546 = ~n29544;
  assign n29526 = ~n29557;
  assign n29548 = n29570 ^ n29571;
  assign n29572 = ~n29570;
  assign n29594 = n29611 & n29612;
  assign n29608 = ~n29623;
  assign n29501 = n446 ^ n29524;
  assign n29534 = n29546 & n29547;
  assign n29503 = n29548 ^ n29549;
  assign n29558 = n29572 & n29573;
  assign n29576 = n29594 ^ n26977;
  assign n25692 = n29608 ^ n29609;
  assign n29595 = ~n29594;
  assign n28347 = n29500 ^ n29501;
  assign n29464 = n29501 & n29500;
  assign n29527 = n29503 & n6018;
  assign n29525 = ~n29534;
  assign n29528 = ~n29503;
  assign n29550 = ~n29558;
  assign n29556 = n25692 & n29563;
  assign n25564 = n29575 ^ n29576;
  assign n28412 = n27119 ^ n25692;
  assign n29590 = n29595 & n29596;
  assign n25638 = ~n25692;
  assign n29486 = ~n28347;
  assign n29515 = n25564 & n29522;
  assign n29502 = n29525 & n29526;
  assign n29505 = ~n29527;
  assign n29516 = n29528 & n445;
  assign n29529 = n29550 & n29551;
  assign n28446 = ~n29556;
  assign n29506 = n28412 ^ n28355;
  assign n29562 = n25638 & n28443;
  assign n25617 = ~n25564;
  assign n29577 = ~n29590;
  assign n29487 = n29502 ^ n29503;
  assign n28426 = ~n29515;
  assign n29504 = ~n29502;
  assign n29489 = ~n29516;
  assign n29507 = n29529 ^ n29530;
  assign n29523 = n25617 & n28400;
  assign n29531 = ~n29529;
  assign n29552 = n29506 & n29530;
  assign n28373 = n25617 ^ n26977;
  assign n29553 = ~n29506;
  assign n28474 = ~n29562;
  assign n29559 = n29577 & n29578;
  assign n29465 = n445 ^ n29487;
  assign n29499 = n29504 & n29505;
  assign n29467 = n29506 ^ n29507;
  assign n28403 = ~n29523;
  assign n29471 = n28353 ^ n28373;
  assign n29532 = ~n29552;
  assign n29535 = n29553 & n29554;
  assign n29536 = n29559 ^ n26908;
  assign n29560 = ~n29559;
  assign n28291 = n29464 ^ n29465;
  assign n29434 = n29465 & n29464;
  assign n29490 = n29467 & n5930;
  assign n29488 = ~n29499;
  assign n29491 = ~n29467;
  assign n29513 = n29471 & n29518;
  assign n29517 = n29531 & n29532;
  assign n29514 = ~n29471;
  assign n29509 = ~n29535;
  assign n25541 = n29536 ^ n29537;
  assign n29555 = n29560 & n29561;
  assign n29451 = ~n28291;
  assign n29437 = ~n29434;
  assign n29477 = n25541 & n29486;
  assign n29466 = n29488 & n29489;
  assign n29469 = ~n29490;
  assign n29478 = n29491 & n444;
  assign n29473 = ~n29513;
  assign n29510 = n29514 & n29493;
  assign n29508 = ~n29517;
  assign n28320 = n26975 ^ n25541;
  assign n25490 = ~n25541;
  assign n29538 = ~n29555;
  assign n29452 = n29466 ^ n29467;
  assign n28377 = ~n29477;
  assign n29468 = ~n29466;
  assign n29454 = ~n29478;
  assign n29485 = n25490 & n28347;
  assign n29443 = n28320 ^ n28239;
  assign n29492 = n29508 & n29509;
  assign n29495 = ~n29510;
  assign n29519 = n29538 & n29539;
  assign n29435 = n444 ^ n29452;
  assign n29463 = n29468 & n29469;
  assign n28350 = ~n29485;
  assign n29470 = n29492 ^ n29493;
  assign n29480 = n29443 & n29458;
  assign n29481 = ~n29443;
  assign n29494 = ~n29492;
  assign n28265 = n29519 ^ n29520;
  assign n29521 = n29519 & n29533;
  assign n28233 = n29434 ^ n29435;
  assign n29436 = ~n29435;
  assign n29453 = ~n29463;
  assign n29439 = n29470 ^ n29471;
  assign n29445 = ~n29480;
  assign n29475 = n29481 & n29482;
  assign n29479 = n29494 & n29495;
  assign n29419 = n28265 ^ n28230;
  assign n25420 = n28265 ^ n26842;
  assign n29511 = ~n29521;
  assign n29410 = n29436 & n29437;
  assign n29447 = n25420 & n29451;
  assign n29438 = n29453 & n29454;
  assign n29456 = n29439 & n443;
  assign n29455 = ~n29439;
  assign n29460 = ~n29475;
  assign n29472 = ~n29479;
  assign n29484 = n29419 & n29496;
  assign n29483 = ~n29419;
  assign n25465 = ~n25420;
  assign n29497 = n29511 & n29512;
  assign n29413 = ~n29410;
  assign n29424 = n29438 ^ n29439;
  assign n28325 = ~n29447;
  assign n29440 = ~n29438;
  assign n29448 = n29455 & n5860;
  assign n29426 = ~n29456;
  assign n29450 = n25465 & n28291;
  assign n29457 = n29472 & n29473;
  assign n29476 = n29483 & n29430;
  assign n29421 = ~n29484;
  assign n26860 = n29497 ^ n29498;
  assign n29411 = n443 ^ n29424;
  assign n29441 = ~n29448;
  assign n28294 = ~n29450;
  assign n29442 = n29457 ^ n29458;
  assign n29459 = ~n29457;
  assign n29461 = n29474 ^ n26860;
  assign n29432 = ~n29476;
  assign n27511 = n29410 ^ n29411;
  assign n29412 = ~n29411;
  assign n29433 = n29440 & n29441;
  assign n29415 = n29442 ^ n29443;
  assign n29449 = n29459 & n29460;
  assign n28205 = n29461 ^ n29462;
  assign n29399 = n28460 ^ n27511;
  assign n29388 = n27511 ^ n29402;
  assign n26604 = n27490 ^ n27511;
  assign n29361 = n27511 & n27490;
  assign n29389 = n29412 & n29413;
  assign n29427 = n29415 & n5793;
  assign n29425 = ~n29433;
  assign n29428 = ~n29415;
  assign n29398 = n28205 ^ n29446;
  assign n29444 = ~n29449;
  assign n27903 = n7 ^ n29388;
  assign n29343 = n29399 & n29400;
  assign n29294 = n29388 & n7;
  assign n29392 = ~n29389;
  assign n29414 = n29425 & n29426;
  assign n29417 = ~n29427;
  assign n29422 = n29428 & n442;
  assign n29429 = n29444 & n29445;
  assign n29385 = n29343 & n29335;
  assign n29052 = ~n27903;
  assign n29383 = ~n29343;
  assign n29403 = n29414 ^ n29415;
  assign n29416 = ~n29414;
  assign n29405 = ~n29422;
  assign n29418 = n29429 ^ n29430;
  assign n29431 = ~n29429;
  assign n29377 = n29383 & n29384;
  assign n29342 = ~n29385;
  assign n29390 = n442 ^ n29403;
  assign n29409 = n29416 & n29417;
  assign n29394 = n29418 ^ n29419;
  assign n29423 = n29431 & n29432;
  assign n29348 = ~n29377;
  assign n29386 = n29389 ^ n29390;
  assign n29391 = ~n29390;
  assign n29407 = n29394 & n441;
  assign n29404 = ~n29409;
  assign n29406 = ~n29394;
  assign n29420 = ~n29423;
  assign n29378 = n29386 & n27416;
  assign n29379 = ~n29386;
  assign n29370 = n29391 & n29392;
  assign n29393 = n29404 & n29405;
  assign n29401 = n29406 & n5708;
  assign n29382 = ~n29407;
  assign n29408 = n29420 & n29421;
  assign n29369 = ~n29378;
  assign n29376 = n29379 & n27434;
  assign n29373 = ~n29370;
  assign n29380 = n29393 ^ n29394;
  assign n29395 = ~n29393;
  assign n29396 = ~n29401;
  assign n29397 = n440 ^ n29408;
  assign n29368 = n29369 & n29361;
  assign n29367 = ~n29376;
  assign n29371 = n441 ^ n29380;
  assign n29387 = n29395 & n29396;
  assign n29375 = n29397 ^ n29398;
  assign n29366 = ~n29368;
  assign n29360 = n29367 & n29369;
  assign n29349 = n29370 ^ n29371;
  assign n29372 = ~n29371;
  assign n29381 = ~n29387;
  assign n26483 = n29360 ^ n29361;
  assign n29358 = n29366 & n29367;
  assign n29363 = n29349 & n27325;
  assign n29362 = ~n29349;
  assign n29364 = n29372 & n29373;
  assign n29374 = n29381 & n29382;
  assign n29344 = n26483 ^ n29353;
  assign n29350 = n29358 ^ n27333;
  assign n26470 = ~n26483;
  assign n29354 = ~n29358;
  assign n29359 = n29362 & n27333;
  assign n29347 = ~n29363;
  assign n29365 = n29374 ^ n29375;
  assign n29334 = n29343 ^ n29344;
  assign n29345 = n29344 & n29348;
  assign n26379 = n29349 ^ n29350;
  assign n29355 = ~n29359;
  assign n29325 = n29364 ^ n29365;
  assign n29329 = n29334 ^ n29335;
  assign n29312 = n29340 ^ n26379;
  assign n29341 = ~n29345;
  assign n26430 = ~n26379;
  assign n29351 = n29354 & n29355;
  assign n29356 = n29325 & n27221;
  assign n29357 = ~n29325;
  assign n29322 = n29329 & n6;
  assign n29331 = n29312 & n29332;
  assign n29321 = ~n29329;
  assign n29330 = ~n29312;
  assign n29336 = n29341 & n29342;
  assign n29346 = ~n29351;
  assign n29328 = ~n29356;
  assign n29352 = n29357 & n27246;
  assign n29320 = n29321 & n21721;
  assign n29296 = ~n29322;
  assign n29323 = n29330 & n29324;
  assign n29318 = ~n29331;
  assign n29319 = ~n29336;
  assign n29337 = n29346 & n29347;
  assign n29339 = ~n29352;
  assign n29317 = n29318 & n29319;
  assign n29310 = ~n29320;
  assign n29307 = ~n29323;
  assign n29311 = n29319 ^ n29324;
  assign n29326 = n29337 ^ n27246;
  assign n29338 = ~n29337;
  assign n29308 = n29310 & n29294;
  assign n29293 = n29310 & n29296;
  assign n29279 = n29311 ^ n29312;
  assign n29306 = ~n29317;
  assign n26336 = n29325 ^ n29326;
  assign n29333 = n29338 & n29339;
  assign n27847 = n29293 ^ n29294;
  assign n29297 = n29279 & n21670;
  assign n29289 = n29306 & n29307;
  assign n29295 = ~n29308;
  assign n29298 = ~n29279;
  assign n29275 = n29313 ^ n26336;
  assign n26330 = ~n26336;
  assign n29327 = ~n29333;
  assign n29274 = n29289 ^ n29290;
  assign n27870 = ~n27847;
  assign n29278 = n29295 & n29296;
  assign n29281 = ~n29297;
  assign n29291 = n29298 & n5;
  assign n29286 = ~n29289;
  assign n29301 = n29275 & n29290;
  assign n29299 = ~n29275;
  assign n29314 = n29327 & n29328;
  assign n29251 = n29274 ^ n29275;
  assign n29263 = n29278 ^ n29279;
  assign n29280 = ~n29278;
  assign n29265 = ~n29291;
  assign n29292 = n29299 & n29300;
  assign n29287 = ~n29301;
  assign n29303 = n29314 ^ n27146;
  assign n29315 = ~n29314;
  assign n29259 = n29251 & n21468;
  assign n29247 = n5 ^ n29263;
  assign n29260 = ~n29251;
  assign n29276 = n29280 & n29281;
  assign n29282 = n29286 & n29287;
  assign n29271 = ~n29292;
  assign n26235 = n29302 ^ n29303;
  assign n29309 = n29315 & n29316;
  assign n27819 = n29247 ^ n27847;
  assign n29216 = n29247 & n27847;
  assign n29248 = ~n29259;
  assign n29254 = n29260 & n4;
  assign n29264 = ~n29276;
  assign n29270 = ~n29282;
  assign n29239 = n29283 ^ n26235;
  assign n26232 = ~n26235;
  assign n29304 = ~n29309;
  assign n28978 = ~n27819;
  assign n29219 = ~n29216;
  assign n29234 = ~n29254;
  assign n29250 = n29264 & n29265;
  assign n29255 = n29270 & n29271;
  assign n29266 = n29239 & n29272;
  assign n29267 = ~n29239;
  assign n29288 = n29304 & n29305;
  assign n29232 = n29250 ^ n29251;
  assign n29238 = n29255 ^ n29256;
  assign n29249 = ~n29250;
  assign n29252 = ~n29255;
  assign n29236 = ~n29266;
  assign n29261 = n29267 & n29256;
  assign n29285 = n29288 & n27075;
  assign n29284 = ~n29288;
  assign n29217 = n4 ^ n29232;
  assign n29221 = n29238 ^ n29239;
  assign n29243 = n29248 & n29249;
  assign n29253 = ~n29261;
  assign n29277 = n29284 & n27115;
  assign n29269 = ~n29285;
  assign n28940 = n29216 ^ n29217;
  assign n29218 = ~n29217;
  assign n29226 = n29221 & n3;
  assign n29225 = ~n29221;
  assign n29233 = ~n29243;
  assign n29244 = n29252 & n29253;
  assign n29268 = n29269 & n29273;
  assign n29258 = ~n29277;
  assign n27786 = ~n28940;
  assign n29184 = n29218 & n29219;
  assign n29222 = n29225 & n21407;
  assign n29190 = ~n29226;
  assign n29220 = n29233 & n29234;
  assign n29235 = ~n29244;
  assign n29257 = ~n29268;
  assign n29262 = n29258 & n29269;
  assign n29201 = n29220 ^ n29221;
  assign n29206 = ~n29222;
  assign n29207 = ~n29220;
  assign n29223 = n29235 & n29236;
  assign n29240 = n29257 & n29258;
  assign n29245 = ~n29262;
  assign n29185 = n3 ^ n29201;
  assign n29202 = n29206 & n29207;
  assign n29203 = n29223 ^ n29215;
  assign n29200 = ~n29223;
  assign n29227 = n29240 ^ n27040;
  assign n26216 = n29245 ^ n29246;
  assign n29241 = ~n29240;
  assign n27752 = n29184 ^ n29185;
  assign n29145 = n29185 & n29184;
  assign n29189 = ~n29202;
  assign n26158 = n29227 ^ n29228;
  assign n29204 = n29231 ^ n26216;
  assign n29237 = n29241 & n29242;
  assign n26143 = ~n26216;
  assign n28901 = ~n27752;
  assign n29174 = n29189 & n29190;
  assign n29175 = n29203 ^ n29204;
  assign n29149 = n29208 ^ n26158;
  assign n29213 = n29204 & n29224;
  assign n26074 = ~n26158;
  assign n29214 = ~n29204;
  assign n29229 = ~n29237;
  assign n29158 = n29174 ^ n29175;
  assign n29172 = ~n29174;
  assign n29187 = n29175 & n2;
  assign n29186 = ~n29175;
  assign n29191 = n29149 & n29165;
  assign n29192 = ~n29149;
  assign n29183 = ~n29213;
  assign n29209 = n29214 & n29215;
  assign n29210 = n29229 & n29230;
  assign n29146 = n2 ^ n29158;
  assign n29181 = n29186 & n21353;
  assign n29156 = ~n29187;
  assign n29154 = ~n29191;
  assign n29188 = n29192 & n29193;
  assign n29199 = ~n29209;
  assign n29194 = n29210 ^ n26932;
  assign n29211 = ~n29210;
  assign n28878 = n29145 ^ n29146;
  assign n29094 = n29146 & n29145;
  assign n29171 = ~n29181;
  assign n29170 = ~n29188;
  assign n26056 = n29194 ^ n29195;
  assign n29196 = n29199 & n29200;
  assign n29205 = n29211 & n29212;
  assign n28888 = ~n28878;
  assign n29168 = n29171 & n29172;
  assign n29123 = n29176 ^ n26056;
  assign n25998 = ~n26056;
  assign n29182 = ~n29196;
  assign n29197 = ~n29205;
  assign n29155 = ~n29168;
  assign n29160 = n29123 & n29169;
  assign n29159 = ~n29123;
  assign n29177 = n29182 & n29183;
  assign n29178 = n29197 & n29198;
  assign n29128 = n29155 & n29156;
  assign n29157 = n29159 & n29141;
  assign n29125 = ~n29160;
  assign n29164 = ~n29177;
  assign n29162 = n29178 ^ n26832;
  assign n29179 = ~n29178;
  assign n29117 = ~n29128;
  assign n29143 = ~n29157;
  assign n26002 = n29162 ^ n29163;
  assign n29148 = n29164 ^ n29165;
  assign n29161 = n29170 & n29164;
  assign n29173 = n29179 & n29180;
  assign n29090 = n29147 ^ n26002;
  assign n29129 = n29148 ^ n29149;
  assign n25925 = ~n26002;
  assign n29153 = ~n29161;
  assign n29166 = ~n29173;
  assign n29115 = n29128 ^ n29129;
  assign n29132 = n29090 & n29139;
  assign n29133 = n29129 & n1;
  assign n29131 = ~n29090;
  assign n29130 = ~n29129;
  assign n29140 = n29153 & n29154;
  assign n29150 = n29166 & n29167;
  assign n29095 = n1 ^ n29115;
  assign n29126 = n29130 & n21237;
  assign n29127 = n29131 & n29110;
  assign n29092 = ~n29132;
  assign n29098 = ~n29133;
  assign n29122 = n29140 ^ n29141;
  assign n29142 = ~n29140;
  assign n29135 = n29150 ^ n26773;
  assign n29151 = ~n29150;
  assign n28824 = n29094 ^ n29095;
  assign n29044 = n29095 & n29094;
  assign n29084 = n29122 ^ n29123;
  assign n29116 = ~n29126;
  assign n29112 = ~n29127;
  assign n25855 = n29135 ^ n29136;
  assign n29134 = n29142 & n29143;
  assign n29144 = n29151 & n29152;
  assign n27706 = ~n28824;
  assign n29107 = n29084 & n0;
  assign n29106 = ~n29084;
  assign n29113 = n29116 & n29117;
  assign n29057 = n29118 ^ n25855;
  assign n25853 = ~n25855;
  assign n29124 = ~n29134;
  assign n29137 = ~n29144;
  assign n29096 = n29106 & n21168;
  assign n29063 = ~n29107;
  assign n29099 = n29057 & n29108;
  assign n29097 = ~n29113;
  assign n29100 = ~n29057;
  assign n29109 = n29124 & n29125;
  assign n29119 = n29137 & n29138;
  assign n29081 = ~n29096;
  assign n29083 = n29097 & n29098;
  assign n29059 = ~n29099;
  assign n29093 = n29100 & n29076;
  assign n29089 = n29109 ^ n29110;
  assign n29111 = ~n29109;
  assign n29103 = n29119 ^ n26722;
  assign n29120 = ~n29119;
  assign n29061 = n29083 ^ n29084;
  assign n29047 = n29089 ^ n29090;
  assign n29082 = ~n29083;
  assign n29078 = ~n29093;
  assign n25747 = n29102 ^ n29103;
  assign n29101 = n29111 & n29112;
  assign n29114 = n29120 & n29121;
  assign n29045 = n0 ^ n29061;
  assign n29073 = n29047 & n15;
  assign n29079 = n29081 & n29082;
  assign n29072 = ~n29047;
  assign n29019 = n29085 ^ n25747;
  assign n25745 = ~n25747;
  assign n29091 = ~n29101;
  assign n29104 = ~n29114;
  assign n28782 = n29044 ^ n29045;
  assign n29008 = n29045 & n29044;
  assign n29064 = n29072 & n21044;
  assign n29025 = ~n29073;
  assign n29065 = n29019 & n29074;
  assign n29062 = ~n29079;
  assign n29066 = ~n29019;
  assign n29075 = n29091 & n29092;
  assign n29086 = n29104 & n29105;
  assign n27650 = ~n28782;
  assign n29046 = n29062 & n29063;
  assign n29049 = ~n29064;
  assign n29021 = ~n29065;
  assign n29060 = n29066 & n29038;
  assign n29056 = n29075 ^ n29076;
  assign n29077 = ~n29075;
  assign n29069 = n29086 ^ n26706;
  assign n29087 = ~n29086;
  assign n29023 = n29046 ^ n29047;
  assign n29011 = n29056 ^ n29057;
  assign n29048 = ~n29046;
  assign n29040 = ~n29060;
  assign n25751 = n29068 ^ n29069;
  assign n29067 = n29077 & n29078;
  assign n29080 = n29087 & n29088;
  assign n29009 = n15 ^ n29023;
  assign n29035 = n29011 & n14;
  assign n29041 = n29048 & n29049;
  assign n29034 = ~n29011;
  assign n28984 = n29050 ^ n25751;
  assign n29051 = n25751 & n27903;
  assign n25645 = ~n25751;
  assign n29058 = ~n29067;
  assign n29070 = ~n29080;
  assign n27616 = n29008 ^ n29009;
  assign n28971 = n29009 & n29008;
  assign n29026 = n29034 & n20935;
  assign n28990 = ~n29035;
  assign n29027 = n28984 & n29036;
  assign n29024 = ~n29041;
  assign n29028 = ~n28984;
  assign n27905 = ~n29051;
  assign n29042 = n25645 & n29052;
  assign n29037 = n29058 & n29059;
  assign n29053 = n29070 & n29071;
  assign n28744 = ~n27616;
  assign n29010 = n29024 & n29025;
  assign n29013 = ~n29026;
  assign n28986 = ~n29027;
  assign n29022 = n29028 & n29003;
  assign n29018 = n29037 ^ n29038;
  assign n27923 = ~n29042;
  assign n29039 = ~n29037;
  assign n29031 = n29053 ^ n26635;
  assign n29054 = ~n29053;
  assign n28988 = n29010 ^ n29011;
  assign n28974 = n29018 ^ n29019;
  assign n29012 = ~n29010;
  assign n29005 = ~n29022;
  assign n25574 = n29030 ^ n29031;
  assign n29029 = n29039 & n29040;
  assign n29043 = n29054 & n29055;
  assign n28972 = n14 ^ n28988;
  assign n29001 = n28974 & n13;
  assign n29006 = n29012 & n29013;
  assign n29000 = ~n28974;
  assign n28946 = n29014 ^ n25574;
  assign n25669 = ~n25574;
  assign n29020 = ~n29029;
  assign n29032 = ~n29043;
  assign n28705 = n28971 ^ n28972;
  assign n28933 = n28972 & n28971;
  assign n28991 = n29000 & n20920;
  assign n28952 = ~n29001;
  assign n28992 = n28946 & n28965;
  assign n28989 = ~n29006;
  assign n28993 = ~n28946;
  assign n29002 = n29020 & n29021;
  assign n29015 = n29032 & n29033;
  assign n27575 = ~n28705;
  assign n28973 = n28989 & n28990;
  assign n28976 = ~n28991;
  assign n28967 = ~n28992;
  assign n28987 = n28993 & n28994;
  assign n28983 = n29002 ^ n29003;
  assign n29004 = ~n29002;
  assign n28996 = n29015 ^ n26592;
  assign n29016 = ~n29015;
  assign n28950 = n28973 ^ n28974;
  assign n28936 = n28983 ^ n28984;
  assign n28975 = ~n28973;
  assign n28948 = ~n28987;
  assign n25589 = n28996 ^ n28997;
  assign n28995 = n29004 & n29005;
  assign n29007 = n29016 & n29017;
  assign n28934 = n13 ^ n28950;
  assign n28963 = n28936 & n12;
  assign n28968 = n28975 & n28976;
  assign n28962 = ~n28936;
  assign n28908 = n25589 ^ n28977;
  assign n28979 = n25589 & n27819;
  assign n25497 = ~n25589;
  assign n28985 = ~n28995;
  assign n28998 = ~n29007;
  assign n27534 = n28933 ^ n28934;
  assign n28893 = n28934 & n28933;
  assign n28953 = n28962 & n20836;
  assign n28914 = ~n28963;
  assign n28954 = n28908 & n28927;
  assign n28951 = ~n28968;
  assign n28955 = ~n28908;
  assign n28969 = n25497 & n28978;
  assign n27821 = ~n28979;
  assign n28964 = n28985 & n28986;
  assign n28980 = n28998 & n28999;
  assign n28673 = ~n27534;
  assign n28896 = ~n28893;
  assign n28935 = n28951 & n28952;
  assign n28938 = ~n28953;
  assign n28910 = ~n28954;
  assign n28949 = n28955 & n28956;
  assign n28945 = n28964 ^ n28965;
  assign n27835 = ~n28969;
  assign n28966 = ~n28964;
  assign n28959 = n28980 ^ n26550;
  assign n28981 = ~n28980;
  assign n28912 = n28935 ^ n28936;
  assign n28898 = n28945 ^ n28946;
  assign n28937 = ~n28935;
  assign n28929 = ~n28949;
  assign n25502 = n28958 ^ n28959;
  assign n28957 = n28966 & n28967;
  assign n28970 = n28981 & n28982;
  assign n28894 = n12 ^ n28912;
  assign n28924 = n28898 & n20775;
  assign n28930 = n28937 & n28938;
  assign n28925 = ~n28898;
  assign n28864 = n28939 ^ n25502;
  assign n28941 = n25502 & n27786;
  assign n25427 = ~n25502;
  assign n28947 = ~n28957;
  assign n28960 = ~n28970;
  assign n27502 = n28893 ^ n28894;
  assign n28895 = ~n28894;
  assign n28900 = ~n28924;
  assign n28915 = n28925 & n11;
  assign n28918 = n28864 & n28885;
  assign n28913 = ~n28930;
  assign n28916 = ~n28864;
  assign n28931 = n25427 & n28940;
  assign n27789 = ~n28941;
  assign n28926 = n28947 & n28948;
  assign n28942 = n28960 & n28961;
  assign n28627 = ~n27502;
  assign n28850 = n28895 & n28896;
  assign n28897 = n28913 & n28914;
  assign n28873 = ~n28915;
  assign n28911 = n28916 & n28917;
  assign n28887 = ~n28918;
  assign n28907 = n28926 ^ n28927;
  assign n27804 = ~n28931;
  assign n28928 = ~n28926;
  assign n28920 = n28942 ^ n26516;
  assign n28943 = ~n28942;
  assign n28871 = n28897 ^ n28898;
  assign n28853 = n28907 ^ n28908;
  assign n28899 = ~n28897;
  assign n28866 = ~n28911;
  assign n25364 = n28920 ^ n28921;
  assign n28919 = n28928 & n28929;
  assign n28932 = n28943 & n28944;
  assign n28851 = n11 ^ n28871;
  assign n28882 = n28853 & n20683;
  assign n28889 = n28899 & n28900;
  assign n28883 = ~n28853;
  assign n28902 = n25364 & n27752;
  assign n25443 = ~n25364;
  assign n28909 = ~n28919;
  assign n28922 = ~n28932;
  assign n27453 = n28850 ^ n28851;
  assign n28814 = n28851 & n28850;
  assign n28854 = ~n28882;
  assign n28874 = n28883 & n10;
  assign n28872 = ~n28889;
  assign n28829 = n28890 ^ n25443;
  assign n28891 = n25443 & n28901;
  assign n27772 = ~n28902;
  assign n28884 = n28909 & n28910;
  assign n28903 = n28922 & n28923;
  assign n28596 = ~n27453;
  assign n28817 = ~n28814;
  assign n28852 = n28872 & n28873;
  assign n28834 = ~n28874;
  assign n28868 = n28829 & n28875;
  assign n28863 = n28884 ^ n28885;
  assign n28869 = ~n28829;
  assign n27755 = ~n28891;
  assign n28886 = ~n28884;
  assign n25286 = n28903 ^ n28904;
  assign n28905 = ~n28903;
  assign n28832 = n28852 ^ n28853;
  assign n28819 = n28863 ^ n28864;
  assign n28855 = ~n28852;
  assign n28831 = ~n28868;
  assign n28867 = n28869 & n28843;
  assign n28808 = n28877 ^ n25286;
  assign n28876 = n28886 & n28887;
  assign n28879 = n25286 & n28888;
  assign n25377 = ~n25286;
  assign n28892 = n28905 & n28906;
  assign n28815 = n10 ^ n28832;
  assign n28840 = n28819 & n20607;
  assign n28846 = n28854 & n28855;
  assign n28841 = ~n28819;
  assign n28856 = n28808 & n28789;
  assign n28845 = ~n28867;
  assign n28857 = ~n28808;
  assign n28865 = ~n28876;
  assign n28870 = n25377 & n28878;
  assign n27722 = ~n28879;
  assign n28880 = ~n28892;
  assign n28566 = n28814 ^ n28815;
  assign n28816 = ~n28815;
  assign n28821 = ~n28840;
  assign n28835 = n28841 & n9;
  assign n28833 = ~n28846;
  assign n28791 = ~n28856;
  assign n28847 = n28857 & n28858;
  assign n28842 = n28865 & n28866;
  assign n27740 = ~n28870;
  assign n28859 = n28880 & n28881;
  assign n28576 = ~n28566;
  assign n28775 = n28816 & n28817;
  assign n28818 = n28833 & n28834;
  assign n28795 = ~n28835;
  assign n28828 = n28842 ^ n28843;
  assign n28810 = ~n28847;
  assign n28844 = ~n28842;
  assign n28848 = n27740 & n27722;
  assign n28837 = n28859 ^ n28860;
  assign n28861 = ~n28859;
  assign n28787 = ~n28775;
  assign n28793 = n28818 ^ n28819;
  assign n28778 = n28828 ^ n28829;
  assign n28820 = ~n28818;
  assign n25234 = n28837 ^ n26404;
  assign n28836 = n28844 & n28845;
  assign n27738 = ~n28848;
  assign n28849 = n28861 & n28862;
  assign n28776 = n9 ^ n28793;
  assign n28806 = n28778 & n8;
  assign n28811 = n28820 & n28821;
  assign n28805 = ~n28778;
  assign n28769 = n28822 ^ n25234;
  assign n28823 = n25234 & n27706;
  assign n25267 = ~n25234;
  assign n28830 = ~n28836;
  assign n28838 = ~n28849;
  assign n27375 = n28775 ^ n28776;
  assign n28737 = n28776 & n28787;
  assign n28796 = n28805 & n20542;
  assign n28756 = ~n28806;
  assign n28799 = n28769 & n28750;
  assign n28794 = ~n28811;
  assign n28797 = ~n28769;
  assign n27689 = ~n28823;
  assign n28812 = n25267 & n28824;
  assign n28807 = n28830 & n28831;
  assign n28825 = n28838 & n28839;
  assign n28518 = ~n27375;
  assign n28777 = n28794 & n28795;
  assign n28780 = ~n28796;
  assign n28792 = n28797 & n28798;
  assign n28771 = ~n28799;
  assign n28788 = n28807 ^ n28808;
  assign n27708 = ~n28812;
  assign n28809 = ~n28807;
  assign n28802 = n28825 ^ n26344;
  assign n28826 = ~n28825;
  assign n28754 = n28777 ^ n28778;
  assign n28716 = n28788 ^ n28789;
  assign n28779 = ~n28777;
  assign n28752 = ~n28792;
  assign n25194 = n28801 ^ n28802;
  assign n28800 = n28809 & n28810;
  assign n28813 = n28826 & n28827;
  assign n28738 = n8 ^ n28754;
  assign n28766 = n28716 & n20485;
  assign n28772 = n28779 & n28780;
  assign n28767 = ~n28716;
  assign n28731 = n28781 ^ n25194;
  assign n28783 = n25194 & n27650;
  assign n25293 = ~n25194;
  assign n28790 = ~n28800;
  assign n28803 = ~n28813;
  assign n27310 = n28737 ^ n28738;
  assign n28739 = ~n28738;
  assign n28742 = ~n28766;
  assign n28757 = n28767 & n23;
  assign n28760 = n28731 & n28711;
  assign n28755 = ~n28772;
  assign n28758 = ~n28731;
  assign n28773 = n25293 & n28782;
  assign n27652 = ~n28783;
  assign n28768 = n28790 & n28791;
  assign n28784 = n28803 & n28804;
  assign n28470 = ~n27310;
  assign n28696 = n28739 & n28737;
  assign n28740 = n28755 & n28756;
  assign n28718 = ~n28757;
  assign n28753 = n28758 & n28759;
  assign n28713 = ~n28760;
  assign n28749 = n28768 ^ n28769;
  assign n27672 = ~n28773;
  assign n28770 = ~n28768;
  assign n28762 = n28784 ^ n26278;
  assign n28785 = ~n28784;
  assign n28699 = ~n28696;
  assign n28715 = n23 ^ n28740;
  assign n28701 = n28749 ^ n28750;
  assign n28741 = ~n28740;
  assign n28733 = ~n28753;
  assign n25178 = n28762 ^ n28763;
  assign n28761 = n28770 & n28771;
  assign n28774 = n28785 & n28786;
  assign n28697 = n28715 ^ n28716;
  assign n28728 = n28701 & n20442;
  assign n28734 = n28741 & n28742;
  assign n28729 = ~n28701;
  assign n28670 = n28743 ^ n25178;
  assign n28745 = n25178 & n27616;
  assign n25180 = ~n25178;
  assign n28751 = ~n28761;
  assign n28764 = ~n28774;
  assign n27206 = n28696 ^ n28697;
  assign n28698 = ~n28697;
  assign n28703 = ~n28728;
  assign n28719 = n28729 & n22;
  assign n28720 = n28670 & n28690;
  assign n28717 = ~n28734;
  assign n28721 = ~n28670;
  assign n28735 = n25180 & n28744;
  assign n27636 = ~n28745;
  assign n28730 = n28751 & n28752;
  assign n28746 = n28764 & n28765;
  assign n28431 = ~n27206;
  assign n28657 = n28698 & n28699;
  assign n28700 = n28717 & n28718;
  assign n28677 = ~n28719;
  assign n28692 = ~n28720;
  assign n28714 = n28721 & n28722;
  assign n28710 = n28730 ^ n28731;
  assign n27619 = ~n28735;
  assign n28732 = ~n28730;
  assign n28724 = n28746 ^ n26171;
  assign n28747 = ~n28746;
  assign n28668 = ~n28657;
  assign n28675 = n28700 ^ n28701;
  assign n28660 = n28710 ^ n28711;
  assign n28702 = ~n28700;
  assign n28672 = ~n28714;
  assign n25182 = n28724 ^ n28725;
  assign n28723 = n28732 & n28733;
  assign n28736 = n28747 & n28748;
  assign n28658 = n22 ^ n28675;
  assign n28686 = n28660 & n20379;
  assign n28693 = n28702 & n28703;
  assign n28687 = ~n28660;
  assign n28632 = n25182 ^ n28704;
  assign n28706 = n25182 & n27575;
  assign n25129 = ~n25182;
  assign n28712 = ~n28723;
  assign n28726 = ~n28736;
  assign n27140 = n28657 ^ n28658;
  assign n28619 = n28658 & n28668;
  assign n28662 = ~n28686;
  assign n28678 = n28687 & n21;
  assign n28680 = n28632 & n28688;
  assign n28676 = ~n28693;
  assign n28679 = ~n28632;
  assign n28694 = n25129 & n28705;
  assign n27577 = ~n28706;
  assign n28689 = n28712 & n28713;
  assign n28707 = n28726 & n28727;
  assign n28383 = ~n27140;
  assign n28659 = n28676 & n28677;
  assign n28638 = ~n28678;
  assign n28674 = n28679 & n28651;
  assign n28634 = ~n28680;
  assign n28669 = n28689 ^ n28690;
  assign n27600 = ~n28694;
  assign n28691 = ~n28689;
  assign n28683 = n28707 ^ n26099;
  assign n28708 = ~n28707;
  assign n28636 = n28659 ^ n28660;
  assign n28622 = n28669 ^ n28670;
  assign n28661 = ~n28659;
  assign n28653 = ~n28674;
  assign n25088 = n28682 ^ n28683;
  assign n28681 = n28691 & n28692;
  assign n28695 = n28708 & n28709;
  assign n28620 = n21 ^ n28636;
  assign n28647 = n28622 & n20341;
  assign n28654 = n28661 & n28662;
  assign n28648 = ~n28622;
  assign n28593 = n28663 ^ n25088;
  assign n28664 = n25088 & n28673;
  assign n25144 = ~n25088;
  assign n28671 = ~n28681;
  assign n28684 = ~n28695;
  assign n27066 = n28619 ^ n28620;
  assign n28580 = n28620 & n28619;
  assign n28623 = ~n28647;
  assign n28639 = n28648 & n20;
  assign n28640 = n28593 & n28649;
  assign n28637 = ~n28654;
  assign n28641 = ~n28593;
  assign n28655 = n25144 & n27534;
  assign n27537 = ~n28664;
  assign n28650 = n28671 & n28672;
  assign n28665 = n28684 & n28685;
  assign n28321 = ~n27066;
  assign n28621 = n28637 & n28638;
  assign n28600 = ~n28639;
  assign n28595 = ~n28640;
  assign n28635 = n28641 & n28613;
  assign n28631 = n28650 ^ n28651;
  assign n27559 = ~n28655;
  assign n28652 = ~n28650;
  assign n28643 = n28665 ^ n26016;
  assign n28666 = ~n28665;
  assign n28598 = n28621 ^ n28622;
  assign n28583 = n28631 ^ n28632;
  assign n28624 = ~n28621;
  assign n28615 = ~n28635;
  assign n25056 = n28643 ^ n28644;
  assign n28642 = n28652 & n28653;
  assign n28656 = n28666 & n28667;
  assign n28581 = n20 ^ n28598;
  assign n28610 = n28583 & n19;
  assign n28616 = n28623 & n28624;
  assign n28609 = ~n28583;
  assign n28552 = n28625 ^ n25056;
  assign n28626 = n25056 & n27502;
  assign n25100 = ~n25056;
  assign n28633 = ~n28642;
  assign n28645 = ~n28656;
  assign n26993 = n28580 ^ n28581;
  assign n28539 = n28581 & n28580;
  assign n28601 = n28609 & n20295;
  assign n28560 = ~n28610;
  assign n28603 = n28552 & n28611;
  assign n28599 = ~n28616;
  assign n28602 = ~n28552;
  assign n27504 = ~n28626;
  assign n28617 = n25100 & n28627;
  assign n28612 = n28633 & n28634;
  assign n28628 = n28645 & n28646;
  assign n28272 = ~n26993;
  assign n28582 = n28599 & n28600;
  assign n28585 = ~n28601;
  assign n28597 = n28602 & n28573;
  assign n28554 = ~n28603;
  assign n28592 = n28612 ^ n28613;
  assign n27516 = ~n28617;
  assign n28614 = ~n28612;
  assign n28605 = n28628 ^ n25989;
  assign n28629 = ~n28628;
  assign n28558 = n28582 ^ n28583;
  assign n28543 = n28592 ^ n28593;
  assign n28584 = ~n28582;
  assign n28575 = ~n28597;
  assign n25012 = n28605 ^ n28606;
  assign n28604 = n28614 & n28615;
  assign n28618 = n28629 & n28630;
  assign n28540 = n19 ^ n28558;
  assign n28571 = n28543 & n18;
  assign n28577 = n28584 & n28585;
  assign n28570 = ~n28543;
  assign n28515 = n28586 ^ n25012;
  assign n28587 = n25012 & n28596;
  assign n25049 = ~n25012;
  assign n28594 = ~n28604;
  assign n28607 = ~n28618;
  assign n26925 = n28539 ^ n28540;
  assign n28541 = ~n28540;
  assign n28561 = n28570 & n20271;
  assign n28521 = ~n28571;
  assign n28562 = n28515 & n28530;
  assign n28559 = ~n28577;
  assign n28563 = ~n28515;
  assign n27480 = ~n28587;
  assign n28578 = n25049 & n27453;
  assign n28572 = n28594 & n28595;
  assign n28588 = n28607 & n28608;
  assign n28502 = n28541 & n28539;
  assign n28542 = n28559 & n28560;
  assign n28544 = ~n28561;
  assign n28532 = ~n28562;
  assign n28555 = n28563 & n28564;
  assign n28551 = n28572 ^ n28573;
  assign n27456 = ~n28578;
  assign n28574 = ~n28572;
  assign n24958 = n28588 ^ n28589;
  assign n28590 = ~n28588;
  assign n28513 = ~n28502;
  assign n28519 = n28542 ^ n28543;
  assign n28505 = n28551 ^ n28552;
  assign n28545 = ~n28542;
  assign n28517 = ~n28555;
  assign n28565 = n28574 & n28575;
  assign n28567 = n24958 & n28576;
  assign n25044 = ~n24958;
  assign n28579 = n28590 & n28591;
  assign n28503 = n18 ^ n28519;
  assign n28528 = n28505 & n17;
  assign n28534 = n28544 & n28545;
  assign n28527 = ~n28505;
  assign n28496 = n28556 ^ n25044;
  assign n28553 = ~n28565;
  assign n28557 = n25044 & n28566;
  assign n27402 = ~n28567;
  assign n28568 = ~n28579;
  assign n26628 = n28502 ^ n28503;
  assign n28461 = n28503 & n28513;
  assign n28522 = n28527 & n20212;
  assign n28483 = ~n28528;
  assign n28520 = ~n28534;
  assign n28535 = n28496 & n28546;
  assign n28529 = n28553 & n28554;
  assign n28536 = ~n28496;
  assign n27432 = ~n28557;
  assign n28547 = n28568 & n28569;
  assign n24728 = n26604 ^ n26628;
  assign n28458 = n28480 ^ n26628;
  assign n28389 = n26628 & n26604;
  assign n28464 = ~n28461;
  assign n28504 = n28520 & n28521;
  assign n28507 = ~n28522;
  assign n28514 = n28529 ^ n28530;
  assign n28498 = ~n28535;
  assign n28533 = n28536 & n28476;
  assign n28531 = ~n28529;
  assign n28537 = n27432 & n27402;
  assign n28524 = n28547 ^ n28548;
  assign n28549 = ~n28547;
  assign n26535 = n103 ^ n28458;
  assign n28160 = n28458 & n103;
  assign n28459 = ~n28458;
  assign n28481 = n28504 ^ n28505;
  assign n28466 = n28514 ^ n28515;
  assign n28506 = ~n28504;
  assign n24924 = n28524 ^ n25833;
  assign n28523 = n28531 & n28532;
  assign n28478 = ~n28533;
  assign n27430 = ~n28537;
  assign n28538 = n28549 & n28550;
  assign n27728 = ~n26535;
  assign n28251 = n28459 & n28460;
  assign n28462 = n17 ^ n28481;
  assign n28493 = n28466 & n20204;
  assign n28499 = n28506 & n28507;
  assign n28494 = ~n28466;
  assign n28452 = n28508 ^ n24924;
  assign n28509 = n24924 & n28518;
  assign n25023 = ~n24924;
  assign n28516 = ~n28523;
  assign n28525 = ~n28538;
  assign n28447 = n28461 ^ n28462;
  assign n28463 = ~n28462;
  assign n28468 = ~n28493;
  assign n28484 = n28494 & n16;
  assign n28485 = n28452 & n28428;
  assign n28482 = ~n28499;
  assign n28486 = ~n28452;
  assign n28500 = n25023 & n27375;
  assign n27346 = ~n28509;
  assign n28495 = n28516 & n28517;
  assign n28510 = n28525 & n28526;
  assign n28435 = n28447 & n26483;
  assign n28434 = ~n28447;
  assign n28416 = n28463 & n28464;
  assign n28465 = n28482 & n28483;
  assign n28438 = ~n28484;
  assign n28430 = ~n28485;
  assign n28479 = n28486 & n28487;
  assign n28475 = n28495 ^ n28496;
  assign n27377 = ~n28500;
  assign n28497 = ~n28495;
  assign n28489 = n28510 ^ n25769;
  assign n28511 = ~n28510;
  assign n28432 = n28434 & n26470;
  assign n28391 = ~n28435;
  assign n28419 = ~n28416;
  assign n28436 = n28465 ^ n28466;
  assign n28395 = n28475 ^ n28476;
  assign n28467 = ~n28465;
  assign n28454 = ~n28479;
  assign n24882 = n28489 ^ n28490;
  assign n28488 = n28497 & n28498;
  assign n28501 = n28511 & n28512;
  assign n28415 = ~n28432;
  assign n28417 = n16 ^ n28436;
  assign n28449 = n28395 & n31;
  assign n28455 = n28467 & n28468;
  assign n28448 = ~n28395;
  assign n28407 = n28469 ^ n24882;
  assign n28471 = n24882 & n27310;
  assign n24982 = ~n24882;
  assign n28477 = ~n28488;
  assign n28491 = ~n28501;
  assign n28410 = n28415 & n28389;
  assign n28388 = n28415 & n28391;
  assign n28334 = n28416 ^ n28417;
  assign n28418 = ~n28417;
  assign n28439 = n28448 & n20137;
  assign n28397 = ~n28449;
  assign n28440 = n28407 & n28450;
  assign n28437 = ~n28455;
  assign n28441 = ~n28407;
  assign n28456 = n24982 & n28470;
  assign n27312 = ~n28471;
  assign n28451 = n28477 & n28478;
  assign n28472 = n28491 & n28492;
  assign n24675 = n28388 ^ n28389;
  assign n28392 = n28334 & n26430;
  assign n28390 = ~n28410;
  assign n28393 = ~n28334;
  assign n28365 = n28418 & n28419;
  assign n28420 = n28437 & n28438;
  assign n28422 = ~n28439;
  assign n28409 = ~n28440;
  assign n28433 = n28441 & n28379;
  assign n28427 = n28451 ^ n28452;
  assign n27280 = ~n28456;
  assign n28453 = ~n28451;
  assign n28444 = n28472 ^ n25692;
  assign n28473 = ~n28472;
  assign n27443 = n26483 ^ n24675;
  assign n24715 = ~n24675;
  assign n28362 = n28390 & n28391;
  assign n28363 = ~n28392;
  assign n28384 = n28393 & n26379;
  assign n28368 = ~n28365;
  assign n28394 = n31 ^ n28420;
  assign n28370 = n28427 ^ n28428;
  assign n28421 = ~n28420;
  assign n28381 = ~n28433;
  assign n24865 = n28443 ^ n28444;
  assign n28442 = n28453 & n28454;
  assign n28457 = n28473 & n28474;
  assign n28326 = n27443 ^ n27434;
  assign n28335 = n28362 ^ n26379;
  assign n28364 = ~n28362;
  assign n28337 = ~n28384;
  assign n28366 = n28394 ^ n28395;
  assign n28404 = n28370 & n20098;
  assign n28411 = n28421 & n28422;
  assign n28405 = ~n28370;
  assign n28423 = n24865 & n28431;
  assign n24908 = ~n24865;
  assign n28429 = ~n28442;
  assign n28445 = ~n28457;
  assign n28308 = n28326 & n28327;
  assign n28306 = ~n28326;
  assign n24670 = n28334 ^ n28335;
  assign n28358 = n28363 & n28364;
  assign n28277 = n28365 ^ n28366;
  assign n28367 = ~n28366;
  assign n28372 = ~n28404;
  assign n28398 = n28405 & n30;
  assign n28396 = ~n28411;
  assign n28329 = n28412 ^ n24908;
  assign n27209 = ~n28423;
  assign n28413 = n24908 & n27206;
  assign n28406 = n28429 & n28430;
  assign n28424 = n28445 & n28446;
  assign n28301 = n28306 & n28307;
  assign n28253 = ~n28308;
  assign n27364 = n24670 ^ n26379;
  assign n24666 = ~n24670;
  assign n28339 = n28277 & n26336;
  assign n28336 = ~n28358;
  assign n28338 = ~n28277;
  assign n28312 = n28367 & n28368;
  assign n28369 = n28396 & n28397;
  assign n28342 = ~n28398;
  assign n28387 = n28329 & n28355;
  assign n28378 = n28406 ^ n28407;
  assign n28385 = ~n28329;
  assign n27243 = ~n28413;
  assign n28408 = ~n28406;
  assign n28401 = n28424 ^ n25564;
  assign n28425 = ~n28424;
  assign n28183 = n27364 ^ n27325;
  assign n28276 = ~n28301;
  assign n28309 = n28336 & n28337;
  assign n28332 = n28338 & n26330;
  assign n28280 = ~n28339;
  assign n28315 = ~n28312;
  assign n28340 = n28369 ^ n28370;
  assign n28317 = n28378 ^ n28379;
  assign n28371 = ~n28369;
  assign n28382 = n28385 & n28386;
  assign n28357 = ~n28387;
  assign n24916 = n28400 ^ n28401;
  assign n28399 = n28408 & n28409;
  assign n28414 = n28425 & n28426;
  assign n28247 = n28183 & n28213;
  assign n28248 = ~n28183;
  assign n28273 = n28276 & n28251;
  assign n28250 = n28276 & n28253;
  assign n28278 = n28309 ^ n26330;
  assign n28310 = ~n28309;
  assign n28311 = ~n28332;
  assign n28313 = n30 ^ n28340;
  assign n28352 = n28317 & n29;
  assign n28359 = n28371 & n28372;
  assign n28351 = ~n28317;
  assign n28269 = n28373 ^ n24916;
  assign n28331 = ~n28382;
  assign n28374 = n24916 & n28383;
  assign n24828 = ~n24916;
  assign n28380 = ~n28399;
  assign n28402 = ~n28414;
  assign n28189 = ~n28247;
  assign n28242 = n28248 & n28249;
  assign n28235 = n28250 ^ n28251;
  assign n28252 = ~n28273;
  assign n24620 = n28277 ^ n28278;
  assign n28302 = n28310 & n28311;
  assign n28219 = n28312 ^ n28313;
  assign n28314 = ~n28313;
  assign n28343 = n28351 & n20052;
  assign n28285 = ~n28352;
  assign n28345 = n28269 & n28353;
  assign n28341 = ~n28359;
  assign n28344 = ~n28269;
  assign n28360 = n24828 & n27140;
  assign n27142 = ~n28374;
  assign n28354 = n28380 & n28381;
  assign n28375 = n28402 & n28403;
  assign n28218 = n28235 & n102;
  assign n28216 = ~n28242;
  assign n28217 = ~n28235;
  assign n28243 = n28252 & n28253;
  assign n27281 = n26336 ^ n24620;
  assign n24630 = ~n24620;
  assign n28282 = n28219 & n26232;
  assign n28279 = ~n28302;
  assign n28281 = ~n28219;
  assign n28257 = n28314 & n28315;
  assign n28316 = n28341 & n28342;
  assign n28319 = ~n28343;
  assign n28333 = n28344 & n28298;
  assign n28271 = ~n28345;
  assign n28328 = n28354 ^ n28355;
  assign n27174 = ~n28360;
  assign n28356 = ~n28354;
  assign n28348 = n28375 ^ n25541;
  assign n28376 = ~n28375;
  assign n28211 = n28217 & n14810;
  assign n28164 = ~n28218;
  assign n28128 = n27281 ^ n27221;
  assign n28212 = ~n28243;
  assign n28254 = n28279 & n28280;
  assign n28274 = n28281 & n26235;
  assign n28255 = ~n28282;
  assign n28260 = ~n28257;
  assign n28283 = n28316 ^ n28317;
  assign n28262 = n28328 ^ n28329;
  assign n28318 = ~n28316;
  assign n28300 = ~n28333;
  assign n24831 = n28347 ^ n28348;
  assign n28346 = n28356 & n28357;
  assign n28361 = n28376 & n28377;
  assign n28193 = n28128 & n28158;
  assign n28190 = ~n28211;
  assign n28191 = ~n28128;
  assign n28182 = n28212 ^ n28213;
  assign n28210 = n28216 & n28212;
  assign n28220 = n28254 ^ n26235;
  assign n28256 = ~n28254;
  assign n28222 = ~n28274;
  assign n28258 = n29 ^ n28283;
  assign n28295 = n28262 & n20006;
  assign n28303 = n28318 & n28319;
  assign n28296 = ~n28262;
  assign n28207 = n28320 ^ n24831;
  assign n28322 = n24831 & n27066;
  assign n24795 = ~n24831;
  assign n28330 = ~n28346;
  assign n28349 = ~n28361;
  assign n28124 = n28182 ^ n28183;
  assign n28184 = n28190 & n28160;
  assign n28159 = n28190 & n28164;
  assign n28185 = n28191 & n28192;
  assign n28132 = ~n28193;
  assign n28188 = ~n28210;
  assign n24591 = n28219 ^ n28220;
  assign n28244 = n28255 & n28256;
  assign n28166 = n28257 ^ n28258;
  assign n28259 = ~n28258;
  assign n28264 = ~n28295;
  assign n28286 = n28296 & n28;
  assign n28287 = n28207 & n28239;
  assign n28284 = ~n28303;
  assign n28288 = ~n28207;
  assign n28304 = n24795 & n28321;
  assign n27068 = ~n28322;
  assign n28297 = n28330 & n28331;
  assign n28323 = n28349 & n28350;
  assign n28153 = n28124 & n101;
  assign n28130 = n28159 ^ n28160;
  assign n28152 = ~n28124;
  assign n28163 = ~n28184;
  assign n28161 = ~n28185;
  assign n28157 = n28188 & n28189;
  assign n27213 = n24591 ^ n26235;
  assign n24588 = ~n24591;
  assign n28223 = n28166 & n26216;
  assign n28221 = ~n28244;
  assign n28224 = ~n28166;
  assign n28197 = n28259 & n28260;
  assign n28261 = n28284 & n28285;
  assign n28227 = ~n28286;
  assign n28241 = ~n28287;
  assign n28275 = n28288 & n28289;
  assign n28268 = n28297 ^ n28298;
  assign n27108 = ~n28304;
  assign n28299 = ~n28297;
  assign n28292 = n28323 ^ n25465;
  assign n28324 = ~n28323;
  assign n26490 = n28130 ^ n27728;
  assign n28067 = n28130 & n26535;
  assign n28147 = n28152 & n14752;
  assign n28099 = ~n28153;
  assign n28129 = n28157 ^ n28158;
  assign n28155 = n28163 & n28164;
  assign n28076 = n27213 ^ n27146;
  assign n28162 = ~n28157;
  assign n28194 = n28221 & n28222;
  assign n28168 = ~n28223;
  assign n28214 = n28224 & n26143;
  assign n28200 = ~n28197;
  assign n28225 = n28261 ^ n28262;
  assign n28202 = n28268 ^ n28269;
  assign n28263 = ~n28261;
  assign n28209 = ~n28275;
  assign n24766 = n28291 ^ n28292;
  assign n28290 = n28299 & n28300;
  assign n28305 = n28324 & n28325;
  assign n27679 = ~n26490;
  assign n28065 = n28128 ^ n28129;
  assign n28071 = ~n28067;
  assign n28122 = ~n28147;
  assign n28133 = n28076 & n28105;
  assign n28123 = ~n28155;
  assign n28134 = ~n28076;
  assign n28154 = n28161 & n28162;
  assign n28165 = n28194 ^ n26143;
  assign n28195 = ~n28194;
  assign n28196 = ~n28214;
  assign n28198 = n28 ^ n28225;
  assign n28237 = n28202 & n27;
  assign n28245 = n28263 & n28264;
  assign n28236 = ~n28202;
  assign n28149 = n28265 ^ n24766;
  assign n28266 = n24766 & n28272;
  assign n24836 = ~n24766;
  assign n28270 = ~n28290;
  assign n28293 = ~n28305;
  assign n28102 = n28065 & n14710;
  assign n28103 = ~n28065;
  assign n28118 = n28122 & n28123;
  assign n28097 = n28123 ^ n28124;
  assign n28107 = ~n28133;
  assign n28125 = n28134 & n28135;
  assign n28131 = ~n28154;
  assign n24536 = n28165 ^ n28166;
  assign n28186 = n28195 & n28196;
  assign n28108 = n28197 ^ n28198;
  assign n28199 = ~n28198;
  assign n28228 = n28236 & n19971;
  assign n28173 = ~n28237;
  assign n28231 = n28149 & n28179;
  assign n28226 = ~n28245;
  assign n28229 = ~n28149;
  assign n28246 = n24836 & n26993;
  assign n27034 = ~n28266;
  assign n28238 = n28270 & n28271;
  assign n28267 = n28293 & n28294;
  assign n28068 = n101 ^ n28097;
  assign n28069 = ~n28102;
  assign n28096 = n28103 & n100;
  assign n28098 = ~n28118;
  assign n28078 = ~n28125;
  assign n28104 = n28131 & n28132;
  assign n27130 = n24536 ^ n26216;
  assign n24566 = ~n24536;
  assign n28169 = n28108 & n26074;
  assign n28167 = ~n28186;
  assign n28170 = ~n28108;
  assign n28139 = n28199 & n28200;
  assign n28201 = n28226 & n28227;
  assign n28204 = ~n28228;
  assign n28215 = n28229 & n28230;
  assign n28181 = ~n28231;
  assign n28206 = n28238 ^ n28239;
  assign n26996 = ~n28246;
  assign n28240 = ~n28238;
  assign n28234 = n28267 ^ n26860;
  assign n26405 = n28067 ^ n28068;
  assign n28070 = ~n28068;
  assign n28045 = ~n28096;
  assign n28092 = n28098 & n28099;
  assign n28075 = n28104 ^ n28105;
  assign n28029 = n27130 ^ n27115;
  assign n28106 = ~n28104;
  assign n28136 = n28167 & n28168;
  assign n28137 = ~n28169;
  assign n28156 = n28170 & n26158;
  assign n28142 = ~n28139;
  assign n28171 = n28201 ^ n28202;
  assign n28144 = n28206 ^ n28207;
  assign n28203 = ~n28201;
  assign n28151 = ~n28215;
  assign n24783 = n28233 ^ n28234;
  assign n28232 = n28240 & n28241;
  assign n27643 = ~n26405;
  assign n28017 = n28070 & n28071;
  assign n28023 = n28075 ^ n28076;
  assign n28064 = ~n28092;
  assign n28079 = n28029 & n28093;
  assign n28080 = ~n28029;
  assign n28100 = n28106 & n28107;
  assign n28109 = n28136 ^ n26158;
  assign n28138 = ~n28136;
  assign n28111 = ~n28156;
  assign n28140 = n27 ^ n28171;
  assign n28176 = n28144 & n19943;
  assign n28187 = n28203 & n28204;
  assign n28177 = ~n28144;
  assign n28095 = n28205 ^ n24783;
  assign n28208 = ~n28232;
  assign n28049 = n28023 & n14678;
  assign n28020 = ~n28017;
  assign n28043 = n28064 ^ n28065;
  assign n28063 = n28069 & n28064;
  assign n28050 = ~n28023;
  assign n28031 = ~n28079;
  assign n28072 = n28080 & n28052;
  assign n28077 = ~n28100;
  assign n24540 = n28108 ^ n28109;
  assign n28126 = n28137 & n28138;
  assign n28056 = n28139 ^ n28140;
  assign n28141 = ~n28140;
  assign n28146 = ~n28176;
  assign n28174 = n28177 & n26;
  assign n28172 = ~n28187;
  assign n28178 = n28208 & n28209;
  assign n28018 = n100 ^ n28043;
  assign n28024 = ~n28049;
  assign n28046 = n28050 & n99;
  assign n28044 = ~n28063;
  assign n28054 = ~n28072;
  assign n28051 = n28077 & n28078;
  assign n27056 = n24540 ^ n26158;
  assign n24509 = ~n24540;
  assign n28112 = n28056 & n26056;
  assign n28110 = ~n28126;
  assign n28113 = ~n28056;
  assign n28084 = n28141 & n28142;
  assign n28143 = n28172 & n28173;
  assign n28116 = ~n28174;
  assign n28148 = n28178 ^ n28179;
  assign n28180 = ~n28178;
  assign n26347 = n28017 ^ n28018;
  assign n28019 = ~n28018;
  assign n28022 = n28044 & n28045;
  assign n27999 = ~n28046;
  assign n28028 = n28051 ^ n28052;
  assign n27986 = n27056 ^ n27040;
  assign n28053 = ~n28051;
  assign n28081 = n28110 & n28111;
  assign n28058 = ~n28112;
  assign n28101 = n28113 & n25998;
  assign n28087 = ~n28084;
  assign n28114 = n28143 ^ n28144;
  assign n28089 = n28148 ^ n28149;
  assign n28145 = ~n28143;
  assign n28175 = n28180 & n28181;
  assign n27608 = ~n26347;
  assign n27976 = n28019 & n28020;
  assign n27997 = n28022 ^ n28023;
  assign n27979 = n28028 ^ n28029;
  assign n28025 = ~n28022;
  assign n28032 = n27986 & n28006;
  assign n28033 = ~n27986;
  assign n28047 = n28053 & n28054;
  assign n28055 = n28081 ^ n25998;
  assign n28082 = ~n28081;
  assign n28083 = ~n28101;
  assign n28085 = n26 ^ n28114;
  assign n28119 = n28089 & n19881;
  assign n28127 = n28145 & n28146;
  assign n28120 = ~n28089;
  assign n28150 = ~n28175;
  assign n27977 = n99 ^ n27997;
  assign n28004 = n27979 & n98;
  assign n28021 = n28024 & n28025;
  assign n28003 = ~n27979;
  assign n27988 = ~n28032;
  assign n28026 = n28033 & n28034;
  assign n28030 = ~n28047;
  assign n24507 = n28055 ^ n28056;
  assign n28073 = n28082 & n28083;
  assign n28066 = n28084 ^ n28085;
  assign n28086 = ~n28085;
  assign n28091 = ~n28119;
  assign n28117 = n28120 & n25;
  assign n28115 = ~n28127;
  assign n28121 = n28150 & n28151;
  assign n26279 = n27976 ^ n27977;
  assign n27942 = n27977 & n27976;
  assign n28000 = n28003 & n14640;
  assign n27962 = ~n28004;
  assign n27998 = ~n28021;
  assign n28008 = ~n28026;
  assign n28005 = n28030 & n28031;
  assign n26969 = n24507 ^ n26056;
  assign n24479 = ~n24507;
  assign n28059 = n28066 & n25925;
  assign n28057 = ~n28073;
  assign n28009 = ~n28066;
  assign n28038 = n28086 & n28087;
  assign n28088 = n28115 & n28116;
  assign n28062 = ~n28117;
  assign n28094 = n24 ^ n28121;
  assign n27556 = ~n26279;
  assign n27978 = n27998 & n27999;
  assign n27981 = ~n28000;
  assign n27985 = n28005 ^ n28006;
  assign n27954 = n26969 ^ n26912;
  assign n28007 = ~n28005;
  assign n28035 = n28057 & n28058;
  assign n28037 = ~n28059;
  assign n28048 = n28009 & n26002;
  assign n28060 = n28088 ^ n28089;
  assign n28042 = n28094 ^ n28095;
  assign n28090 = ~n28088;
  assign n27960 = n27978 ^ n27979;
  assign n27946 = n27985 ^ n27986;
  assign n27980 = ~n27978;
  assign n27989 = n27954 & n27968;
  assign n27990 = ~n27954;
  assign n28001 = n28007 & n28008;
  assign n28010 = n28035 ^ n26002;
  assign n28036 = ~n28035;
  assign n28012 = ~n28048;
  assign n28039 = n25 ^ n28060;
  assign n28074 = n28090 & n28091;
  assign n27943 = n98 ^ n27960;
  assign n27965 = n27946 & n14600;
  assign n27975 = n27980 & n27981;
  assign n27966 = ~n27946;
  assign n27956 = ~n27989;
  assign n27982 = n27990 & n27991;
  assign n27987 = ~n28001;
  assign n24444 = n28009 ^ n28010;
  assign n28027 = n28036 & n28037;
  assign n27972 = n28038 ^ n28039;
  assign n28040 = ~n28039;
  assign n28061 = ~n28074;
  assign n26244 = n27942 ^ n27943;
  assign n27944 = ~n27943;
  assign n27948 = ~n27965;
  assign n27963 = n27966 & n97;
  assign n27961 = ~n27975;
  assign n27970 = ~n27982;
  assign n27967 = n27987 & n27988;
  assign n24470 = ~n24444;
  assign n28014 = n27972 & n25855;
  assign n28011 = ~n28027;
  assign n28013 = ~n27972;
  assign n28015 = n28040 & n28038;
  assign n28041 = n28061 & n28062;
  assign n27532 = ~n26244;
  assign n27907 = n27944 & n27942;
  assign n27945 = n27961 & n27962;
  assign n27928 = ~n27963;
  assign n27953 = n27967 ^ n27968;
  assign n27969 = ~n27967;
  assign n26900 = n24470 ^ n26002;
  assign n27992 = n28011 & n28012;
  assign n28002 = n28013 & n25853;
  assign n27974 = ~n28014;
  assign n28016 = n28041 ^ n28042;
  assign n27926 = n27945 ^ n27946;
  assign n27910 = n27953 ^ n27954;
  assign n27947 = ~n27945;
  assign n27918 = n26900 ^ n26877;
  assign n27964 = n27969 & n27970;
  assign n27971 = n27992 ^ n25853;
  assign n27993 = ~n27992;
  assign n27994 = ~n28002;
  assign n27936 = n28015 ^ n28016;
  assign n27908 = n97 ^ n27926;
  assign n27932 = n27910 & n14563;
  assign n27940 = n27947 & n27948;
  assign n27933 = ~n27910;
  assign n27951 = n27918 & n27935;
  assign n27949 = ~n27918;
  assign n27955 = ~n27964;
  assign n24442 = n27971 ^ n27972;
  assign n27983 = n27993 & n27994;
  assign n27995 = n27936 & n25747;
  assign n27996 = ~n27936;
  assign n26136 = n27907 ^ n27908;
  assign n27871 = n27908 & n27907;
  assign n27912 = ~n27932;
  assign n27929 = n27933 & n96;
  assign n27927 = ~n27940;
  assign n27941 = n27949 & n27950;
  assign n27914 = ~n27951;
  assign n27934 = n27955 & n27956;
  assign n26835 = n25855 ^ n24442;
  assign n24410 = ~n24442;
  assign n27973 = ~n27983;
  assign n27939 = ~n27995;
  assign n27984 = n27996 & n25745;
  assign n27476 = ~n26136;
  assign n27874 = ~n27871;
  assign n27909 = n27927 & n27928;
  assign n27894 = ~n27929;
  assign n27917 = n27934 ^ n27935;
  assign n27880 = n26835 ^ n26813;
  assign n27931 = ~n27941;
  assign n27930 = ~n27934;
  assign n27957 = n27973 & n27974;
  assign n27959 = ~n27984;
  assign n27892 = n27909 ^ n27910;
  assign n27876 = n27917 ^ n27918;
  assign n27911 = ~n27909;
  assign n27919 = n27880 & n27924;
  assign n27925 = n27930 & n27931;
  assign n27920 = ~n27880;
  assign n27937 = n27957 ^ n25747;
  assign n27958 = ~n27957;
  assign n27872 = n96 ^ n27892;
  assign n27900 = n27876 & n14517;
  assign n27906 = n27911 & n27912;
  assign n27901 = ~n27876;
  assign n27882 = ~n27919;
  assign n27915 = n27920 & n27897;
  assign n27913 = ~n27925;
  assign n24372 = n27936 ^ n27937;
  assign n27952 = n27958 & n27959;
  assign n26065 = n27871 ^ n27872;
  assign n27873 = ~n27872;
  assign n27878 = ~n27900;
  assign n27895 = n27901 & n111;
  assign n27893 = ~n27906;
  assign n27896 = n27913 & n27914;
  assign n27899 = ~n27915;
  assign n26776 = n24372 ^ n25747;
  assign n24408 = ~n24372;
  assign n27938 = ~n27952;
  assign n27441 = ~n26065;
  assign n27836 = n27873 & n27874;
  assign n27875 = n27893 & n27894;
  assign n27859 = ~n27895;
  assign n27879 = n27896 ^ n27897;
  assign n27843 = n26776 ^ n26722;
  assign n27898 = ~n27896;
  assign n27921 = n27938 & n27939;
  assign n27849 = ~n27836;
  assign n27857 = n27875 ^ n27876;
  assign n27839 = n27879 ^ n27880;
  assign n27877 = ~n27875;
  assign n27885 = n27843 & n27889;
  assign n27890 = n27898 & n27899;
  assign n27886 = ~n27843;
  assign n27902 = n27921 ^ n25645;
  assign n27922 = ~n27921;
  assign n27837 = n111 ^ n27857;
  assign n27861 = n27839 & n110;
  assign n27860 = ~n27839;
  assign n27869 = n27877 & n27878;
  assign n27845 = ~n27885;
  assign n27883 = n27886 & n27863;
  assign n27881 = ~n27890;
  assign n24333 = n27902 ^ n27903;
  assign n27916 = n27922 & n27923;
  assign n25992 = n27836 ^ n27837;
  assign n27805 = n27837 & n27849;
  assign n27852 = n27860 & n14497;
  assign n27824 = ~n27861;
  assign n27858 = ~n27869;
  assign n27862 = n27881 & n27882;
  assign n27865 = ~n27883;
  assign n26725 = n25751 ^ n24333;
  assign n24359 = ~n24333;
  assign n27904 = ~n27916;
  assign n27408 = ~n25992;
  assign n27841 = ~n27852;
  assign n27838 = n27858 & n27859;
  assign n27842 = n27862 ^ n27863;
  assign n27813 = n26725 ^ n26706;
  assign n27864 = ~n27862;
  assign n27891 = n27904 & n27905;
  assign n27822 = n27838 ^ n27839;
  assign n27809 = n27842 ^ n27843;
  assign n27840 = ~n27838;
  assign n27850 = n27813 & n27853;
  assign n27854 = n27864 & n27865;
  assign n27851 = ~n27813;
  assign n27888 = n27891 & n25669;
  assign n27887 = ~n27891;
  assign n27806 = n110 ^ n27822;
  assign n27826 = n27809 & n109;
  assign n27825 = ~n27809;
  assign n27832 = n27840 & n27841;
  assign n27815 = ~n27850;
  assign n27846 = n27851 & n27828;
  assign n27844 = ~n27854;
  assign n27884 = n27887 & n25574;
  assign n27868 = ~n27888;
  assign n25955 = n27805 ^ n27806;
  assign n27807 = ~n27806;
  assign n27816 = n27825 & n14444;
  assign n27792 = ~n27826;
  assign n27823 = ~n27832;
  assign n27827 = n27844 & n27845;
  assign n27830 = ~n27846;
  assign n27867 = n27868 & n27870;
  assign n27856 = ~n27884;
  assign n27323 = ~n25955;
  assign n27773 = n27807 & n27805;
  assign n27811 = ~n27816;
  assign n27808 = n27823 & n27824;
  assign n27812 = n27827 ^ n27828;
  assign n27829 = ~n27827;
  assign n27855 = ~n27867;
  assign n27866 = n27856 & n27868;
  assign n27790 = n27808 ^ n27809;
  assign n27777 = n27812 ^ n27813;
  assign n27810 = ~n27808;
  assign n27817 = n27829 & n27830;
  assign n27833 = n27855 & n27856;
  assign n27848 = ~n27866;
  assign n27774 = n109 ^ n27790;
  assign n27794 = n27777 & n108;
  assign n27793 = ~n27777;
  assign n27801 = n27810 & n27811;
  assign n27814 = ~n27817;
  assign n27818 = n27833 ^ n25497;
  assign n24331 = n27847 ^ n27848;
  assign n27834 = ~n27833;
  assign n25842 = n27773 ^ n27774;
  assign n27775 = ~n27774;
  assign n27784 = n27793 & n14397;
  assign n27758 = ~n27794;
  assign n27791 = ~n27801;
  assign n27795 = n27814 & n27815;
  assign n24291 = n27818 ^ n27819;
  assign n26679 = n25574 ^ n24331;
  assign n27831 = n27834 & n27835;
  assign n24293 = ~n24331;
  assign n27240 = ~n25842;
  assign n27741 = n27775 & n27773;
  assign n27779 = ~n27784;
  assign n27776 = n27791 & n27792;
  assign n27781 = n27795 ^ n27796;
  assign n27783 = ~n27795;
  assign n26638 = n25589 ^ n24291;
  assign n27780 = n26679 ^ n26666;
  assign n24251 = ~n24291;
  assign n27820 = ~n27831;
  assign n27756 = n27776 ^ n27777;
  assign n27745 = n27780 ^ n27781;
  assign n27778 = ~n27776;
  assign n27719 = n26638 ^ n26622;
  assign n27797 = n27780 & n27796;
  assign n27798 = ~n27780;
  assign n27802 = n27820 & n27821;
  assign n27742 = n108 ^ n27756;
  assign n27759 = n27745 & n14377;
  assign n27760 = ~n27745;
  assign n27765 = n27778 & n27779;
  assign n27766 = n27719 & n27736;
  assign n27767 = ~n27719;
  assign n27762 = ~n27797;
  assign n27785 = n27798 & n27799;
  assign n27787 = n27802 ^ n25502;
  assign n27803 = ~n27802;
  assign n25808 = n27741 ^ n27742;
  assign n27743 = ~n27742;
  assign n27747 = ~n27759;
  assign n27750 = n27760 & n107;
  assign n27757 = ~n27765;
  assign n27727 = ~n27766;
  assign n27763 = n27767 & n27768;
  assign n27782 = ~n27785;
  assign n24239 = n27786 ^ n27787;
  assign n27800 = n27803 & n27804;
  assign n27186 = ~n25808;
  assign n27709 = n27743 & n27741;
  assign n27725 = ~n27750;
  assign n27744 = n27757 & n27758;
  assign n27749 = ~n27763;
  assign n26595 = n25502 ^ n24239;
  assign n27769 = n27782 & n27783;
  assign n24211 = ~n24239;
  assign n27788 = ~n27800;
  assign n27712 = ~n27709;
  assign n27723 = n27744 ^ n27745;
  assign n27746 = ~n27744;
  assign n27691 = n26595 ^ n26550;
  assign n27761 = ~n27769;
  assign n27770 = n27788 & n27789;
  assign n27710 = n107 ^ n27723;
  assign n27731 = n27746 & n27747;
  assign n27733 = n27691 & n27748;
  assign n27732 = ~n27691;
  assign n27751 = n27761 & n27762;
  assign n27753 = n27770 ^ n25364;
  assign n27771 = ~n27770;
  assign n27124 = n27709 ^ n27710;
  assign n27711 = ~n27710;
  assign n27724 = ~n27731;
  assign n27729 = n27732 & n27714;
  assign n27693 = ~n27733;
  assign n27735 = ~n27751;
  assign n24171 = n27752 ^ n27753;
  assign n27764 = n27771 & n27772;
  assign n25694 = ~n27124;
  assign n27660 = n27711 & n27712;
  assign n27700 = n27724 & n27725;
  assign n27716 = ~n27729;
  assign n27718 = n27735 ^ n27736;
  assign n27734 = n27749 & n27735;
  assign n24198 = ~n24171;
  assign n27754 = ~n27764;
  assign n27684 = ~n27700;
  assign n27701 = n27718 ^ n27719;
  assign n26533 = n24198 ^ n25364;
  assign n27726 = ~n27734;
  assign n27737 = n27754 & n27755;
  assign n27682 = n27700 ^ n27701;
  assign n27703 = n27701 & n106;
  assign n27654 = n26533 ^ n26497;
  assign n27702 = ~n27701;
  assign n27713 = n27726 & n27727;
  assign n24111 = n27737 ^ n27738;
  assign n27739 = ~n27737;
  assign n27661 = n106 ^ n27682;
  assign n27695 = n27702 & n14316;
  assign n27698 = n27654 & n27676;
  assign n27664 = ~n27703;
  assign n27690 = n27713 ^ n27714;
  assign n27696 = ~n27654;
  assign n27715 = ~n27713;
  assign n26488 = n25377 ^ n24111;
  assign n27720 = n24111 & n27728;
  assign n24169 = ~n24111;
  assign n27730 = n27739 & n27740;
  assign n25618 = n27660 ^ n27661;
  assign n27620 = n27661 & n27660;
  assign n27648 = n27690 ^ n27691;
  assign n27683 = ~n27695;
  assign n27694 = n27696 & n27697;
  assign n27677 = ~n27698;
  assign n27640 = n26488 ^ n26412;
  assign n27704 = n27715 & n27716;
  assign n26514 = ~n27720;
  assign n27717 = n24169 & n26535;
  assign n27721 = ~n27730;
  assign n27050 = ~n25618;
  assign n27611 = ~n27620;
  assign n27674 = n27648 & n105;
  assign n27673 = ~n27648;
  assign n27680 = n27683 & n27684;
  assign n27656 = ~n27694;
  assign n27687 = n27640 & n27623;
  assign n27685 = ~n27640;
  assign n27692 = ~n27704;
  assign n26537 = ~n27717;
  assign n27705 = n27721 & n27722;
  assign n27662 = n27673 & n14279;
  assign n27630 = ~n27674;
  assign n27663 = ~n27680;
  assign n27681 = n27685 & n27686;
  assign n27642 = ~n27687;
  assign n27675 = n27692 & n27693;
  assign n26437 = n27705 ^ n27706;
  assign n27707 = ~n27705;
  assign n27645 = ~n27662;
  assign n27647 = n27663 & n27664;
  assign n27653 = n27675 ^ n27676;
  assign n27625 = ~n27681;
  assign n27678 = ~n27675;
  assign n24071 = n26437 ^ n25267;
  assign n27605 = n26437 ^ n26404;
  assign n27699 = n27707 & n27708;
  assign n27628 = n27647 ^ n27648;
  assign n27613 = n27653 ^ n27654;
  assign n27646 = ~n27647;
  assign n27665 = n27677 & n27678;
  assign n27666 = n24071 & n27679;
  assign n27669 = n27605 & n27586;
  assign n24129 = ~n24071;
  assign n27667 = ~n27605;
  assign n27688 = ~n27699;
  assign n27621 = n105 ^ n27628;
  assign n27637 = n27613 & n14245;
  assign n27644 = n27645 & n27646;
  assign n27638 = ~n27613;
  assign n27655 = ~n27665;
  assign n26461 = ~n27666;
  assign n27657 = n24129 & n26490;
  assign n27658 = n27667 & n27668;
  assign n27607 = ~n27669;
  assign n27670 = n27688 & n27689;
  assign n25543 = n27620 ^ n27621;
  assign n27610 = ~n27621;
  assign n27614 = ~n27637;
  assign n27631 = n27638 & n104;
  assign n27629 = ~n27644;
  assign n27639 = n27655 & n27656;
  assign n26492 = ~n27657;
  assign n27584 = ~n27658;
  assign n27649 = n27670 ^ n25293;
  assign n27671 = ~n27670;
  assign n26961 = ~n25543;
  assign n27578 = n27610 & n27611;
  assign n27612 = n27629 & n27630;
  assign n27591 = ~n27631;
  assign n27622 = n27639 ^ n27640;
  assign n27641 = ~n27639;
  assign n24080 = n27649 ^ n27650;
  assign n27659 = n27671 & n27672;
  assign n27601 = n27612 ^ n27613;
  assign n27561 = n27622 ^ n27623;
  assign n27615 = ~n27612;
  assign n26369 = n24080 ^ n25194;
  assign n27632 = n27641 & n27642;
  assign n27633 = n24080 & n27643;
  assign n24029 = ~n24080;
  assign n27651 = ~n27659;
  assign n27579 = n104 ^ n27601;
  assign n27602 = n27561 & n14200;
  assign n27609 = n27614 & n27615;
  assign n27603 = ~n27561;
  assign n27570 = n26369 ^ n26344;
  assign n27624 = ~n27632;
  assign n26408 = ~n27633;
  assign n27626 = n24029 & n26405;
  assign n27634 = n27651 & n27652;
  assign n25467 = n27578 ^ n27579;
  assign n27538 = n27579 & n27578;
  assign n27581 = ~n27602;
  assign n27592 = n27603 & n119;
  assign n27593 = n27570 & n27547;
  assign n27590 = ~n27609;
  assign n27594 = ~n27570;
  assign n27604 = n27624 & n27625;
  assign n26440 = ~n27626;
  assign n27617 = n27634 ^ n25178;
  assign n27635 = ~n27634;
  assign n27541 = ~n27538;
  assign n27580 = n27590 & n27591;
  assign n27563 = ~n27592;
  assign n27549 = ~n27593;
  assign n27587 = n27594 & n27595;
  assign n27585 = n27604 ^ n27605;
  assign n27606 = ~n27604;
  assign n24010 = n27616 ^ n27617;
  assign n27627 = n27635 & n27636;
  assign n27560 = n119 ^ n27580;
  assign n27543 = n27585 ^ n27586;
  assign n27582 = ~n27580;
  assign n27572 = ~n27587;
  assign n27596 = n27606 & n27607;
  assign n27597 = n24010 & n27608;
  assign n24037 = ~n24010;
  assign n27618 = ~n27627;
  assign n27539 = n27560 ^ n27561;
  assign n27567 = n27543 & n14171;
  assign n27573 = n27581 & n27582;
  assign n27568 = ~n27543;
  assign n26309 = n24037 ^ n25180;
  assign n27583 = ~n27596;
  assign n26375 = ~n27597;
  assign n27588 = n24037 & n26347;
  assign n27598 = n27618 & n27619;
  assign n24740 = n27538 ^ n27539;
  assign n27540 = ~n27539;
  assign n27545 = ~n27567;
  assign n27564 = n27568 & n118;
  assign n27506 = n26309 ^ n26239;
  assign n27562 = ~n27573;
  assign n27569 = n27583 & n27584;
  assign n26350 = ~n27588;
  assign n27574 = n27598 ^ n25129;
  assign n27599 = ~n27598;
  assign n27510 = ~n24740;
  assign n27494 = n27540 & n27541;
  assign n27542 = n27562 & n27563;
  assign n27519 = ~n27564;
  assign n27553 = n27506 & n27565;
  assign n27554 = ~n27506;
  assign n27546 = n27569 ^ n27570;
  assign n27571 = ~n27569;
  assign n24008 = n27574 ^ n27575;
  assign n27589 = n27599 & n27600;
  assign n26601 = n26604 ^ n27510;
  assign n27487 = n27510 ^ n27511;
  assign n27491 = n27510 & n24728;
  assign n27517 = n27542 ^ n27543;
  assign n27498 = n27546 ^ n27547;
  assign n27544 = ~n27542;
  assign n27508 = ~n27553;
  assign n27550 = n27554 & n27529;
  assign n26242 = n24008 ^ n25182;
  assign n27555 = n24008 & n26279;
  assign n27566 = n27571 & n27572;
  assign n23970 = ~n24008;
  assign n27576 = ~n27589;
  assign n23792 = n26601 ^ n26628;
  assign n25102 = n199 ^ n27487;
  assign n27361 = n26601 & n27490;
  assign n27264 = n27487 & n199;
  assign n27466 = n27491 ^ n24675;
  assign n27493 = n27491 & n24675;
  assign n27492 = ~n27491;
  assign n27495 = n118 ^ n27517;
  assign n27525 = n27498 & n14111;
  assign n27533 = n27544 & n27545;
  assign n27526 = ~n27498;
  assign n27458 = n26242 ^ n26227;
  assign n27530 = ~n27550;
  assign n26282 = ~n27555;
  assign n27551 = n23970 & n27556;
  assign n27548 = ~n27566;
  assign n27557 = n27576 & n27577;
  assign n25132 = ~n25102;
  assign n27488 = n27492 & n24715;
  assign n27445 = ~n27493;
  assign n27465 = n27494 ^ n27495;
  assign n27496 = ~n27495;
  assign n27500 = ~n27525;
  assign n27520 = n27526 & n117;
  assign n27522 = n27458 & n27527;
  assign n27518 = ~n27533;
  assign n27521 = ~n27458;
  assign n27528 = n27548 & n27549;
  assign n26312 = ~n27551;
  assign n27535 = n27557 ^ n25088;
  assign n27558 = ~n27557;
  assign n23638 = n27465 ^ n27466;
  assign n27467 = ~n27488;
  assign n27446 = n27496 & n27494;
  assign n27497 = n27518 & n27519;
  assign n27470 = ~n27520;
  assign n27512 = n27521 & n27484;
  assign n27460 = ~n27522;
  assign n27505 = n27528 ^ n27529;
  assign n23906 = n27534 ^ n27535;
  assign n27531 = ~n27528;
  assign n27552 = n27558 & n27559;
  assign n27433 = n27443 ^ n23638;
  assign n23621 = ~n23638;
  assign n27461 = n27467 & n27465;
  assign n27468 = n27497 ^ n27498;
  assign n27450 = n27505 ^ n27506;
  assign n27499 = ~n27497;
  assign n27486 = ~n27512;
  assign n26161 = n23906 ^ n25088;
  assign n27523 = n27530 & n27531;
  assign n27524 = n23906 & n27532;
  assign n23968 = ~n23906;
  assign n27536 = ~n27552;
  assign n27414 = n27433 & n27434;
  assign n27415 = ~n27433;
  assign n27444 = ~n27461;
  assign n27447 = n117 ^ n27468;
  assign n27482 = n27450 & n116;
  assign n27489 = n27499 & n27500;
  assign n27481 = ~n27450;
  assign n27405 = n26161 ^ n26099;
  assign n27507 = ~n27523;
  assign n26210 = ~n27524;
  assign n27513 = n23968 & n26244;
  assign n27514 = n27536 & n27537;
  assign n27363 = ~n27414;
  assign n27409 = n27415 & n27416;
  assign n27417 = n27444 & n27445;
  assign n27392 = n27446 ^ n27447;
  assign n27448 = ~n27447;
  assign n27471 = n27481 & n14072;
  assign n27422 = ~n27482;
  assign n27474 = n27405 & n27438;
  assign n27469 = ~n27489;
  assign n27472 = ~n27405;
  assign n27483 = n27507 & n27508;
  assign n26246 = ~n27513;
  assign n27501 = n27514 ^ n25100;
  assign n27515 = ~n27514;
  assign n27390 = ~n27409;
  assign n27391 = n27417 ^ n24666;
  assign n27419 = n27417 & n24666;
  assign n27418 = ~n27417;
  assign n27394 = n27448 & n27446;
  assign n27449 = n27469 & n27470;
  assign n27452 = ~n27471;
  assign n27462 = n27472 & n27473;
  assign n27407 = ~n27474;
  assign n27457 = n27483 ^ n27484;
  assign n27485 = ~n27483;
  assign n23937 = n27501 ^ n27502;
  assign n27509 = n27515 & n27516;
  assign n27387 = n27390 & n27361;
  assign n27360 = n27390 & n27363;
  assign n23564 = n27391 ^ n27392;
  assign n27410 = n27418 & n24670;
  assign n27403 = ~n27419;
  assign n27420 = n27449 ^ n27450;
  assign n27397 = n27457 ^ n27458;
  assign n27451 = ~n27449;
  assign n27440 = ~n27462;
  assign n26100 = n25056 ^ n23937;
  assign n27475 = n27485 & n27486;
  assign n27477 = n23937 & n26136;
  assign n23933 = ~n23937;
  assign n27503 = ~n27509;
  assign n27347 = n27360 ^ n27361;
  assign n27288 = n23564 ^ n27364;
  assign n27362 = ~n27387;
  assign n23550 = ~n23564;
  assign n27393 = n27403 & n27392;
  assign n27379 = ~n27410;
  assign n27395 = n116 ^ n27420;
  assign n27436 = n27397 & n115;
  assign n27442 = n27451 & n27452;
  assign n27435 = ~n27397;
  assign n27352 = n26100 ^ n26064;
  assign n27459 = ~n27475;
  assign n27463 = n23933 & n27476;
  assign n26139 = ~n27477;
  assign n27478 = n27503 & n27504;
  assign n27330 = n27347 & n198;
  assign n27331 = n27288 & n27325;
  assign n27329 = ~n27347;
  assign n27332 = ~n27288;
  assign n27356 = n27362 & n27363;
  assign n27378 = ~n27393;
  assign n27313 = n27394 ^ n27395;
  assign n27335 = n27395 & n27394;
  assign n27423 = n27435 & n14061;
  assign n27369 = ~n27436;
  assign n27424 = n27352 & n27384;
  assign n27421 = ~n27442;
  assign n27425 = ~n27352;
  assign n27437 = n27459 & n27460;
  assign n26176 = ~n27463;
  assign n27454 = n27478 ^ n25012;
  assign n27479 = ~n27478;
  assign n27324 = n27329 & n8617;
  assign n27266 = ~n27330;
  assign n27268 = ~n27331;
  assign n27326 = n27332 & n27333;
  assign n27297 = ~n27356;
  assign n27348 = n27378 & n27379;
  assign n27365 = n27313 & n24630;
  assign n27366 = ~n27313;
  assign n27338 = ~n27335;
  assign n27396 = n27421 & n27422;
  assign n27398 = ~n27423;
  assign n27354 = ~n27424;
  assign n27411 = n27425 & n27426;
  assign n27404 = n27437 ^ n27438;
  assign n27439 = ~n27437;
  assign n23909 = n27453 ^ n27454;
  assign n27464 = n27479 & n27480;
  assign n27295 = ~n27324;
  assign n27287 = n27297 ^ n27325;
  assign n27296 = ~n27326;
  assign n27314 = n27348 ^ n24620;
  assign n27350 = ~n27348;
  assign n27349 = ~n27365;
  assign n27357 = n27366 & n24620;
  assign n27367 = n27396 ^ n27397;
  assign n27340 = n27404 ^ n27405;
  assign n27399 = ~n27396;
  assign n27386 = ~n27411;
  assign n26026 = n25049 ^ n23909;
  assign n27427 = n27439 & n27440;
  assign n27428 = n23909 & n27441;
  assign n23850 = ~n23909;
  assign n27455 = ~n27464;
  assign n27220 = n27287 ^ n27288;
  assign n27289 = n27295 & n27264;
  assign n27263 = n27295 & n27266;
  assign n27290 = n27296 & n27297;
  assign n23520 = n27313 ^ n27314;
  assign n27334 = n27349 & n27350;
  assign n27316 = ~n27357;
  assign n27336 = n115 ^ n27367;
  assign n27380 = n27340 & n14006;
  assign n27388 = n27398 & n27399;
  assign n27381 = ~n27340;
  assign n27284 = n26026 ^ n25941;
  assign n27406 = ~n27427;
  assign n26068 = ~n27428;
  assign n27412 = n23850 & n26065;
  assign n27429 = n27455 & n27456;
  assign n27258 = n27220 & n197;
  assign n27226 = n27263 ^ n27264;
  assign n27257 = ~n27220;
  assign n27191 = n27281 ^ n23520;
  assign n27265 = ~n27289;
  assign n27267 = ~n27290;
  assign n23516 = ~n23520;
  assign n27315 = ~n27334;
  assign n27249 = n27335 ^ n27336;
  assign n27337 = ~n27336;
  assign n27342 = ~n27380;
  assign n27370 = n27381 & n114;
  assign n27372 = n27284 & n27382;
  assign n27368 = ~n27388;
  assign n27371 = ~n27284;
  assign n27383 = n27406 & n27407;
  assign n26103 = ~n27412;
  assign n23788 = n27429 ^ n27430;
  assign n27431 = ~n27429;
  assign n25953 = n27226 ^ n25102;
  assign n27153 = n27226 & n25102;
  assign n27244 = n27257 & n8554;
  assign n27189 = ~n27258;
  assign n27247 = n27191 & n27221;
  assign n27259 = n27265 & n27266;
  assign n27260 = n27267 & n27268;
  assign n27245 = ~n27191;
  assign n27282 = n27315 & n27316;
  assign n27299 = n27249 & n24591;
  assign n27298 = ~n27249;
  assign n27271 = n27337 & n27338;
  assign n27339 = n27368 & n27369;
  assign n27302 = ~n27370;
  assign n27358 = n27371 & n27320;
  assign n27286 = ~n27372;
  assign n27351 = n27383 ^ n27384;
  assign n27385 = ~n27383;
  assign n25951 = n24958 ^ n23788;
  assign n27400 = n23788 & n27408;
  assign n23848 = ~n23788;
  assign n27413 = n27431 & n27432;
  assign n25967 = ~n25953;
  assign n27156 = ~n27153;
  assign n27218 = ~n27244;
  assign n27227 = n27245 & n27246;
  assign n27177 = ~n27247;
  assign n27219 = ~n27259;
  assign n27212 = ~n27260;
  assign n27248 = n27282 ^ n24588;
  assign n27269 = ~n27282;
  assign n27291 = n27298 & n24588;
  assign n27229 = ~n27299;
  assign n27274 = ~n27271;
  assign n27300 = n27339 ^ n27340;
  assign n27276 = n27351 ^ n27352;
  assign n27341 = ~n27339;
  assign n27322 = ~n27358;
  assign n27254 = n25951 ^ n25929;
  assign n27373 = n27385 & n27386;
  assign n27389 = n23848 & n25992;
  assign n25994 = ~n27400;
  assign n27401 = ~n27413;
  assign n27210 = n27218 & n27219;
  assign n27187 = n27219 ^ n27220;
  assign n27190 = n27212 ^ n27221;
  assign n27211 = ~n27227;
  assign n23415 = n27248 ^ n27249;
  assign n27270 = ~n27291;
  assign n27272 = n114 ^ n27300;
  assign n27317 = n27276 & n13964;
  assign n27327 = n27341 & n27342;
  assign n27318 = ~n27276;
  assign n27344 = n27254 & n27355;
  assign n27343 = ~n27254;
  assign n27353 = ~n27373;
  assign n26029 = ~n27389;
  assign n27374 = n27401 & n27402;
  assign n27154 = n197 ^ n27187;
  assign n27143 = n27190 ^ n27191;
  assign n27188 = ~n27210;
  assign n27195 = n27211 & n27212;
  assign n27111 = n27213 ^ n23415;
  assign n23449 = ~n23415;
  assign n27261 = n27269 & n27270;
  assign n27250 = n27271 ^ n27272;
  assign n27273 = ~n27272;
  assign n27278 = ~n27317;
  assign n27303 = n27318 & n113;
  assign n27301 = ~n27327;
  assign n27328 = n27343 & n27215;
  assign n27256 = ~n27344;
  assign n27319 = n27353 & n27354;
  assign n25871 = n27374 ^ n27375;
  assign n27376 = ~n27374;
  assign n25060 = n27153 ^ n27154;
  assign n27158 = n27143 & n196;
  assign n27155 = ~n27154;
  assign n27157 = ~n27143;
  assign n27175 = n27188 & n27189;
  assign n27179 = n27111 & n27192;
  assign n27176 = ~n27195;
  assign n27178 = ~n27111;
  assign n27230 = n27250 & n24566;
  assign n27228 = ~n27261;
  assign n27163 = ~n27250;
  assign n27199 = n27273 & n27274;
  assign n27275 = n27301 & n27302;
  assign n27233 = ~n27303;
  assign n27283 = n27319 ^ n27320;
  assign n27217 = ~n27328;
  assign n27321 = ~n27319;
  assign n27183 = n25871 ^ n25833;
  assign n23809 = n25871 ^ n24924;
  assign n27359 = n27376 & n27377;
  assign n25891 = ~n25060;
  assign n27069 = n27155 & n27156;
  assign n27144 = n27157 & n8495;
  assign n27084 = ~n27158;
  assign n27126 = ~n27175;
  assign n27145 = n27176 & n27177;
  assign n27161 = n27178 & n27146;
  assign n27114 = ~n27179;
  assign n27196 = n27228 & n27229;
  assign n27222 = n27163 & n24536;
  assign n27198 = ~n27230;
  assign n27231 = n27275 ^ n27276;
  assign n27203 = n27283 ^ n27284;
  assign n27277 = ~n27275;
  assign n27304 = n27321 & n27322;
  assign n27305 = n27183 & n27150;
  assign n27308 = n23809 & n27323;
  assign n27306 = ~n27183;
  assign n23796 = ~n23809;
  assign n27345 = ~n27359;
  assign n27082 = ~n27069;
  assign n27109 = n27126 ^ n27143;
  assign n27125 = ~n27144;
  assign n27110 = n27145 ^ n27146;
  assign n27148 = ~n27145;
  assign n27147 = ~n27161;
  assign n27162 = n27196 ^ n24566;
  assign n27197 = ~n27196;
  assign n27165 = ~n27222;
  assign n27200 = n113 ^ n27231;
  assign n27252 = n27203 & n112;
  assign n27262 = n27277 & n27278;
  assign n27251 = ~n27203;
  assign n27285 = ~n27304;
  assign n27152 = ~n27305;
  assign n27292 = n27306 & n27307;
  assign n25918 = ~n27308;
  assign n27293 = n23796 & n25955;
  assign n27309 = n27345 & n27346;
  assign n27070 = n196 ^ n27109;
  assign n27039 = n27110 ^ n27111;
  assign n27112 = n27125 & n27126;
  assign n27129 = n27147 & n27148;
  assign n23409 = n27162 ^ n27163;
  assign n27193 = n27197 & n27198;
  assign n27093 = n27199 ^ n27200;
  assign n27201 = ~n27200;
  assign n27234 = n27251 & n13918;
  assign n27168 = ~n27252;
  assign n27232 = ~n27262;
  assign n27253 = n27285 & n27286;
  assign n27185 = ~n27292;
  assign n25957 = ~n27293;
  assign n25804 = n27309 ^ n27310;
  assign n27311 = ~n27309;
  assign n25018 = n27069 ^ n27070;
  assign n26963 = n27070 & n27082;
  assign n27072 = n27039 & n195;
  assign n27071 = ~n27039;
  assign n27083 = ~n27112;
  assign n27113 = ~n27129;
  assign n27038 = n27130 ^ n23409;
  assign n23368 = ~n23409;
  assign n27164 = ~n27193;
  assign n27134 = n27201 & n27199;
  assign n27202 = n27232 & n27233;
  assign n27204 = ~n27234;
  assign n27214 = n27253 ^ n27254;
  assign n27255 = ~n27253;
  assign n27121 = n25804 ^ n25675;
  assign n23743 = n25804 ^ n24882;
  assign n27294 = n27311 & n27312;
  assign n25805 = ~n25018;
  assign n27053 = n27071 & n8474;
  assign n26999 = ~n27072;
  assign n27073 = n27083 & n27084;
  assign n27074 = n27113 & n27114;
  assign n27090 = n27038 & n27115;
  assign n27091 = ~n27038;
  assign n27131 = n27164 & n27165;
  assign n27166 = n27202 ^ n27203;
  assign n27098 = n27214 ^ n27215;
  assign n27205 = ~n27202;
  assign n27235 = n27255 & n27256;
  assign n27238 = n27121 & n27079;
  assign n27239 = n23743 & n25842;
  assign n27236 = ~n27121;
  assign n23759 = ~n23743;
  assign n27279 = ~n27294;
  assign n27035 = ~n27053;
  assign n27036 = ~n27073;
  assign n27037 = n27074 ^ n27075;
  assign n27054 = ~n27074;
  assign n27017 = ~n27090;
  assign n27085 = n27091 & n27075;
  assign n27092 = n27131 ^ n24509;
  assign n27133 = n27131 & n24509;
  assign n27132 = ~n27131;
  assign n27135 = n112 ^ n27166;
  assign n27181 = n27098 & n127;
  assign n27194 = n27204 & n27205;
  assign n27180 = ~n27098;
  assign n27216 = ~n27235;
  assign n27223 = n27236 & n27237;
  assign n27123 = ~n27238;
  assign n25881 = ~n27239;
  assign n27224 = n23759 & n27240;
  assign n27241 = n27279 & n27280;
  assign n27015 = n27035 & n27036;
  assign n26966 = n27037 ^ n27038;
  assign n26997 = n27036 ^ n27039;
  assign n27055 = ~n27085;
  assign n23353 = n27092 ^ n27093;
  assign n27127 = n27132 & n24540;
  assign n27116 = ~n27133;
  assign n27002 = n27134 ^ n27135;
  assign n27057 = n27135 & n27134;
  assign n27169 = n27180 & n13893;
  assign n27100 = ~n27181;
  assign n27167 = ~n27194;
  assign n27182 = n27216 & n27217;
  assign n27081 = ~n27223;
  assign n25845 = ~n27224;
  assign n27207 = n27241 ^ n24865;
  assign n27242 = ~n27241;
  assign n26964 = n195 ^ n26997;
  assign n27001 = n26966 & n194;
  assign n26998 = ~n27015;
  assign n27000 = ~n26966;
  assign n27051 = n27054 & n27055;
  assign n26947 = n27056 ^ n23353;
  assign n23348 = ~n23353;
  assign n27094 = n27116 & n27093;
  assign n27096 = n27002 & n24479;
  assign n27077 = ~n27127;
  assign n27095 = ~n27002;
  assign n27060 = ~n27057;
  assign n27136 = n27167 & n27168;
  assign n27138 = ~n27169;
  assign n27149 = n27182 ^ n27183;
  assign n27184 = ~n27182;
  assign n23734 = n27206 ^ n27207;
  assign n27225 = n27242 & n27243;
  assign n24961 = n26963 ^ n26964;
  assign n26893 = n26964 & n26963;
  assign n26965 = n26998 & n26999;
  assign n26982 = n27000 & n8425;
  assign n26929 = ~n27001;
  assign n27018 = n26947 & n27040;
  assign n27016 = ~n27051;
  assign n27019 = ~n26947;
  assign n27076 = ~n27094;
  assign n27086 = n27095 & n24507;
  assign n27043 = ~n27096;
  assign n27097 = n127 ^ n27136;
  assign n27062 = n27149 ^ n27150;
  assign n27137 = ~n27136;
  assign n25729 = n23734 ^ n24865;
  assign n27170 = n27184 & n27185;
  assign n27171 = n23734 & n27186;
  assign n23656 = ~n23734;
  assign n27208 = ~n27225;
  assign n25743 = ~n24961;
  assign n26927 = n26965 ^ n26966;
  assign n26968 = ~n26965;
  assign n26967 = ~n26982;
  assign n26983 = n27016 & n27017;
  assign n26949 = ~n27018;
  assign n27010 = n27019 & n26984;
  assign n27041 = n27076 & n27077;
  assign n27005 = ~n27086;
  assign n27058 = n27097 ^ n27098;
  assign n27117 = n27062 & n13832;
  assign n27128 = n27137 & n27138;
  assign n27118 = ~n27062;
  assign n27007 = n25729 ^ n25692;
  assign n27151 = ~n27170;
  assign n25773 = ~n27171;
  assign n27159 = n23656 & n25808;
  assign n27172 = n27208 & n27209;
  assign n26894 = n194 ^ n26927;
  assign n26945 = n26967 & n26968;
  assign n26946 = n26983 ^ n26984;
  assign n26985 = ~n26983;
  assign n26986 = ~n27010;
  assign n27003 = n27041 ^ n24507;
  assign n27042 = ~n27041;
  assign n26933 = n27057 ^ n27058;
  assign n27059 = ~n27058;
  assign n27064 = ~n27117;
  assign n27101 = n27118 & n126;
  assign n27102 = n27007 & n27119;
  assign n27099 = ~n27128;
  assign n27103 = ~n27007;
  assign n27120 = n27151 & n27152;
  assign n25810 = ~n27159;
  assign n27139 = n27172 ^ n24828;
  assign n27173 = ~n27172;
  assign n24945 = n26893 ^ n26894;
  assign n26895 = ~n26894;
  assign n26928 = ~n26945;
  assign n26897 = n26946 ^ n26947;
  assign n26980 = n26985 & n26986;
  assign n23268 = n27002 ^ n27003;
  assign n27020 = n27042 & n27043;
  assign n27022 = n26933 & n24470;
  assign n27021 = ~n26933;
  assign n26987 = n27059 & n27060;
  assign n27061 = n27099 & n27100;
  assign n27025 = ~n27101;
  assign n27009 = ~n27102;
  assign n27087 = n27103 & n27047;
  assign n27078 = n27120 ^ n27121;
  assign n27122 = ~n27120;
  assign n23670 = n27139 ^ n27140;
  assign n27160 = n27173 & n27174;
  assign n25664 = ~n24945;
  assign n26827 = n26895 & n26893;
  assign n26896 = n26928 & n26929;
  assign n26915 = n26897 & n193;
  assign n26914 = ~n26897;
  assign n26876 = n26969 ^ n23268;
  assign n26948 = ~n26980;
  assign n23319 = ~n23268;
  assign n27004 = ~n27020;
  assign n27011 = n27021 & n24444;
  assign n26936 = ~n27022;
  assign n27023 = n27061 ^ n27062;
  assign n26990 = n27078 ^ n27079;
  assign n27063 = ~n27061;
  assign n27049 = ~n27087;
  assign n25653 = n24916 ^ n23670;
  assign n27104 = n27122 & n27123;
  assign n27105 = n23670 & n27124;
  assign n23686 = ~n23670;
  assign n27141 = ~n27160;
  assign n26861 = n26896 ^ n26897;
  assign n26881 = ~n26896;
  assign n26911 = n26914 & n8392;
  assign n26849 = ~n26915;
  assign n26930 = n26876 & n26912;
  assign n26941 = n26948 & n26949;
  assign n26931 = ~n26876;
  assign n26970 = n27004 & n27005;
  assign n26972 = ~n27011;
  assign n26988 = n126 ^ n27023;
  assign n27044 = n26990 & n13776;
  assign n27052 = n27063 & n27064;
  assign n27045 = ~n26990;
  assign n26938 = n25653 ^ n25564;
  assign n27080 = ~n27104;
  assign n27088 = n23686 & n25694;
  assign n25733 = ~n27105;
  assign n27106 = n27141 & n27142;
  assign n26828 = n193 ^ n26861;
  assign n26880 = ~n26911;
  assign n26863 = ~n26930;
  assign n26916 = n26931 & n26932;
  assign n26899 = ~n26941;
  assign n26934 = n26970 ^ n24444;
  assign n26971 = ~n26970;
  assign n26867 = n26987 ^ n26988;
  assign n26917 = n26988 & n26987;
  assign n26992 = ~n27044;
  assign n27026 = n27045 & n125;
  assign n27027 = n26938 & n26977;
  assign n27024 = ~n27052;
  assign n27028 = ~n26938;
  assign n27046 = n27080 & n27081;
  assign n25697 = ~n27088;
  assign n27065 = n27106 ^ n24795;
  assign n27107 = ~n27106;
  assign n24886 = n26827 ^ n26828;
  assign n26829 = ~n26828;
  assign n26874 = n26880 & n26881;
  assign n26875 = n26899 ^ n26912;
  assign n26898 = ~n26916;
  assign n23230 = n26933 ^ n26934;
  assign n26950 = n26971 & n26972;
  assign n26952 = n26867 & n24442;
  assign n26951 = ~n26867;
  assign n26920 = ~n26917;
  assign n26989 = n27024 & n27025;
  assign n26955 = ~n27026;
  assign n26940 = ~n27027;
  assign n27012 = n27028 & n27029;
  assign n27006 = n27046 ^ n27047;
  assign n27048 = ~n27046;
  assign n23582 = n27065 ^ n27066;
  assign n27089 = n27107 & n27108;
  assign n25591 = ~n24886;
  assign n26757 = n26829 & n26827;
  assign n26848 = ~n26874;
  assign n26816 = n26875 ^ n26876;
  assign n26882 = n26898 & n26899;
  assign n26797 = n26900 ^ n23230;
  assign n23275 = ~n23230;
  assign n26935 = ~n26950;
  assign n26942 = n26951 & n24410;
  assign n26869 = ~n26952;
  assign n26953 = n26989 ^ n26990;
  assign n26922 = n27006 ^ n27007;
  assign n26991 = ~n26989;
  assign n26979 = ~n27012;
  assign n25583 = n24831 ^ n23582;
  assign n27030 = n27048 & n27049;
  assign n27031 = n23582 & n27050;
  assign n23541 = ~n23582;
  assign n27067 = ~n27089;
  assign n26815 = n26848 & n26849;
  assign n26846 = n26816 & n192;
  assign n26845 = ~n26816;
  assign n26864 = n26797 & n26877;
  assign n26862 = ~n26882;
  assign n26865 = ~n26797;
  assign n26901 = n26935 & n26936;
  assign n26903 = ~n26942;
  assign n26918 = n125 ^ n26953;
  assign n26974 = n26922 & n124;
  assign n26981 = n26991 & n26992;
  assign n26973 = ~n26922;
  assign n26871 = n25583 ^ n25490;
  assign n27008 = ~n27030;
  assign n25621 = ~n27031;
  assign n27013 = n23541 & n25618;
  assign n27032 = n27067 & n27068;
  assign n26786 = n26815 ^ n26816;
  assign n26811 = ~n26815;
  assign n26830 = n26845 & n8358;
  assign n26784 = ~n26846;
  assign n26831 = n26862 & n26863;
  assign n26800 = ~n26864;
  assign n26850 = n26865 & n26832;
  assign n26866 = n26901 ^ n24410;
  assign n26902 = ~n26901;
  assign n26804 = n26917 ^ n26918;
  assign n26919 = ~n26918;
  assign n26956 = n26973 & n13745;
  assign n26888 = ~n26974;
  assign n26957 = n26871 & n26975;
  assign n26954 = ~n26981;
  assign n26958 = ~n26871;
  assign n26976 = n27008 & n27009;
  assign n25657 = ~n27013;
  assign n26994 = n27032 ^ n24766;
  assign n27033 = ~n27032;
  assign n26758 = n192 ^ n26786;
  assign n26812 = ~n26830;
  assign n26796 = n26831 ^ n26832;
  assign n26833 = ~n26831;
  assign n26834 = ~n26850;
  assign n23237 = n26866 ^ n26867;
  assign n26883 = n26902 & n26903;
  assign n26885 = n26804 & n24372;
  assign n26884 = ~n26804;
  assign n26851 = n26919 & n26920;
  assign n26921 = n26954 & n26955;
  assign n26924 = ~n26956;
  assign n26873 = ~n26957;
  assign n26943 = n26958 & n26908;
  assign n26937 = n26976 ^ n26977;
  assign n26978 = ~n26976;
  assign n23485 = n26993 ^ n26994;
  assign n27014 = n27033 & n27034;
  assign n24869 = n26757 ^ n26758;
  assign n26759 = ~n26758;
  assign n26744 = n26796 ^ n26797;
  assign n26798 = n26811 & n26812;
  assign n26817 = n26833 & n26834;
  assign n26743 = n26835 ^ n23237;
  assign n23217 = ~n23237;
  assign n26868 = ~n26883;
  assign n26878 = n26884 & n24408;
  assign n26838 = ~n26885;
  assign n26854 = ~n26851;
  assign n26886 = n26921 ^ n26922;
  assign n26856 = n26937 ^ n26938;
  assign n26923 = ~n26921;
  assign n26910 = ~n26943;
  assign n25505 = n23485 ^ n24766;
  assign n26959 = n26978 & n26979;
  assign n26960 = n23485 & n25543;
  assign n23556 = ~n23485;
  assign n26995 = ~n27014;
  assign n25513 = ~n24869;
  assign n25437 = n26759 & n26757;
  assign n26770 = n26744 & n207;
  assign n26769 = ~n26744;
  assign n26783 = ~n26798;
  assign n26802 = n26743 & n26813;
  assign n26799 = ~n26817;
  assign n26801 = ~n26743;
  assign n26836 = n26868 & n26869;
  assign n26806 = ~n26878;
  assign n26852 = n124 ^ n26886;
  assign n26904 = n26856 & n13696;
  assign n26913 = n26923 & n26924;
  assign n26905 = ~n26856;
  assign n26808 = n25505 ^ n25420;
  assign n26939 = ~n26959;
  assign n25545 = ~n26960;
  assign n26944 = n23556 & n26961;
  assign n26962 = n26995 & n26996;
  assign n26690 = ~n25437;
  assign n26760 = n26769 & n8317;
  assign n26718 = ~n26770;
  assign n26771 = n26783 & n26784;
  assign n26772 = n26799 & n26800;
  assign n26787 = n26801 & n26773;
  assign n26746 = ~n26802;
  assign n26803 = n26836 ^ n24408;
  assign n26837 = ~n26836;
  assign n26751 = n26851 ^ n26852;
  assign n26853 = ~n26852;
  assign n26858 = ~n26904;
  assign n26889 = n26905 & n123;
  assign n26891 = n26808 & n26906;
  assign n26887 = ~n26913;
  assign n26890 = ~n26808;
  assign n26907 = n26939 & n26940;
  assign n25587 = ~n26944;
  assign n26926 = n26962 ^ n24783;
  assign n26740 = ~n26760;
  assign n26741 = ~n26771;
  assign n26742 = n26772 ^ n26773;
  assign n26774 = ~n26772;
  assign n26775 = ~n26787;
  assign n23249 = n26803 ^ n26804;
  assign n26818 = n26837 & n26838;
  assign n26819 = n26751 & n24333;
  assign n26820 = ~n26751;
  assign n26788 = n26853 & n26854;
  assign n26855 = n26887 & n26888;
  assign n26823 = ~n26889;
  assign n26879 = n26890 & n26842;
  assign n26810 = ~n26891;
  assign n26870 = n26907 ^ n26908;
  assign n26909 = ~n26907;
  assign n24799 = n26925 ^ n26926;
  assign n26730 = n26740 & n26741;
  assign n26692 = n26742 ^ n26743;
  assign n26716 = n26741 ^ n26744;
  assign n26761 = n26774 & n26775;
  assign n26696 = n26776 ^ n23249;
  assign n23183 = ~n23249;
  assign n26805 = ~n26818;
  assign n26753 = ~n26819;
  assign n26814 = n26820 & n24359;
  assign n26791 = ~n26788;
  assign n26821 = n26855 ^ n26856;
  assign n26793 = n26870 ^ n26871;
  assign n26857 = ~n26855;
  assign n26844 = ~n26879;
  assign n26859 = n24799 ^ n24783;
  assign n26892 = n26909 & n26910;
  assign n25396 = n207 ^ n26716;
  assign n26720 = n26692 & n206;
  assign n26717 = ~n26730;
  assign n26719 = ~n26692;
  assign n26749 = n26696 & n26722;
  assign n26745 = ~n26761;
  assign n26747 = ~n26696;
  assign n26777 = n26805 & n26806;
  assign n26779 = ~n26814;
  assign n26789 = n123 ^ n26821;
  assign n26840 = n26793 & n122;
  assign n26847 = n26857 & n26858;
  assign n26839 = ~n26793;
  assign n25436 = n26859 ^ n26860;
  assign n26872 = ~n26892;
  assign n26689 = ~n25396;
  assign n26691 = n26717 & n26718;
  assign n26708 = n26719 & n8278;
  assign n26672 = ~n26720;
  assign n26721 = n26745 & n26746;
  assign n26731 = n26747 & n26748;
  assign n26724 = ~n26749;
  assign n26750 = n26777 ^ n24359;
  assign n26778 = ~n26777;
  assign n26701 = n26788 ^ n26789;
  assign n26790 = ~n26789;
  assign n26755 = n25436 ^ n26825;
  assign n26824 = n26839 & n13622;
  assign n26767 = ~n26840;
  assign n26822 = ~n26847;
  assign n26841 = n26872 & n26873;
  assign n26646 = n26689 & n26690;
  assign n26670 = n26691 ^ n26692;
  assign n26694 = ~n26691;
  assign n26693 = ~n26708;
  assign n26695 = n26721 ^ n26722;
  assign n26723 = ~n26721;
  assign n26698 = ~n26731;
  assign n23211 = n26750 ^ n26751;
  assign n26762 = n26778 & n26779;
  assign n26764 = n26701 & n24293;
  assign n26763 = ~n26701;
  assign n26732 = n26790 & n26791;
  assign n26792 = n26822 & n26823;
  assign n26795 = ~n26824;
  assign n26807 = n26841 ^ n26842;
  assign n26843 = ~n26841;
  assign n26647 = n206 ^ n26670;
  assign n26649 = ~n26646;
  assign n26685 = n26693 & n26694;
  assign n26651 = n26695 ^ n26696;
  assign n26709 = n26723 & n26724;
  assign n26655 = n26725 ^ n23211;
  assign n23151 = ~n23211;
  assign n26752 = ~n26762;
  assign n26756 = n26763 & n24331;
  assign n26728 = ~n26764;
  assign n26735 = ~n26732;
  assign n26765 = n26792 ^ n26793;
  assign n26737 = n26807 ^ n26808;
  assign n26794 = ~n26792;
  assign n26826 = n26843 & n26844;
  assign n23802 = n26646 ^ n26647;
  assign n26648 = ~n26647;
  assign n26673 = n26651 & n8239;
  assign n26671 = ~n26685;
  assign n26674 = ~n26651;
  assign n26700 = n26655 & n26706;
  assign n26697 = ~n26709;
  assign n26699 = ~n26655;
  assign n26726 = n26752 & n26753;
  assign n26704 = ~n26756;
  assign n26733 = n122 ^ n26765;
  assign n26781 = n26737 & n121;
  assign n26785 = n26794 & n26795;
  assign n26780 = ~n26737;
  assign n26809 = ~n26826;
  assign n26602 = n23802 ^ n26628;
  assign n26542 = n23802 & n23792;
  assign n26605 = n26648 & n26649;
  assign n26650 = n26671 & n26672;
  assign n26653 = ~n26673;
  assign n26667 = n26674 & n205;
  assign n26675 = n26697 & n26698;
  assign n26686 = n26699 & n26676;
  assign n26657 = ~n26700;
  assign n26702 = n26726 ^ n24331;
  assign n26727 = ~n26726;
  assign n26661 = n26732 ^ n26733;
  assign n26734 = ~n26733;
  assign n26768 = n26780 & n13583;
  assign n26715 = ~n26781;
  assign n26766 = ~n26785;
  assign n26782 = n26809 & n26810;
  assign n22814 = n26601 ^ n26602;
  assign n24615 = n295 ^ n26602;
  assign n26332 = n26602 & n295;
  assign n26603 = ~n26602;
  assign n26608 = ~n26605;
  assign n26629 = n26650 ^ n26651;
  assign n26652 = ~n26650;
  assign n26631 = ~n26667;
  assign n26654 = n26675 ^ n26676;
  assign n26677 = ~n26675;
  assign n26678 = ~n26686;
  assign n23146 = n26701 ^ n26702;
  assign n26710 = n26727 & n26728;
  assign n26711 = n26661 & n24291;
  assign n26712 = ~n26661;
  assign n26687 = n26734 & n26735;
  assign n26736 = n26766 & n26767;
  assign n26739 = ~n26768;
  assign n26754 = n120 ^ n26782;
  assign n24636 = ~n24615;
  assign n26418 = n26603 & n26604;
  assign n26606 = n205 ^ n26629;
  assign n26644 = n26652 & n26653;
  assign n26610 = n26654 ^ n26655;
  assign n26668 = n26677 & n26678;
  assign n26614 = n26679 ^ n23146;
  assign n23114 = ~n23146;
  assign n26703 = ~n26710;
  assign n26665 = ~n26711;
  assign n26707 = n26712 & n24251;
  assign n26705 = ~n26687;
  assign n26713 = n26736 ^ n26737;
  assign n26663 = n26754 ^ n26755;
  assign n26738 = ~n26736;
  assign n26596 = n26605 ^ n26606;
  assign n26607 = ~n26606;
  assign n26633 = n26610 & n204;
  assign n26630 = ~n26644;
  assign n26632 = ~n26610;
  assign n26658 = n26614 & n26666;
  assign n26656 = ~n26668;
  assign n26659 = ~n26614;
  assign n26680 = n26703 & n26704;
  assign n26682 = ~n26707;
  assign n26688 = n121 ^ n26713;
  assign n26729 = n26738 & n26739;
  assign n26584 = n26596 & n23621;
  assign n26585 = ~n26596;
  assign n26564 = n26607 & n26608;
  assign n26609 = n26630 & n26631;
  assign n26624 = n26632 & n8227;
  assign n26588 = ~n26633;
  assign n26634 = n26656 & n26657;
  assign n26616 = ~n26658;
  assign n26645 = n26659 & n26635;
  assign n26660 = n26680 ^ n24251;
  assign n26681 = ~n26680;
  assign n26619 = n26687 ^ n26688;
  assign n26684 = n26688 & n26705;
  assign n26714 = ~n26729;
  assign n26563 = ~n26584;
  assign n26581 = n26585 & n23638;
  assign n26586 = n26609 ^ n26610;
  assign n26612 = ~n26609;
  assign n26611 = ~n26624;
  assign n26613 = n26634 ^ n26635;
  assign n26636 = ~n26634;
  assign n26637 = ~n26645;
  assign n23128 = n26660 ^ n26661;
  assign n26669 = n26681 & n26682;
  assign n26683 = n26714 & n26715;
  assign n26562 = n26563 & n26542;
  assign n26554 = ~n26581;
  assign n26565 = n204 ^ n26586;
  assign n26599 = n26611 & n26612;
  assign n26567 = n26613 ^ n26614;
  assign n26625 = n26636 & n26637;
  assign n26571 = n26638 ^ n23128;
  assign n23076 = ~n23128;
  assign n26664 = ~n26669;
  assign n26662 = n26683 ^ n26684;
  assign n26553 = ~n26562;
  assign n26541 = n26563 & n26554;
  assign n26555 = n26564 ^ n26565;
  assign n26519 = n26565 & n26564;
  assign n26590 = n26567 & n203;
  assign n26587 = ~n26599;
  assign n26589 = ~n26567;
  assign n26618 = n26571 & n26622;
  assign n26615 = ~n26625;
  assign n26617 = ~n26571;
  assign n26556 = n26662 ^ n26663;
  assign n26641 = n26664 & n26665;
  assign n22698 = n26541 ^ n26542;
  assign n26530 = n26553 & n26554;
  assign n26543 = n26555 & n23550;
  assign n26507 = ~n26555;
  assign n26566 = n26587 & n26588;
  assign n26582 = n26589 & n8167;
  assign n26546 = ~n26590;
  assign n26591 = n26615 & n26616;
  assign n26600 = n26617 & n26592;
  assign n26573 = ~n26618;
  assign n26620 = n26641 ^ n24239;
  assign n26639 = n26556 & n24198;
  assign n26643 = n26641 & n24239;
  assign n26640 = ~n26556;
  assign n26642 = ~n26641;
  assign n24694 = n22698 ^ n23638;
  assign n26506 = n26530 ^ n23550;
  assign n22689 = ~n22698;
  assign n26532 = ~n26530;
  assign n26538 = n26507 & n23564;
  assign n26531 = ~n26543;
  assign n26544 = n26566 ^ n26567;
  assign n26568 = ~n26566;
  assign n26569 = ~n26582;
  assign n26570 = n26591 ^ n26592;
  assign n26593 = ~n26591;
  assign n26594 = ~n26600;
  assign n23095 = n26619 ^ n26620;
  assign n26559 = ~n26639;
  assign n26626 = n26640 & n24171;
  assign n26627 = n26642 & n24211;
  assign n26623 = ~n26643;
  assign n26482 = n24694 ^ n24675;
  assign n22589 = n26506 ^ n26507;
  assign n26518 = n26531 & n26532;
  assign n26509 = ~n26538;
  assign n26520 = n203 ^ n26544;
  assign n26560 = n26568 & n26569;
  assign n26522 = n26570 ^ n26571;
  assign n26583 = n26593 & n26594;
  assign n26526 = n26595 ^ n23095;
  assign n23082 = ~n23095;
  assign n26621 = n26623 & n26619;
  assign n26580 = ~n26626;
  assign n26598 = ~n26627;
  assign n26471 = n26482 & n26483;
  assign n24676 = n23564 ^ n22589;
  assign n26469 = ~n26482;
  assign n22628 = ~n22589;
  assign n26508 = ~n26518;
  assign n26453 = n26519 ^ n26520;
  assign n26473 = n26520 & n26519;
  assign n26548 = n26522 & n202;
  assign n26545 = ~n26560;
  assign n26547 = ~n26522;
  assign n26574 = n26526 & n26550;
  assign n26572 = ~n26583;
  assign n26575 = ~n26526;
  assign n26597 = ~n26621;
  assign n26352 = n24676 ^ n24670;
  assign n26462 = n26469 & n26470;
  assign n26420 = ~n26471;
  assign n26484 = n26508 & n26509;
  assign n26499 = n26453 & n23516;
  assign n26498 = ~n26453;
  assign n26476 = ~n26473;
  assign n26521 = n26545 & n26546;
  assign n26539 = n26547 & n8128;
  assign n26502 = ~n26548;
  assign n26549 = n26572 & n26573;
  assign n26552 = ~n26574;
  assign n26561 = n26575 & n26576;
  assign n26578 = n26597 & n26598;
  assign n26431 = n26352 & n26379;
  assign n26429 = ~n26352;
  assign n26448 = ~n26462;
  assign n26454 = n26484 ^ n23520;
  assign n26486 = ~n26484;
  assign n26493 = n26498 & n23520;
  assign n26485 = ~n26499;
  assign n26500 = n26521 ^ n26522;
  assign n26523 = ~n26521;
  assign n26524 = ~n26539;
  assign n26525 = n26549 ^ n26550;
  assign n26551 = ~n26549;
  assign n26528 = ~n26561;
  assign n26557 = n26578 ^ n24171;
  assign n26579 = ~n26578;
  assign n26416 = n26429 & n26430;
  assign n26364 = ~n26431;
  assign n26441 = n26448 & n26418;
  assign n26417 = n26448 & n26420;
  assign n22488 = n26453 ^ n26454;
  assign n26472 = n26485 & n26486;
  assign n26456 = ~n26493;
  assign n26474 = n202 ^ n26500;
  assign n26515 = n26523 & n26524;
  assign n26478 = n26525 ^ n26526;
  assign n26540 = n26551 & n26552;
  assign n23072 = n26556 ^ n26557;
  assign n26577 = n26579 & n26580;
  assign n26389 = ~n26416;
  assign n26398 = n26417 ^ n26418;
  assign n24645 = n23520 ^ n22488;
  assign n26419 = ~n26441;
  assign n22577 = ~n22488;
  assign n26455 = ~n26472;
  assign n26400 = n26473 ^ n26474;
  assign n26475 = ~n26474;
  assign n26503 = n26478 & n8107;
  assign n26501 = ~n26515;
  assign n26504 = ~n26478;
  assign n26465 = n26533 ^ n23072;
  assign n26527 = ~n26540;
  assign n23060 = ~n23072;
  assign n26558 = ~n26577;
  assign n26391 = n26398 & n294;
  assign n26296 = n24645 ^ n24620;
  assign n26390 = ~n26398;
  assign n26409 = n26419 & n26420;
  assign n26432 = n26455 & n26456;
  assign n26422 = n26475 & n26476;
  assign n26477 = n26501 & n26502;
  assign n26480 = ~n26503;
  assign n26494 = n26504 & n201;
  assign n26510 = n26465 & n26516;
  assign n26517 = n26527 & n26528;
  assign n26511 = ~n26465;
  assign n26534 = n26558 & n26559;
  assign n26377 = n26390 & n2545;
  assign n26334 = ~n26391;
  assign n26378 = ~n26409;
  assign n26399 = n26432 ^ n23449;
  assign n26434 = n26432 & n23449;
  assign n26433 = ~n26432;
  assign n26449 = n26477 ^ n26478;
  assign n26479 = ~n26477;
  assign n26451 = ~n26494;
  assign n26495 = ~n26510;
  assign n26505 = n26511 & n26497;
  assign n26496 = ~n26517;
  assign n26512 = n26534 ^ n26535;
  assign n26536 = ~n26534;
  assign n26365 = ~n26377;
  assign n26351 = n26378 ^ n26379;
  assign n26376 = n26389 & n26378;
  assign n22455 = n26399 ^ n26400;
  assign n26421 = n26433 & n23415;
  assign n26410 = ~n26434;
  assign n26423 = n201 ^ n26449;
  assign n26463 = n26479 & n26480;
  assign n26487 = n26495 & n26496;
  assign n26464 = n26496 ^ n26497;
  assign n26467 = ~n26505;
  assign n23017 = n24111 ^ n26512;
  assign n26529 = n26536 & n26537;
  assign n26285 = n26351 ^ n26352;
  assign n26353 = n26365 & n26332;
  assign n26331 = n26365 & n26334;
  assign n24600 = n22455 ^ n23415;
  assign n26363 = ~n26376;
  assign n22493 = ~n22455;
  assign n26401 = n26410 & n26400;
  assign n26381 = ~n26421;
  assign n26318 = n26422 ^ n26423;
  assign n26366 = n26423 & n26422;
  assign n26450 = ~n26463;
  assign n26425 = n26464 ^ n26465;
  assign n26466 = ~n26487;
  assign n26445 = n26488 ^ n23017;
  assign n23005 = ~n23017;
  assign n26513 = ~n26529;
  assign n26314 = n26285 & n293;
  assign n26297 = n26331 ^ n26332;
  assign n26194 = n24600 ^ n24591;
  assign n26313 = ~n26285;
  assign n26333 = ~n26353;
  assign n26329 = n26363 & n26364;
  assign n26380 = ~n26401;
  assign n26392 = n26318 & n23409;
  assign n26393 = ~n26318;
  assign n26424 = n26450 & n26451;
  assign n26442 = n26425 & n8067;
  assign n26443 = ~n26425;
  assign n26444 = n26466 & n26467;
  assign n26458 = n26445 & n26468;
  assign n26457 = ~n26445;
  assign n26489 = n26513 & n26514;
  assign n24597 = n26297 ^ n24615;
  assign n26211 = n26297 & n24615;
  assign n26305 = n26313 & n2430;
  assign n26251 = ~n26314;
  assign n26295 = n26329 ^ n26330;
  assign n26315 = n26333 & n26334;
  assign n26337 = n26329 & n26330;
  assign n26335 = ~n26329;
  assign n26354 = n26380 & n26381;
  assign n26320 = ~n26392;
  assign n26382 = n26393 & n23368;
  assign n26394 = n26424 ^ n26425;
  assign n26427 = ~n26424;
  assign n26426 = ~n26442;
  assign n26435 = n26443 & n200;
  assign n26411 = n26444 ^ n26445;
  assign n26446 = ~n26444;
  assign n26452 = n26457 & n26412;
  assign n26447 = ~n26458;
  assign n26459 = n26489 ^ n26490;
  assign n26491 = ~n26489;
  assign n26264 = ~n24597;
  assign n26197 = n26295 ^ n26296;
  assign n26283 = ~n26305;
  assign n26284 = ~n26315;
  assign n26316 = n26335 & n26336;
  assign n26304 = ~n26337;
  assign n26317 = n26354 ^ n23368;
  assign n26355 = ~n26354;
  assign n26356 = ~n26382;
  assign n26367 = n200 ^ n26394;
  assign n26341 = n26411 ^ n26412;
  assign n26413 = n26426 & n26427;
  assign n26396 = ~n26435;
  assign n26436 = n26446 & n26447;
  assign n26415 = ~n26452;
  assign n22911 = n24071 ^ n26459;
  assign n26481 = n26491 & n26492;
  assign n26263 = n26197 & n292;
  assign n26262 = ~n26197;
  assign n26271 = n26283 & n26284;
  assign n26249 = n26284 ^ n26285;
  assign n26298 = n26304 & n26296;
  assign n26270 = ~n26316;
  assign n22416 = n26317 ^ n26318;
  assign n26345 = n26355 & n26356;
  assign n26253 = n26366 ^ n26367;
  assign n26299 = n26367 & n26366;
  assign n26384 = n26341 & n215;
  assign n26383 = ~n26341;
  assign n26395 = ~n26413;
  assign n26414 = ~n26436;
  assign n26386 = n26437 ^ n22911;
  assign n22960 = ~n22911;
  assign n26460 = ~n26481;
  assign n26212 = n293 ^ n26249;
  assign n26247 = n26262 & n2338;
  assign n26180 = ~n26263;
  assign n26265 = n22416 & n24597;
  assign n26250 = ~n26271;
  assign n24581 = n23409 ^ n22416;
  assign n26269 = ~n26298;
  assign n22403 = ~n22416;
  assign n26319 = ~n26345;
  assign n26338 = n26253 & n23353;
  assign n26339 = ~n26253;
  assign n26371 = n26383 & n8015;
  assign n26323 = ~n26384;
  assign n26368 = n26395 & n26396;
  assign n26385 = n26414 & n26415;
  assign n26402 = n26386 & n26360;
  assign n26403 = ~n26386;
  assign n26438 = n26460 & n26461;
  assign n24568 = n26211 ^ n26212;
  assign n26122 = n26212 & n26211;
  assign n26213 = ~n26247;
  assign n26233 = n26250 & n26251;
  assign n26107 = n24581 ^ n24566;
  assign n26248 = n22403 & n26264;
  assign n24599 = ~n26265;
  assign n26231 = n26269 & n26270;
  assign n26286 = n26319 & n26320;
  assign n26255 = ~n26338;
  assign n26321 = n26339 & n23348;
  assign n26340 = n215 ^ n26368;
  assign n26357 = ~n26371;
  assign n26358 = ~n26368;
  assign n26359 = n26385 ^ n26386;
  assign n26388 = ~n26385;
  assign n26387 = ~n26402;
  assign n26397 = n26403 & n26404;
  assign n26406 = n26438 ^ n24080;
  assign n26439 = ~n26438;
  assign n26177 = ~n24568;
  assign n26127 = ~n26122;
  assign n26217 = n26107 & n26143;
  assign n26193 = n26231 ^ n26232;
  assign n26196 = ~n26233;
  assign n26215 = ~n26107;
  assign n24608 = ~n26248;
  assign n26236 = n26231 & n26232;
  assign n26234 = ~n26231;
  assign n26252 = n26286 ^ n23348;
  assign n26287 = ~n26286;
  assign n26288 = ~n26321;
  assign n26300 = n26340 ^ n26341;
  assign n26346 = n26357 & n26358;
  assign n26290 = n26359 ^ n26360;
  assign n26372 = n26387 & n26388;
  assign n26362 = ~n26397;
  assign n22871 = n26405 ^ n26406;
  assign n26428 = n26439 & n26440;
  assign n26141 = n26193 ^ n26194;
  assign n26166 = n26196 ^ n26197;
  assign n26195 = n26213 & n26196;
  assign n26199 = n26215 & n26216;
  assign n26145 = ~n26217;
  assign n26228 = n26234 & n26235;
  assign n26214 = ~n26236;
  assign n22354 = n26252 ^ n26253;
  assign n26272 = n26287 & n26288;
  assign n26184 = n26299 ^ n26300;
  assign n26301 = ~n26300;
  assign n26324 = n26290 & n7981;
  assign n26322 = ~n26346;
  assign n26325 = ~n26290;
  assign n26361 = ~n26372;
  assign n22941 = ~n22871;
  assign n26407 = ~n26428;
  assign n26123 = n292 ^ n26166;
  assign n26164 = n26141 & n291;
  assign n26178 = n22354 & n24568;
  assign n26163 = ~n26141;
  assign n26179 = ~n26195;
  assign n26109 = ~n26199;
  assign n26198 = n26214 & n26194;
  assign n24547 = n23353 ^ n22354;
  assign n26182 = ~n26228;
  assign n22285 = ~n22354;
  assign n26254 = ~n26272;
  assign n26267 = n26184 & n23319;
  assign n26266 = ~n26184;
  assign n26221 = n26301 & n26299;
  assign n26289 = n26322 & n26323;
  assign n26291 = ~n26324;
  assign n26306 = n26325 & n214;
  assign n26326 = n26361 & n26362;
  assign n26327 = n26369 ^ n22941;
  assign n26373 = n26407 & n26408;
  assign n26104 = n26122 ^ n26123;
  assign n26126 = ~n26123;
  assign n26157 = n26163 & n2210;
  assign n26095 = ~n26164;
  assign n26165 = n22285 & n26177;
  assign n24571 = ~n26178;
  assign n26140 = n26179 & n26180;
  assign n26034 = n24547 ^ n24540;
  assign n26181 = ~n26198;
  assign n26218 = n26254 & n26255;
  assign n26256 = n26266 & n23268;
  assign n26220 = ~n26267;
  assign n26257 = n26289 ^ n26290;
  assign n26292 = ~n26289;
  assign n26259 = ~n26306;
  assign n26293 = n26326 ^ n26327;
  assign n26308 = ~n26326;
  assign n26342 = n26327 & n26294;
  assign n26343 = ~n26327;
  assign n26348 = n26373 ^ n24010;
  assign n26374 = ~n26373;
  assign n24533 = ~n26104;
  assign n26069 = n26126 & n26127;
  assign n26105 = n26140 ^ n26141;
  assign n26124 = ~n26157;
  assign n26146 = n26034 & n26158;
  assign n24585 = ~n26165;
  assign n26125 = ~n26140;
  assign n26147 = ~n26034;
  assign n26142 = n26181 & n26182;
  assign n26183 = n26218 ^ n23319;
  assign n26219 = ~n26218;
  assign n26186 = ~n26256;
  assign n26222 = n214 ^ n26257;
  assign n26273 = n26291 & n26292;
  assign n26224 = n26293 ^ n26294;
  assign n26307 = ~n26342;
  assign n26328 = n26343 & n26344;
  assign n22827 = n26347 ^ n26348;
  assign n26370 = n26374 & n26375;
  assign n26070 = n291 ^ n26105;
  assign n26118 = n26124 & n26125;
  assign n26106 = n26142 ^ n26143;
  assign n26036 = ~n26146;
  assign n26129 = n26147 & n26074;
  assign n26144 = ~n26142;
  assign n22209 = n26183 ^ n26184;
  assign n26200 = n26219 & n26220;
  assign n26111 = n26221 ^ n26222;
  assign n26151 = n26222 & n26221;
  assign n26260 = n26224 & n7930;
  assign n26258 = ~n26273;
  assign n26261 = ~n26224;
  assign n26302 = n26307 & n26308;
  assign n26203 = n26309 ^ n22827;
  assign n26275 = ~n26328;
  assign n22908 = ~n22827;
  assign n26349 = ~n26370;
  assign n24503 = n26069 ^ n26070;
  assign n25968 = n26070 & n26069;
  assign n26093 = n22209 & n26104;
  assign n26045 = n26106 ^ n26107;
  assign n26094 = ~n26118;
  assign n26076 = ~n26129;
  assign n26128 = n26144 & n26145;
  assign n22262 = ~n22209;
  assign n26187 = n26111 & n23230;
  assign n26185 = ~n26200;
  assign n26188 = ~n26111;
  assign n26223 = n26258 & n26259;
  assign n26225 = ~n26260;
  assign n26237 = n26261 & n213;
  assign n26276 = n26203 & n26239;
  assign n26274 = ~n26302;
  assign n26277 = ~n26203;
  assign n26310 = n26349 & n26350;
  assign n26031 = ~n24503;
  assign n26071 = n26045 & n2109;
  assign n24551 = ~n26093;
  assign n26087 = n22262 & n24533;
  assign n26088 = n26094 & n26095;
  assign n26072 = ~n26045;
  assign n26108 = ~n26128;
  assign n24518 = n22262 ^ n23268;
  assign n26148 = n26185 & n26186;
  assign n26113 = ~n26187;
  assign n26167 = n26188 & n23275;
  assign n26189 = n26223 ^ n26224;
  assign n26226 = ~n26223;
  assign n26191 = ~n26237;
  assign n26238 = n26274 & n26275;
  assign n26205 = ~n26276;
  assign n26268 = n26277 & n26278;
  assign n26280 = n26310 ^ n23970;
  assign n26311 = ~n26310;
  assign n26043 = ~n26071;
  assign n26052 = n26072 & n290;
  assign n24538 = ~n26087;
  assign n26044 = ~n26088;
  assign n25961 = n24518 ^ n24479;
  assign n26073 = n26108 & n26109;
  assign n26110 = n26148 ^ n23275;
  assign n26149 = ~n26148;
  assign n26150 = ~n26167;
  assign n26152 = n213 ^ n26189;
  assign n26201 = n26225 & n26226;
  assign n26202 = n26238 ^ n26239;
  assign n26241 = ~n26238;
  assign n26240 = ~n26268;
  assign n22779 = n26279 ^ n26280;
  assign n26303 = n26311 & n26312;
  assign n26032 = n26043 & n26044;
  assign n26009 = n26044 ^ n26045;
  assign n26011 = ~n26052;
  assign n26033 = n26073 ^ n26074;
  assign n26054 = n25961 & n25998;
  assign n26055 = ~n25961;
  assign n26075 = ~n26073;
  assign n22098 = n26110 ^ n26111;
  assign n26130 = n26149 & n26150;
  assign n26038 = n26151 ^ n26152;
  assign n26080 = n26152 & n26151;
  assign n26190 = ~n26201;
  assign n26154 = n26202 ^ n26203;
  assign n26229 = n26240 & n26241;
  assign n26133 = n26242 ^ n22779;
  assign n22869 = ~n22779;
  assign n26281 = ~n26303;
  assign n25969 = n290 ^ n26009;
  assign n26020 = n22098 & n26031;
  assign n26010 = ~n26032;
  assign n25971 = n26033 ^ n26034;
  assign n26000 = ~n26054;
  assign n26046 = n26055 & n26056;
  assign n26053 = n26075 & n26076;
  assign n24482 = n22098 ^ n23230;
  assign n22196 = ~n22098;
  assign n26112 = ~n26130;
  assign n26083 = ~n26080;
  assign n26153 = n26190 & n26191;
  assign n26168 = n26154 & n7900;
  assign n26169 = ~n26154;
  assign n26206 = n26133 & n26227;
  assign n26204 = ~n26229;
  assign n26207 = ~n26133;
  assign n26243 = n26281 & n26282;
  assign n24472 = n25968 ^ n25969;
  assign n25892 = n25969 & n25968;
  assign n25970 = n26010 & n26011;
  assign n25996 = n25971 & n289;
  assign n24505 = ~n26020;
  assign n25995 = ~n25971;
  assign n25887 = n24482 ^ n24444;
  assign n26030 = n22196 & n24503;
  assign n25963 = ~n26046;
  assign n26035 = ~n26053;
  assign n26077 = n26112 & n26113;
  assign n26114 = n26153 ^ n26154;
  assign n26155 = ~n26153;
  assign n26156 = ~n26168;
  assign n26159 = n26169 & n212;
  assign n26170 = n26204 & n26205;
  assign n26135 = ~n26206;
  assign n26192 = n26207 & n26171;
  assign n26208 = n26243 ^ n26244;
  assign n26245 = ~n26243;
  assign n25931 = ~n24472;
  assign n25895 = ~n25892;
  assign n25933 = n25970 ^ n25971;
  assign n25959 = ~n25970;
  assign n25981 = n25995 & n2069;
  assign n25921 = ~n25996;
  assign n26003 = n25887 & n25925;
  assign n26001 = ~n25887;
  assign n24523 = ~n26030;
  assign n25997 = n26035 & n26036;
  assign n26037 = n26077 ^ n23217;
  assign n26079 = n26077 & n23217;
  assign n26078 = ~n26077;
  assign n26081 = n212 ^ n26114;
  assign n26131 = n26155 & n26156;
  assign n26116 = ~n26159;
  assign n26132 = n26170 ^ n26171;
  assign n26173 = ~n26170;
  assign n26172 = ~n26192;
  assign n22760 = n26208 ^ n23968;
  assign n26230 = n26245 & n26246;
  assign n25893 = n289 ^ n25933;
  assign n25958 = ~n25981;
  assign n25960 = n25997 ^ n25998;
  assign n25983 = n26001 & n26002;
  assign n25927 = ~n26003;
  assign n25999 = ~n25997;
  assign n22127 = n26037 ^ n26038;
  assign n26057 = n26078 & n23237;
  assign n26047 = ~n26079;
  assign n25934 = n26080 ^ n26081;
  assign n26082 = ~n26081;
  assign n26115 = ~n26131;
  assign n26085 = n26132 ^ n26133;
  assign n26160 = n26172 & n26173;
  assign n22849 = ~n22760;
  assign n26209 = ~n26230;
  assign n24435 = n25892 ^ n25893;
  assign n25894 = ~n25893;
  assign n25919 = n22127 & n25931;
  assign n25946 = n25958 & n25959;
  assign n25883 = n25960 ^ n25961;
  assign n25889 = ~n25983;
  assign n25982 = n25999 & n26000;
  assign n24450 = n23237 ^ n22127;
  assign n22081 = ~n22127;
  assign n26039 = n26047 & n26038;
  assign n26040 = n25934 & n23183;
  assign n26013 = ~n26057;
  assign n26041 = ~n25934;
  assign n26004 = n26082 & n26083;
  assign n26084 = n26115 & n26116;
  assign n26097 = n26085 & n211;
  assign n26096 = ~n26085;
  assign n26134 = ~n26160;
  assign n26060 = n26161 ^ n22849;
  assign n26174 = n26209 & n26210;
  assign n25859 = ~n24435;
  assign n25811 = n25894 & n25895;
  assign n24475 = ~n25919;
  assign n25922 = n25883 & n2009;
  assign n25932 = n22081 & n24472;
  assign n25920 = ~n25946;
  assign n25923 = ~n25883;
  assign n25818 = n24450 ^ n24442;
  assign n25962 = ~n25982;
  assign n26012 = ~n26039;
  assign n25974 = ~n26040;
  assign n26021 = n26041 & n23249;
  assign n26007 = ~n26004;
  assign n26042 = n26084 ^ n26085;
  assign n26059 = ~n26084;
  assign n26089 = n26096 & n7845;
  assign n26023 = ~n26097;
  assign n26098 = n26134 & n26135;
  assign n26121 = n26060 & n26099;
  assign n26119 = ~n26060;
  assign n26137 = n26174 ^ n23937;
  assign n26175 = ~n26174;
  assign n25882 = n25920 & n25921;
  assign n25885 = ~n25922;
  assign n25906 = n25923 & n288;
  assign n24489 = ~n25932;
  assign n25924 = n25962 & n25963;
  assign n25972 = n26012 & n26013;
  assign n25937 = ~n26021;
  assign n26005 = n211 ^ n26042;
  assign n26058 = ~n26089;
  assign n26061 = n26098 ^ n26099;
  assign n26090 = ~n26098;
  assign n26117 = n26119 & n26120;
  assign n26050 = ~n26121;
  assign n22802 = n26136 ^ n26137;
  assign n26162 = n26175 & n26176;
  assign n25847 = n25882 ^ n25883;
  assign n25884 = ~n25882;
  assign n25849 = ~n25906;
  assign n25886 = n25924 ^ n25925;
  assign n25926 = ~n25924;
  assign n25935 = n25972 ^ n23249;
  assign n25973 = ~n25972;
  assign n25862 = n26004 ^ n26005;
  assign n26006 = ~n26005;
  assign n26048 = n26058 & n26059;
  assign n25985 = n26060 ^ n26061;
  assign n25977 = n26100 ^ n22802;
  assign n26091 = ~n26117;
  assign n22677 = ~n22802;
  assign n26138 = ~n26162;
  assign n25812 = n288 ^ n25847;
  assign n25874 = n25884 & n25885;
  assign n25814 = n25886 ^ n25887;
  assign n25907 = n25926 & n25927;
  assign n22065 = n25934 ^ n25935;
  assign n25964 = n25973 & n25974;
  assign n25965 = n25862 & n23211;
  assign n25966 = ~n25862;
  assign n25908 = n26006 & n26007;
  assign n26024 = n25985 & n7794;
  assign n26022 = ~n26048;
  assign n26025 = ~n25985;
  assign n26062 = n25977 & n26016;
  assign n26086 = n26090 & n26091;
  assign n26063 = ~n25977;
  assign n26101 = n26138 & n26139;
  assign n24400 = n25811 ^ n25812;
  assign n25734 = n25812 & n25811;
  assign n25850 = n25814 & n1922;
  assign n25860 = n22065 & n24435;
  assign n25848 = ~n25874;
  assign n25851 = ~n25814;
  assign n24415 = n22065 ^ n23249;
  assign n25888 = ~n25907;
  assign n22054 = ~n22065;
  assign n25936 = ~n25964;
  assign n25864 = ~n25965;
  assign n25947 = n25966 & n23151;
  assign n25984 = n26022 & n26023;
  assign n25986 = ~n26024;
  assign n26014 = n26025 & n210;
  assign n26018 = ~n26062;
  assign n26051 = n26063 & n26064;
  assign n26049 = ~n26086;
  assign n26066 = n26101 ^ n23909;
  assign n26102 = ~n26101;
  assign n25774 = ~n24400;
  assign n25813 = n25848 & n25849;
  assign n25816 = ~n25850;
  assign n25834 = n25851 & n303;
  assign n25846 = n22054 & n25859;
  assign n24437 = ~n25860;
  assign n25706 = n24415 ^ n24408;
  assign n25852 = n25888 & n25889;
  assign n25896 = n25936 & n25937;
  assign n25898 = ~n25947;
  assign n25948 = n25984 ^ n25985;
  assign n25987 = ~n25984;
  assign n25950 = ~n26014;
  assign n26015 = n26049 & n26050;
  assign n25979 = ~n26051;
  assign n22729 = n26065 ^ n26066;
  assign n26092 = n26102 & n26103;
  assign n25776 = n25813 ^ n25814;
  assign n25815 = ~n25813;
  assign n25778 = ~n25834;
  assign n24453 = ~n25846;
  assign n25817 = n25852 ^ n25853;
  assign n25856 = n25852 & n25853;
  assign n25854 = ~n25852;
  assign n25861 = n25896 ^ n23151;
  assign n25897 = ~n25896;
  assign n25909 = n210 ^ n25948;
  assign n25975 = n25986 & n25987;
  assign n25976 = n26015 ^ n26016;
  assign n25901 = n26026 ^ n22729;
  assign n26017 = ~n26015;
  assign n22717 = ~n22729;
  assign n26067 = ~n26092;
  assign n25735 = n303 ^ n25776;
  assign n25797 = n25815 & n25816;
  assign n25737 = n25817 ^ n25818;
  assign n25835 = n25854 & n25855;
  assign n25822 = ~n25856;
  assign n22010 = n25861 ^ n25862;
  assign n25890 = n25897 & n25898;
  assign n25786 = n25908 ^ n25909;
  assign n25836 = n25909 & n25908;
  assign n25949 = ~n25975;
  assign n25911 = n25976 ^ n25977;
  assign n25990 = n25901 & n25941;
  assign n26008 = n26017 & n26018;
  assign n25988 = ~n25901;
  assign n26027 = n26067 & n26068;
  assign n24363 = n25734 ^ n25735;
  assign n25658 = n25735 & n25734;
  assign n25775 = n22010 & n24400;
  assign n25780 = n25737 & n302;
  assign n25777 = ~n25797;
  assign n25779 = ~n25737;
  assign n25819 = n25822 & n25818;
  assign n24378 = n22010 ^ n23211;
  assign n25784 = ~n25835;
  assign n21971 = ~n22010;
  assign n25863 = ~n25890;
  assign n25910 = n25949 & n25950;
  assign n25938 = n25911 & n7739;
  assign n25939 = ~n25911;
  assign n25980 = n25988 & n25989;
  assign n25903 = ~n25990;
  assign n25978 = ~n26008;
  assign n25991 = n26027 ^ n23848;
  assign n26028 = ~n26027;
  assign n25699 = ~n24363;
  assign n25759 = n21971 & n25774;
  assign n24402 = ~n25775;
  assign n25736 = n25777 & n25778;
  assign n25760 = n25779 & n1874;
  assign n25702 = ~n25780;
  assign n25608 = n24378 ^ n24359;
  assign n25783 = ~n25819;
  assign n25823 = n25863 & n25864;
  assign n25875 = n25910 ^ n25911;
  assign n25912 = ~n25910;
  assign n25913 = ~n25938;
  assign n25928 = n25939 & n209;
  assign n25940 = n25978 & n25979;
  assign n25943 = ~n25980;
  assign n22671 = n25991 ^ n25992;
  assign n26019 = n26028 & n26029;
  assign n25700 = n25736 ^ n25737;
  assign n24418 = ~n25759;
  assign n25738 = ~n25736;
  assign n25739 = ~n25760;
  assign n25749 = n25608 & n25645;
  assign n25750 = ~n25608;
  assign n25744 = n25783 & n25784;
  assign n25785 = n25823 ^ n23114;
  assign n25825 = n25823 & n23114;
  assign n25824 = ~n25823;
  assign n25837 = n209 ^ n25875;
  assign n25899 = n25912 & n25913;
  assign n25877 = ~n25928;
  assign n25900 = n25940 ^ n25941;
  assign n25868 = n25951 ^ n22671;
  assign n25942 = ~n25940;
  assign n25952 = n22671 & n25967;
  assign n22547 = ~n22671;
  assign n25993 = ~n26019;
  assign n25659 = n302 ^ n25700;
  assign n25720 = n25738 & n25739;
  assign n25705 = n25744 ^ n25745;
  assign n25647 = ~n25749;
  assign n25741 = n25750 & n25751;
  assign n25748 = n25744 & n25745;
  assign n25746 = ~n25744;
  assign n21953 = n25785 ^ n25786;
  assign n25820 = n25824 & n23146;
  assign n25798 = ~n25825;
  assign n25684 = n25836 ^ n25837;
  assign n25763 = n25837 & n25836;
  assign n25876 = ~n25899;
  assign n25839 = n25900 ^ n25901;
  assign n25915 = n25868 & n25929;
  assign n25930 = n25942 & n25943;
  assign n25914 = ~n25868;
  assign n25095 = ~n25952;
  assign n25944 = n22547 & n25953;
  assign n25954 = n25993 & n25994;
  assign n24343 = n25658 ^ n25659;
  assign n25660 = ~n25659;
  assign n25698 = n21953 & n24363;
  assign n25643 = n25705 ^ n25706;
  assign n25701 = ~n25720;
  assign n25610 = ~n25741;
  assign n25740 = n25746 & n25747;
  assign n25721 = ~n25748;
  assign n24339 = n21953 ^ n23146;
  assign n21938 = ~n21953;
  assign n25787 = n25798 & n25786;
  assign n25762 = ~n25820;
  assign n25800 = n25684 & n23128;
  assign n25799 = ~n25684;
  assign n25766 = ~n25763;
  assign n25838 = n25876 & n25877;
  assign n25865 = n25839 & n7684;
  assign n25866 = ~n25839;
  assign n25904 = n25914 & n25828;
  assign n25870 = ~n25915;
  assign n25902 = ~n25930;
  assign n25076 = ~n25944;
  assign n25916 = n25954 ^ n25955;
  assign n25956 = ~n25954;
  assign n25623 = ~n24343;
  assign n25569 = n25660 & n25658;
  assign n25666 = n25643 & n301;
  assign n24365 = ~n25698;
  assign n25679 = n21938 & n25699;
  assign n25680 = n25701 & n25702;
  assign n25665 = ~n25643;
  assign n25532 = n24339 ^ n24331;
  assign n25707 = n25721 & n25706;
  assign n25682 = ~n25740;
  assign n25761 = ~n25787;
  assign n25788 = n25799 & n23076;
  assign n25686 = ~n25800;
  assign n25801 = n25838 ^ n25839;
  assign n25840 = ~n25838;
  assign n25841 = ~n25865;
  assign n25857 = n25866 & n208;
  assign n25867 = n25902 & n25903;
  assign n25830 = ~n25904;
  assign n25905 = n25095 & n25076;
  assign n22474 = n25916 ^ n23809;
  assign n25945 = n25956 & n25957;
  assign n25661 = n25665 & n1851;
  assign n25593 = ~n25666;
  assign n24382 = ~n25679;
  assign n25628 = ~n25680;
  assign n25667 = n25532 & n25574;
  assign n25668 = ~n25532;
  assign n25681 = ~n25707;
  assign n25722 = n25761 & n25762;
  assign n25724 = ~n25788;
  assign n25764 = n208 ^ n25801;
  assign n25826 = n25840 & n25841;
  assign n25803 = ~n25857;
  assign n25827 = n25867 ^ n25868;
  assign n25869 = ~n25867;
  assign n25878 = n22474 & n25891;
  assign n25093 = ~n25905;
  assign n22612 = ~n22474;
  assign n25917 = ~n25945;
  assign n25606 = n25628 ^ n25643;
  assign n25627 = ~n25661;
  assign n25534 = ~n25667;
  assign n25662 = n25668 & n25669;
  assign n25644 = n25681 & n25682;
  assign n25683 = n25722 ^ n23076;
  assign n25723 = ~n25722;
  assign n25611 = n25763 ^ n25764;
  assign n25765 = ~n25764;
  assign n25802 = ~n25826;
  assign n25728 = n25827 ^ n25828;
  assign n25858 = n25869 & n25870;
  assign n25792 = n25871 ^ n22612;
  assign n25038 = ~n25878;
  assign n25872 = n22612 & n25060;
  assign n25879 = n25917 & n25918;
  assign n25570 = n301 ^ n25606;
  assign n25624 = n25627 & n25628;
  assign n25607 = n25644 ^ n25645;
  assign n25576 = ~n25662;
  assign n25646 = ~n25644;
  assign n21910 = n25683 ^ n25684;
  assign n25708 = n25723 & n25724;
  assign n25726 = n25611 & n23082;
  assign n25725 = ~n25611;
  assign n25687 = n25765 & n25766;
  assign n25767 = n25802 & n25803;
  assign n25790 = n25728 & n223;
  assign n25789 = ~n25728;
  assign n25831 = n25792 & n25755;
  assign n25829 = ~n25858;
  assign n25832 = ~n25792;
  assign n25062 = ~n25872;
  assign n25843 = n25879 ^ n23743;
  assign n25880 = ~n25879;
  assign n24283 = n25569 ^ n25570;
  assign n25469 = n25570 & n25569;
  assign n25548 = n25607 ^ n25608;
  assign n25605 = n21910 & n25623;
  assign n25592 = ~n25624;
  assign n25629 = n25646 & n25647;
  assign n24299 = n23128 ^ n21910;
  assign n21876 = ~n21910;
  assign n25685 = ~n25708;
  assign n25709 = n25725 & n23095;
  assign n25650 = ~n25726;
  assign n25690 = ~n25687;
  assign n25727 = n223 ^ n25767;
  assign n25752 = ~n25767;
  assign n25781 = n25789 & n7559;
  assign n25711 = ~n25790;
  assign n25791 = n25829 & n25830;
  assign n25794 = ~n25831;
  assign n25821 = n25832 & n25833;
  assign n22444 = n25842 ^ n25843;
  assign n25873 = n25880 & n25881;
  assign n25528 = ~n24283;
  assign n25571 = n25548 & n1797;
  assign n25588 = n25592 & n25593;
  assign n25572 = ~n25548;
  assign n24325 = ~n25605;
  assign n25458 = n24299 ^ n24291;
  assign n25622 = n21876 & n24343;
  assign n25609 = ~n25629;
  assign n25648 = n25685 & n25686;
  assign n25614 = ~n25709;
  assign n25688 = n25727 ^ n25728;
  assign n25753 = ~n25781;
  assign n25754 = n25791 ^ n25792;
  assign n25715 = n22444 ^ n25804;
  assign n25793 = ~n25791;
  assign n25757 = ~n25821;
  assign n25806 = n22444 & n25018;
  assign n22468 = ~n22444;
  assign n25844 = ~n25873;
  assign n25546 = ~n25571;
  assign n25552 = n25572 & n300;
  assign n25547 = ~n25588;
  assign n25577 = n25458 & n25589;
  assign n25578 = ~n25458;
  assign n25573 = n25609 & n25610;
  assign n24345 = ~n25622;
  assign n25612 = n25648 ^ n23095;
  assign n25649 = ~n25648;
  assign n25535 = n25687 ^ n25688;
  assign n25689 = ~n25688;
  assign n25742 = n25752 & n25753;
  assign n25671 = n25754 ^ n25755;
  assign n25770 = n25715 & n25675;
  assign n25782 = n25793 & n25794;
  assign n25768 = ~n25715;
  assign n25795 = n22468 & n25805;
  assign n25020 = ~n25806;
  assign n25807 = n25844 & n25845;
  assign n25530 = n25546 & n25547;
  assign n25508 = n25547 ^ n25548;
  assign n25510 = ~n25552;
  assign n25531 = n25573 ^ n25574;
  assign n25460 = ~n25577;
  assign n25554 = n25578 & n25497;
  assign n25575 = ~n25573;
  assign n21867 = n25611 ^ n25612;
  assign n25630 = n25649 & n25650;
  assign n25651 = n25535 & n23072;
  assign n25652 = ~n25535;
  assign n25594 = n25689 & n25690;
  assign n25712 = n25671 & n7536;
  assign n25710 = ~n25742;
  assign n25713 = ~n25671;
  assign n25758 = n25768 & n25769;
  assign n25717 = ~n25770;
  assign n25756 = ~n25782;
  assign n24999 = ~n25795;
  assign n25771 = n25807 ^ n25808;
  assign n25809 = ~n25807;
  assign n25470 = n300 ^ n25508;
  assign n25509 = ~n25530;
  assign n25473 = n25531 ^ n25532;
  assign n25529 = n21867 & n24283;
  assign n25499 = ~n25554;
  assign n25553 = n25575 & n25576;
  assign n24257 = n21867 ^ n23095;
  assign n21860 = ~n21867;
  assign n25613 = ~n25630;
  assign n25538 = ~n25651;
  assign n25631 = n25652 & n23060;
  assign n25670 = n25710 & n25711;
  assign n25673 = ~n25712;
  assign n25703 = n25713 & n222;
  assign n25714 = n25756 & n25757;
  assign n25677 = ~n25758;
  assign n22334 = n25771 ^ n23656;
  assign n25796 = n25809 & n25810;
  assign n24261 = n25469 ^ n25470;
  assign n25471 = ~n25470;
  assign n25472 = n25509 & n25510;
  assign n25494 = n25473 & n1764;
  assign n25495 = ~n25473;
  assign n25514 = n21860 & n25528;
  assign n24285 = ~n25529;
  assign n25391 = n24257 ^ n24239;
  assign n25533 = ~n25553;
  assign n25579 = n25613 & n25614;
  assign n25581 = ~n25631;
  assign n25632 = n25670 ^ n25671;
  assign n25672 = ~n25670;
  assign n25634 = ~n25703;
  assign n25674 = n25714 ^ n25715;
  assign n25601 = n25729 ^ n22334;
  assign n25716 = ~n25714;
  assign n25730 = n22334 & n25743;
  assign n22469 = ~n22334;
  assign n25772 = ~n25796;
  assign n25439 = ~n24261;
  assign n25397 = n25471 & n25469;
  assign n25440 = n25472 ^ n25473;
  assign n25474 = ~n25472;
  assign n25475 = ~n25494;
  assign n25480 = n25495 & n299;
  assign n25500 = n25391 & n25427;
  assign n24304 = ~n25514;
  assign n25501 = ~n25391;
  assign n25496 = n25533 & n25534;
  assign n25536 = n25579 ^ n23072;
  assign n25580 = ~n25579;
  assign n25595 = n222 ^ n25632;
  assign n25663 = n25672 & n25673;
  assign n25597 = n25674 ^ n25675;
  assign n25693 = n25601 & n25638;
  assign n25704 = n25716 & n25717;
  assign n25691 = ~n25601;
  assign n24986 = ~n25730;
  assign n25718 = n22469 & n24961;
  assign n25731 = n25772 & n25773;
  assign n25398 = n299 ^ n25440;
  assign n25400 = ~n25397;
  assign n25456 = n25474 & n25475;
  assign n25442 = ~n25480;
  assign n25457 = n25496 ^ n25497;
  assign n25429 = ~n25500;
  assign n25482 = n25501 & n25502;
  assign n25498 = ~n25496;
  assign n21771 = n25535 ^ n25536;
  assign n25555 = n25580 & n25581;
  assign n25582 = n25594 ^ n25595;
  assign n25515 = n25595 & n25594;
  assign n25635 = n25597 & n7384;
  assign n25633 = ~n25663;
  assign n25636 = ~n25597;
  assign n25678 = n25691 & n25692;
  assign n25640 = ~n25693;
  assign n25676 = ~n25704;
  assign n24964 = ~n25718;
  assign n25695 = n25731 ^ n23670;
  assign n25732 = ~n25731;
  assign n24202 = n25397 ^ n25398;
  assign n25399 = ~n25398;
  assign n25438 = n21771 & n24261;
  assign n25441 = ~n25456;
  assign n25402 = n25457 ^ n25458;
  assign n25393 = ~n25482;
  assign n25481 = n25498 & n25499;
  assign n24217 = n21771 ^ n23072;
  assign n21803 = ~n21771;
  assign n25537 = ~n25555;
  assign n25557 = n25582 & n23017;
  assign n25556 = ~n25582;
  assign n25518 = ~n25515;
  assign n25596 = n25633 & n25634;
  assign n25598 = ~n25635;
  assign n25625 = n25636 & n221;
  assign n25637 = n25676 & n25677;
  assign n25603 = ~n25678;
  assign n22384 = n25694 ^ n25695;
  assign n25719 = n25732 & n25733;
  assign n25368 = ~n24202;
  assign n25338 = n25399 & n25400;
  assign n24263 = ~n25438;
  assign n25423 = n21803 & n25439;
  assign n25401 = n25441 & n25442;
  assign n25425 = n25402 & n298;
  assign n25424 = ~n25402;
  assign n25334 = n24217 ^ n24171;
  assign n25459 = ~n25481;
  assign n25476 = n25537 & n25538;
  assign n25549 = n25556 & n23005;
  assign n25462 = ~n25557;
  assign n25558 = n25596 ^ n25597;
  assign n25599 = ~n25596;
  assign n25560 = ~n25625;
  assign n25600 = n25637 ^ n25638;
  assign n25524 = n25653 ^ n22384;
  assign n25639 = ~n25637;
  assign n25654 = n22384 & n25664;
  assign n22256 = ~n22384;
  assign n25696 = ~n25719;
  assign n25341 = ~n25338;
  assign n25370 = n25401 ^ n25402;
  assign n24244 = ~n25423;
  assign n25388 = ~n25401;
  assign n25408 = n25424 & n1703;
  assign n25360 = ~n25425;
  assign n25431 = n25334 & n25443;
  assign n25430 = ~n25334;
  assign n25426 = n25459 & n25460;
  assign n25503 = ~n25476;
  assign n25504 = ~n25549;
  assign n25516 = n221 ^ n25558;
  assign n25590 = n25598 & n25599;
  assign n25520 = n25600 ^ n25601;
  assign n25615 = n25524 & n25564;
  assign n25626 = n25639 & n25640;
  assign n25616 = ~n25524;
  assign n25641 = n22256 & n24945;
  assign n24928 = ~n25654;
  assign n25655 = n25696 & n25697;
  assign n25339 = n298 ^ n25370;
  assign n25389 = ~n25408;
  assign n25390 = n25426 ^ n25427;
  assign n25410 = n25430 & n25364;
  assign n25336 = ~n25431;
  assign n25428 = ~n25426;
  assign n25483 = n25503 & n25504;
  assign n25511 = n25504 & n25462;
  assign n25433 = n25515 ^ n25516;
  assign n25517 = ~n25516;
  assign n25561 = n25520 & n7394;
  assign n25559 = ~n25590;
  assign n25562 = ~n25520;
  assign n25566 = ~n25615;
  assign n25604 = n25616 & n25617;
  assign n25602 = ~n25626;
  assign n24947 = ~n25641;
  assign n25619 = n25655 ^ n23582;
  assign n25656 = ~n25655;
  assign n24181 = n25338 ^ n25339;
  assign n25340 = ~n25339;
  assign n25376 = n25388 & n25389;
  assign n25330 = n25390 ^ n25391;
  assign n25366 = ~n25410;
  assign n25409 = n25428 & n25429;
  assign n25461 = ~n25483;
  assign n25477 = ~n25511;
  assign n25404 = ~n25433;
  assign n25445 = n25517 & n25518;
  assign n25519 = n25559 & n25560;
  assign n25522 = ~n25561;
  assign n25550 = n25562 & n220;
  assign n25563 = n25602 & n25603;
  assign n25526 = ~n25604;
  assign n22153 = n25618 ^ n25619;
  assign n25642 = n25656 & n25657;
  assign n25315 = ~n24181;
  assign n25277 = n25340 & n25341;
  assign n25361 = n25330 & n1678;
  assign n25359 = ~n25376;
  assign n25362 = ~n25330;
  assign n25392 = ~n25409;
  assign n25432 = n25461 & n25462;
  assign n21773 = n25476 ^ n25477;
  assign n25463 = ~n25445;
  assign n25484 = n25519 ^ n25520;
  assign n25521 = ~n25519;
  assign n25486 = ~n25550;
  assign n25523 = n25563 ^ n25564;
  assign n25452 = n25583 ^ n22153;
  assign n25565 = ~n25563;
  assign n25584 = n22153 & n25591;
  assign n22271 = ~n22153;
  assign n25620 = ~n25642;
  assign n25280 = ~n25277;
  assign n25329 = n25359 & n25360;
  assign n25332 = ~n25361;
  assign n25348 = n25362 & n297;
  assign n25358 = n25368 & n21773;
  assign n25363 = n25392 & n25393;
  assign n24137 = n25432 ^ n25433;
  assign n24177 = n21773 ^ n23017;
  assign n25435 = n25432 & n22960;
  assign n25434 = ~n25432;
  assign n21764 = ~n21773;
  assign n25446 = n220 ^ n25484;
  assign n25512 = n25521 & n25522;
  assign n25448 = n25523 ^ n25524;
  assign n25539 = n25452 & n25490;
  assign n25551 = n25565 & n25566;
  assign n25540 = ~n25452;
  assign n24888 = ~n25584;
  assign n25567 = n22271 & n24886;
  assign n25585 = n25620 & n25621;
  assign n25306 = n25329 ^ n25330;
  assign n25331 = ~n25329;
  assign n25308 = ~n25348;
  assign n24204 = ~n25358;
  assign n25333 = n25363 ^ n25364;
  assign n25369 = n21764 & n24202;
  assign n25365 = ~n25363;
  assign n25245 = n24137 ^ n24071;
  assign n21607 = n24137 ^ n22911;
  assign n25312 = n24177 ^ n24169;
  assign n25411 = n25434 & n22911;
  assign n25403 = ~n25435;
  assign n25343 = n25445 ^ n25446;
  assign n25378 = n25446 & n25463;
  assign n25487 = n25448 & n7342;
  assign n25485 = ~n25512;
  assign n25488 = ~n25448;
  assign n25454 = ~n25539;
  assign n25527 = n25540 & n25541;
  assign n25525 = ~n25551;
  assign n24914 = ~n25567;
  assign n25542 = n25585 ^ n23556;
  assign n25586 = ~n25585;
  assign n25278 = n297 ^ n25306;
  assign n25316 = n21607 & n24181;
  assign n25320 = n25331 & n25332;
  assign n25282 = n25333 ^ n25334;
  assign n25349 = n25365 & n25366;
  assign n24221 = ~n25369;
  assign n25372 = n25312 & n25377;
  assign n21685 = ~n21607;
  assign n25371 = ~n25312;
  assign n25394 = n25403 & n25404;
  assign n25374 = ~n25411;
  assign n25413 = n25343 & n22941;
  assign n25412 = ~n25343;
  assign n25447 = n25485 & n25486;
  assign n25450 = ~n25487;
  assign n25478 = n25488 & n219;
  assign n25489 = n25525 & n25526;
  assign n25491 = ~n25527;
  assign n22228 = n25542 ^ n25543;
  assign n25568 = n25586 & n25587;
  assign n25265 = n25277 ^ n25278;
  assign n25279 = ~n25278;
  assign n25305 = n21685 & n25315;
  assign n24163 = ~n25316;
  assign n25310 = n25282 & n296;
  assign n25307 = ~n25320;
  assign n25309 = ~n25282;
  assign n25335 = ~n25349;
  assign n25367 = n25371 & n25286;
  assign n25314 = ~n25372;
  assign n25373 = ~n25394;
  assign n25405 = n25412 & n22871;
  assign n25345 = ~n25413;
  assign n25414 = n25447 ^ n25448;
  assign n25449 = ~n25447;
  assign n25416 = ~n25478;
  assign n25451 = n25489 ^ n25490;
  assign n25385 = n25505 ^ n22228;
  assign n25492 = ~n25489;
  assign n25506 = n22228 & n25513;
  assign n22124 = ~n22228;
  assign n25544 = ~n25568;
  assign n24120 = ~n25265;
  assign n25237 = n25279 & n25280;
  assign n24183 = ~n25305;
  assign n25281 = n25307 & n25308;
  assign n25298 = n25309 & n1618;
  assign n25261 = ~n25310;
  assign n25311 = n25335 & n25336;
  assign n25288 = ~n25367;
  assign n25342 = n25373 & n25374;
  assign n25318 = ~n25405;
  assign n25379 = n219 ^ n25414;
  assign n25444 = n25449 & n25450;
  assign n25381 = n25451 ^ n25452;
  assign n25466 = n25385 & n25420;
  assign n25479 = n25491 & n25492;
  assign n25464 = ~n25385;
  assign n25493 = n22124 & n24869;
  assign n24852 = ~n25506;
  assign n25507 = n25544 & n25545;
  assign n25259 = n25281 ^ n25282;
  assign n25283 = ~n25281;
  assign n25284 = ~n25298;
  assign n25285 = n25311 ^ n25312;
  assign n25313 = ~n25311;
  assign n24098 = n25342 ^ n25343;
  assign n25344 = ~n25342;
  assign n25268 = n25378 ^ n25379;
  assign n25321 = n25379 & n25378;
  assign n25417 = n25381 & n7252;
  assign n25415 = ~n25444;
  assign n25418 = ~n25381;
  assign n25455 = n25464 & n25465;
  assign n25422 = ~n25466;
  assign n25453 = ~n25479;
  assign n24871 = ~n25493;
  assign n25468 = n25507 ^ n24799;
  assign n25238 = n296 ^ n25259;
  assign n25272 = n25283 & n25284;
  assign n25222 = n25285 ^ n25286;
  assign n25299 = n25313 & n25314;
  assign n25212 = n24098 ^ n24080;
  assign n21571 = n24098 ^ n22871;
  assign n25337 = n25344 & n25345;
  assign n25350 = n25268 & n22827;
  assign n25351 = ~n25268;
  assign n25380 = n25415 & n25416;
  assign n25383 = ~n25417;
  assign n25406 = n25418 & n218;
  assign n25419 = n25453 & n25454;
  assign n25387 = ~n25455;
  assign n22106 = n25467 ^ n25468;
  assign n24083 = n25237 ^ n25238;
  assign n25203 = n25238 & n25237;
  assign n25250 = n21571 & n24120;
  assign n25263 = n25222 & n311;
  assign n25260 = ~n25272;
  assign n25262 = ~n25222;
  assign n25287 = ~n25299;
  assign n25291 = n25212 & n25194;
  assign n25292 = ~n25212;
  assign n21641 = ~n21571;
  assign n25317 = ~n25337;
  assign n25271 = ~n25350;
  assign n25346 = n25351 & n22908;
  assign n25352 = n25380 ^ n25381;
  assign n25382 = ~n25380;
  assign n25354 = ~n25406;
  assign n25384 = n25419 ^ n25420;
  assign n25328 = n25436 ^ n22106;
  assign n25395 = n25437 ^ n22106;
  assign n25421 = ~n25419;
  assign n25219 = ~n24083;
  assign n25206 = ~n25203;
  assign n24123 = ~n25250;
  assign n25239 = n25260 & n25261;
  assign n25251 = n25262 & n1559;
  assign n25224 = ~n25263;
  assign n25258 = n21641 & n25265;
  assign n25266 = n25287 & n25288;
  assign n25196 = ~n25291;
  assign n25289 = n25292 & n25293;
  assign n25294 = n25317 & n25318;
  assign n25296 = ~n25346;
  assign n25322 = n218 ^ n25352;
  assign n25375 = n25382 & n25383;
  assign n25324 = n25384 ^ n25385;
  assign n24835 = n25395 ^ n25396;
  assign n25407 = n25421 & n25422;
  assign n25221 = n311 ^ n25239;
  assign n25240 = ~n25239;
  assign n25241 = ~n25251;
  assign n24141 = ~n25258;
  assign n25264 = n25266 & n25267;
  assign n25252 = ~n25266;
  assign n25214 = ~n25289;
  assign n25269 = n25294 ^ n22827;
  assign n25295 = ~n25294;
  assign n25227 = n25321 ^ n25322;
  assign n25273 = n25322 & n25321;
  assign n25355 = n25324 & n7185;
  assign n25353 = ~n25375;
  assign n25356 = ~n25324;
  assign n25386 = ~n25407;
  assign n25204 = n25221 ^ n25222;
  assign n25232 = n25240 & n25241;
  assign n25233 = n25252 ^ n25245;
  assign n25253 = n25252 & n25234;
  assign n25244 = ~n25264;
  assign n21583 = n25268 ^ n25269;
  assign n25290 = n25295 & n25296;
  assign n25301 = n25227 & n22779;
  assign n25300 = ~n25227;
  assign n25323 = n25353 & n25354;
  assign n25326 = ~n25355;
  assign n25347 = n25356 & n217;
  assign n25357 = n25386 & n25387;
  assign n24040 = n25203 ^ n25204;
  assign n25205 = ~n25204;
  assign n25220 = n21583 & n24083;
  assign n25223 = ~n25232;
  assign n25192 = n25233 ^ n25234;
  assign n25242 = n25244 & n25245;
  assign n24057 = n21583 ^ n22827;
  assign n25226 = ~n25253;
  assign n21595 = ~n21583;
  assign n25270 = ~n25290;
  assign n25297 = n25300 & n22869;
  assign n25230 = ~n25301;
  assign n25302 = n25323 ^ n25324;
  assign n25325 = ~n25323;
  assign n25304 = ~n25347;
  assign n25327 = n216 ^ n25357;
  assign n25189 = ~n24040;
  assign n25164 = n25205 & n25206;
  assign n25218 = n21595 & n25219;
  assign n24103 = ~n25220;
  assign n25210 = n25223 & n25224;
  assign n25158 = n24057 ^ n24010;
  assign n25225 = ~n25242;
  assign n25246 = n25270 & n25271;
  assign n25248 = ~n25297;
  assign n25274 = n217 ^ n25302;
  assign n25319 = n25325 & n25326;
  assign n25276 = n25327 ^ n25328;
  assign n25207 = n25210 & n1507;
  assign n24085 = ~n25218;
  assign n25201 = ~n25210;
  assign n25211 = n25225 & n25226;
  assign n25228 = n25246 ^ n22779;
  assign n25247 = ~n25246;
  assign n25197 = n25273 ^ n25274;
  assign n25256 = n25274 & n25273;
  assign n25303 = ~n25319;
  assign n25187 = n25201 ^ n25192;
  assign n25202 = n25201 & n310;
  assign n25191 = ~n25207;
  assign n25193 = n25211 ^ n25212;
  assign n25213 = ~n25211;
  assign n21515 = n25227 ^ n25228;
  assign n25243 = n25247 & n25248;
  assign n25255 = n25197 & n22849;
  assign n25254 = ~n25197;
  assign n25275 = n25303 & n25304;
  assign n25165 = n310 ^ n25187;
  assign n25186 = n21515 & n25189;
  assign n25190 = n25191 & n25192;
  assign n25154 = n25193 ^ n25194;
  assign n25174 = ~n25202;
  assign n25208 = n25213 & n25214;
  assign n21523 = ~n21515;
  assign n25229 = ~n25243;
  assign n25249 = n25254 & n22760;
  assign n25200 = ~n25255;
  assign n25257 = n25275 ^ n25276;
  assign n24000 = n25164 ^ n25165;
  assign n25117 = n25165 & n25164;
  assign n24062 = ~n25186;
  assign n25175 = n25154 & n1450;
  assign n25173 = ~n25190;
  assign n25176 = ~n25154;
  assign n25188 = n21523 & n24040;
  assign n25195 = ~n25208;
  assign n24016 = n21523 ^ n22779;
  assign n25215 = n25229 & n25230;
  assign n25217 = ~n25249;
  assign n25160 = n25256 ^ n25257;
  assign n25147 = ~n24000;
  assign n25120 = ~n25117;
  assign n25153 = n25173 & n25174;
  assign n25156 = ~n25175;
  assign n25168 = n25176 & n309;
  assign n24043 = ~n25188;
  assign n25110 = n24008 ^ n24016;
  assign n25177 = n25195 & n25196;
  assign n25198 = n25215 ^ n22760;
  assign n25216 = ~n25215;
  assign n25236 = n25160 & n22802;
  assign n25235 = ~n25160;
  assign n25137 = n25153 ^ n25154;
  assign n25155 = ~n25153;
  assign n25139 = ~n25168;
  assign n25157 = n25177 ^ n25178;
  assign n25171 = n25110 & n25182;
  assign n25181 = n25177 & n25178;
  assign n25170 = ~n25110;
  assign n25179 = ~n25177;
  assign n21461 = n25197 ^ n25198;
  assign n25209 = n25216 & n25217;
  assign n25231 = n25235 & n22677;
  assign n25185 = ~n25236;
  assign n25118 = n309 ^ n25137;
  assign n25148 = n21461 & n24000;
  assign n25152 = n25155 & n25156;
  assign n25122 = n25157 ^ n25158;
  assign n25167 = n25170 & n25129;
  assign n25112 = ~n25171;
  assign n25169 = n25179 & n25180;
  assign n25166 = ~n25181;
  assign n23976 = n21461 ^ n22760;
  assign n21446 = ~n21461;
  assign n25199 = ~n25209;
  assign n25163 = ~n25231;
  assign n25108 = n25117 ^ n25118;
  assign n25119 = ~n25118;
  assign n25136 = n21446 & n25147;
  assign n24002 = ~n25148;
  assign n25141 = n25122 & n308;
  assign n25138 = ~n25152;
  assign n25140 = ~n25122;
  assign n25071 = n23976 ^ n23968;
  assign n25159 = n25166 & n25158;
  assign n25131 = ~n25167;
  assign n25150 = ~n25169;
  assign n25183 = n25199 & n25200;
  assign n25104 = ~n25108;
  assign n25078 = n25119 & n25120;
  assign n24021 = ~n25136;
  assign n25121 = n25138 & n25139;
  assign n25133 = n25140 & n1423;
  assign n25107 = ~n25141;
  assign n25142 = n25071 & n25088;
  assign n25143 = ~n25071;
  assign n25149 = ~n25159;
  assign n25161 = n25183 ^ n22802;
  assign n25184 = ~n25183;
  assign n25081 = ~n25078;
  assign n25105 = n25121 ^ n25122;
  assign n25123 = ~n25121;
  assign n25124 = ~n25133;
  assign n25074 = ~n25142;
  assign n25134 = n25143 & n25144;
  assign n25128 = n25149 & n25150;
  assign n21289 = n25160 ^ n25161;
  assign n25172 = n25184 & n25185;
  assign n25079 = n308 ^ n25105;
  assign n25103 = n21289 & n25108;
  assign n25115 = n25123 & n25124;
  assign n25109 = n25128 ^ n25129;
  assign n25090 = ~n25134;
  assign n25130 = ~n25128;
  assign n21337 = ~n21289;
  assign n25162 = ~n25172;
  assign n25068 = n25078 ^ n25079;
  assign n25080 = ~n25079;
  assign n23981 = ~n25103;
  assign n25096 = n21337 & n25104;
  assign n25077 = n25109 ^ n25110;
  assign n25106 = ~n25115;
  assign n25125 = n25130 & n25131;
  assign n23953 = n21337 ^ n22677;
  assign n25151 = n25162 & n25163;
  assign n25065 = ~n25068;
  assign n25040 = n25080 & n25081;
  assign n23962 = ~n25096;
  assign n25086 = n25077 & n307;
  assign n25097 = n25106 & n25107;
  assign n25085 = ~n25077;
  assign n25031 = n23953 ^ n23937;
  assign n25111 = ~n25125;
  assign n25146 = n25151 & n22717;
  assign n25145 = ~n25151;
  assign n25043 = ~n25040;
  assign n23978 = n23981 & n23962;
  assign n25082 = n25085 & n1356;
  assign n25052 = ~n25086;
  assign n25070 = ~n25097;
  assign n25098 = n25031 & n25056;
  assign n25087 = n25111 & n25112;
  assign n25099 = ~n25031;
  assign n25135 = n25145 & n22729;
  assign n25127 = ~n25146;
  assign n25064 = n25070 ^ n25077;
  assign n25069 = ~n25082;
  assign n25072 = n25087 ^ n25088;
  assign n25033 = ~n25098;
  assign n25091 = n25099 & n25100;
  assign n25089 = ~n25087;
  assign n25126 = n25127 & n25132;
  assign n25114 = ~n25135;
  assign n25041 = n307 ^ n25064;
  assign n25067 = n25069 & n25070;
  assign n25027 = n25071 ^ n25072;
  assign n25083 = n25089 & n25090;
  assign n25058 = ~n25091;
  assign n25113 = ~n25126;
  assign n25116 = n25114 & n25127;
  assign n23896 = n25040 ^ n25041;
  assign n25042 = ~n25041;
  assign n25053 = n25027 & n1286;
  assign n25051 = ~n25067;
  assign n25054 = ~n25027;
  assign n25073 = ~n25083;
  assign n25092 = n25113 & n25114;
  assign n25101 = ~n25116;
  assign n25022 = ~n23896;
  assign n24988 = n25042 & n25043;
  assign n25026 = n25051 & n25052;
  assign n25028 = ~n25053;
  assign n25047 = n25054 & n306;
  assign n25055 = n25073 & n25074;
  assign n21083 = n25092 ^ n25093;
  assign n21272 = n25101 ^ n25102;
  assign n25094 = ~n25092;
  assign n25005 = n21083 & n25022;
  assign n25000 = ~n24988;
  assign n25006 = n25026 ^ n25027;
  assign n25029 = ~n25026;
  assign n25008 = ~n25047;
  assign n25030 = n25055 ^ n25056;
  assign n25057 = ~n25055;
  assign n25066 = n21272 & n25068;
  assign n23857 = n22671 ^ n21083;
  assign n23913 = n22729 ^ n21272;
  assign n21231 = ~n21083;
  assign n25084 = n25094 & n25095;
  assign n21204 = ~n21272;
  assign n23877 = ~n25005;
  assign n24989 = n306 ^ n25006;
  assign n25021 = n21231 & n23896;
  assign n25024 = n25028 & n25029;
  assign n24991 = n25030 ^ n25031;
  assign n25048 = n25057 & n25058;
  assign n24978 = n23857 ^ n23788;
  assign n24995 = n23913 ^ n23909;
  assign n25063 = n21204 & n25065;
  assign n23917 = ~n25066;
  assign n25075 = ~n25084;
  assign n23861 = n24988 ^ n24989;
  assign n24949 = n24989 & n25000;
  assign n23898 = ~n25021;
  assign n25009 = n24991 & n1201;
  assign n25007 = ~n25024;
  assign n25010 = ~n24991;
  assign n25035 = n24978 & n25044;
  assign n25032 = ~n25048;
  assign n25046 = n24995 & n25049;
  assign n25034 = ~n24978;
  assign n25045 = ~n24995;
  assign n23941 = ~n25063;
  assign n25059 = n25075 & n25076;
  assign n24971 = ~n23861;
  assign n24952 = ~n24949;
  assign n24990 = n25007 & n25008;
  assign n24992 = ~n25009;
  assign n25001 = n25010 & n305;
  assign n25011 = n25032 & n25033;
  assign n25025 = n25034 & n24958;
  assign n24980 = ~n25035;
  assign n25036 = n25045 & n25012;
  assign n24997 = ~n25046;
  assign n25039 = n23941 & n23917;
  assign n23817 = n25059 ^ n25060;
  assign n25061 = ~n25059;
  assign n24972 = n24990 ^ n24991;
  assign n24993 = ~n24990;
  assign n24974 = ~n25001;
  assign n24994 = n25011 ^ n25012;
  assign n25013 = ~n25011;
  assign n24960 = ~n25025;
  assign n25014 = ~n25036;
  assign n24941 = n23796 ^ n23817;
  assign n20996 = n22474 ^ n23817;
  assign n23939 = ~n25039;
  assign n25050 = n25061 & n25062;
  assign n24965 = n20996 & n24971;
  assign n24950 = n305 ^ n24972;
  assign n24987 = n24992 & n24993;
  assign n24954 = n24994 ^ n24995;
  assign n25002 = n25013 & n25014;
  assign n25016 = n24941 & n25023;
  assign n25015 = ~n24941;
  assign n21147 = ~n20996;
  assign n25037 = ~n25050;
  assign n23821 = n24949 ^ n24950;
  assign n23843 = ~n24965;
  assign n24951 = ~n24950;
  assign n24970 = n21147 & n23861;
  assign n24976 = n24954 & n304;
  assign n24973 = ~n24987;
  assign n24975 = ~n24954;
  assign n24996 = ~n25002;
  assign n25003 = n25015 & n24924;
  assign n24943 = ~n25016;
  assign n25017 = n25037 & n25038;
  assign n24934 = ~n23821;
  assign n24918 = n24951 & n24952;
  assign n23863 = ~n24970;
  assign n24953 = n24973 & n24974;
  assign n24966 = n24975 & n1168;
  assign n24937 = ~n24976;
  assign n24977 = n24996 & n24997;
  assign n24926 = ~n25003;
  assign n23771 = n25017 ^ n25018;
  assign n25019 = ~n25017;
  assign n24935 = n24953 ^ n24954;
  assign n24955 = ~n24953;
  assign n24956 = ~n24966;
  assign n24957 = n24977 ^ n24978;
  assign n24979 = ~n24977;
  assign n24904 = n23771 ^ n23743;
  assign n20913 = n23771 ^ n22468;
  assign n25004 = n25019 & n25020;
  assign n24929 = n20913 & n24934;
  assign n24919 = n304 ^ n24935;
  assign n24948 = n24955 & n24956;
  assign n24898 = n24957 ^ n24958;
  assign n24967 = n24979 & n24980;
  assign n24983 = n24904 & n24882;
  assign n24981 = ~n24904;
  assign n21055 = ~n20913;
  assign n24998 = ~n25004;
  assign n24915 = n24918 ^ n24919;
  assign n24875 = n24919 & n24918;
  assign n23801 = ~n24929;
  assign n24933 = n21055 & n23821;
  assign n24939 = n24898 & n319;
  assign n24936 = ~n24948;
  assign n24938 = ~n24898;
  assign n24959 = ~n24967;
  assign n24968 = n24981 & n24982;
  assign n24906 = ~n24983;
  assign n24984 = n24998 & n24999;
  assign n24896 = ~n24915;
  assign n23823 = ~n24933;
  assign n24920 = n24936 & n24937;
  assign n24930 = n24938 & n1118;
  assign n24900 = ~n24939;
  assign n24940 = n24959 & n24960;
  assign n24884 = ~n24968;
  assign n24962 = n24984 ^ n22334;
  assign n24985 = ~n24984;
  assign n24897 = n319 ^ n24920;
  assign n24921 = ~n24920;
  assign n24922 = ~n24930;
  assign n24923 = n24940 ^ n24941;
  assign n24942 = ~n24940;
  assign n20962 = n24961 ^ n24962;
  assign n24969 = n24985 & n24986;
  assign n24889 = n20962 & n24896;
  assign n24876 = n24897 ^ n24898;
  assign n24917 = n24921 & n24922;
  assign n24878 = n24923 ^ n24924;
  assign n24931 = n24942 & n24943;
  assign n23745 = n20962 ^ n22469;
  assign n20869 = ~n20962;
  assign n24963 = ~n24969;
  assign n24872 = n24875 ^ n24876;
  assign n24839 = n24876 & n24875;
  assign n23749 = ~n24889;
  assign n24895 = n20869 & n24915;
  assign n24902 = n24878 & n318;
  assign n24899 = ~n24917;
  assign n24901 = ~n24878;
  assign n24848 = n23745 ^ n23734;
  assign n24925 = ~n24931;
  assign n24944 = n24963 & n24964;
  assign n24858 = ~n24872;
  assign n24842 = ~n24839;
  assign n23776 = ~n24895;
  assign n24877 = n24899 & n24900;
  assign n24890 = n24901 & n1025;
  assign n24861 = ~n24902;
  assign n24909 = n24848 & n24865;
  assign n24907 = ~n24848;
  assign n24903 = n24925 & n24926;
  assign n23693 = n24944 ^ n24945;
  assign n24946 = ~n24944;
  assign n24873 = n23776 & n23749;
  assign n24859 = n24877 ^ n24878;
  assign n24879 = ~n24877;
  assign n24880 = ~n24890;
  assign n24881 = n24903 ^ n24904;
  assign n24892 = n24907 & n24908;
  assign n24850 = ~n24909;
  assign n24905 = ~n24903;
  assign n24810 = n23693 ^ n23686;
  assign n20787 = n22384 ^ n23693;
  assign n24932 = n24946 & n24947;
  assign n24853 = n20787 & n24858;
  assign n24840 = n318 ^ n24859;
  assign n23774 = ~n24873;
  assign n24874 = n24879 & n24880;
  assign n24844 = n24881 ^ n24882;
  assign n24867 = ~n24892;
  assign n24891 = n24905 & n24906;
  assign n24910 = n24810 & n24916;
  assign n24911 = ~n24810;
  assign n20885 = ~n20787;
  assign n24927 = ~n24932;
  assign n23644 = n24839 ^ n24840;
  assign n23697 = ~n24853;
  assign n24841 = ~n24840;
  assign n24857 = n20885 & n24872;
  assign n24862 = n24844 & n970;
  assign n24860 = ~n24874;
  assign n24863 = ~n24844;
  assign n24883 = ~n24891;
  assign n24812 = ~n24910;
  assign n24893 = n24911 & n24828;
  assign n24912 = n24927 & n24928;
  assign n24821 = ~n23644;
  assign n24803 = n24841 & n24842;
  assign n23725 = ~n24857;
  assign n24843 = n24860 & n24861;
  assign n24846 = ~n24862;
  assign n24854 = n24863 & n317;
  assign n24864 = n24883 & n24884;
  assign n24830 = ~n24893;
  assign n24885 = n24912 ^ n22271;
  assign n24913 = ~n24912;
  assign n24837 = n23725 & n23697;
  assign n24822 = n24843 ^ n24844;
  assign n24845 = ~n24843;
  assign n24824 = ~n24854;
  assign n24847 = n24864 ^ n24865;
  assign n24866 = ~n24864;
  assign n20692 = n24885 ^ n24886;
  assign n24894 = n24913 & n24914;
  assign n24814 = n20692 & n24821;
  assign n24804 = n317 ^ n24822;
  assign n23723 = ~n24837;
  assign n24838 = n24845 & n24846;
  assign n24806 = n24847 ^ n24848;
  assign n24855 = n24866 & n24867;
  assign n20799 = ~n20692;
  assign n24887 = ~n24894;
  assign n24800 = n24803 ^ n24804;
  assign n24801 = n24804 & n24803;
  assign n23673 = ~n24814;
  assign n24820 = n20799 & n23644;
  assign n24825 = n24806 & n901;
  assign n24823 = ~n24838;
  assign n24826 = ~n24806;
  assign n24849 = ~n24855;
  assign n23613 = n20799 ^ n22271;
  assign n24868 = n24887 & n24888;
  assign n24788 = ~n24800;
  assign n24774 = ~n24801;
  assign n23647 = ~n24820;
  assign n24805 = n24823 & n24824;
  assign n24807 = ~n24825;
  assign n24815 = n24826 & n316;
  assign n24780 = n23613 ^ n23541;
  assign n24827 = n24849 & n24850;
  assign n23585 = n24868 ^ n24869;
  assign n24870 = ~n24868;
  assign n24789 = n24805 ^ n24806;
  assign n24808 = ~n24805;
  assign n24791 = ~n24815;
  assign n24809 = n24827 ^ n24828;
  assign n24818 = n24780 & n24831;
  assign n24817 = ~n24780;
  assign n24829 = ~n24827;
  assign n24755 = n23585 ^ n23485;
  assign n20722 = n23585 ^ n22228;
  assign n24856 = n24870 & n24871;
  assign n24772 = n316 ^ n24789;
  assign n24787 = n20722 & n24800;
  assign n24802 = n24807 & n24808;
  assign n24776 = n24809 ^ n24810;
  assign n24813 = n24817 & n24795;
  assign n24782 = ~n24818;
  assign n24816 = n24829 & n24830;
  assign n24832 = n24755 & n24836;
  assign n24833 = ~n24755;
  assign n20626 = ~n20722;
  assign n24851 = ~n24856;
  assign n24773 = ~n24772;
  assign n23589 = ~n24787;
  assign n24784 = n20626 & n24788;
  assign n24793 = n24776 & n315;
  assign n24790 = ~n24802;
  assign n24792 = ~n24776;
  assign n24797 = ~n24813;
  assign n24811 = ~n24816;
  assign n24757 = ~n24832;
  assign n24819 = n24833 & n24766;
  assign n24834 = n24851 & n24852;
  assign n24748 = n24773 & n24774;
  assign n23618 = ~n24784;
  assign n24775 = n24790 & n24791;
  assign n24785 = n24792 & n840;
  assign n24762 = ~n24793;
  assign n24794 = n24811 & n24812;
  assign n24768 = ~n24819;
  assign n22141 = n24834 ^ n24835;
  assign n24769 = n23618 & n23589;
  assign n24760 = n24775 ^ n24776;
  assign n24777 = ~n24775;
  assign n24778 = ~n24785;
  assign n24779 = n24794 ^ n24795;
  assign n24771 = n24801 ^ n22141;
  assign n24796 = ~n24794;
  assign n24798 = n22141 ^ n22106;
  assign n24749 = n315 ^ n24760;
  assign n23616 = ~n24769;
  assign n23558 = n24771 ^ n24772;
  assign n24770 = n24777 & n24778;
  assign n24751 = n24779 ^ n24780;
  assign n24786 = n24796 & n24797;
  assign n23525 = n24798 ^ n24799;
  assign n22833 = n24748 ^ n24749;
  assign n24729 = n24749 & n24748;
  assign n24764 = n24751 & n314;
  assign n24761 = ~n24770;
  assign n24763 = ~n24751;
  assign n24738 = n23525 ^ n24783;
  assign n24781 = ~n24786;
  assign n24726 = n24740 ^ n22833;
  assign n23778 = ~n22833;
  assign n24732 = ~n24729;
  assign n24750 = n24761 & n24762;
  assign n24758 = n24763 & n792;
  assign n24743 = ~n24764;
  assign n24765 = n24781 & n24782;
  assign n23241 = n391 ^ n24726;
  assign n24662 = n24726 & n391;
  assign n21843 = n22814 ^ n23778;
  assign n24727 = n23792 ^ n23778;
  assign n24701 = n23778 & n22814;
  assign n24741 = n24750 ^ n24751;
  assign n24752 = ~n24750;
  assign n24753 = ~n24758;
  assign n24754 = n24765 ^ n24766;
  assign n24767 = ~n24765;
  assign n24723 = n24662 & n390;
  assign n24393 = ~n23241;
  assign n24682 = n24727 & n24728;
  assign n24722 = ~n24662;
  assign n24730 = n314 ^ n24741;
  assign n24747 = n24752 & n24753;
  assign n24734 = n24754 ^ n24755;
  assign n24759 = n24767 & n24768;
  assign n24713 = n24722 & n16646;
  assign n24716 = n24682 & n24675;
  assign n24656 = ~n24723;
  assign n24714 = ~n24682;
  assign n24724 = n24729 ^ n24730;
  assign n24731 = ~n24730;
  assign n24745 = n24734 & n313;
  assign n24742 = ~n24747;
  assign n24744 = ~n24734;
  assign n24756 = ~n24759;
  assign n24669 = ~n24713;
  assign n24711 = n24714 & n24715;
  assign n24679 = ~n24716;
  assign n24717 = n24724 & n22698;
  assign n24718 = ~n24724;
  assign n24708 = n24731 & n24732;
  assign n24733 = n24742 & n24743;
  assign n24739 = n24744 & n746;
  assign n24721 = ~n24745;
  assign n24746 = n24756 & n24757;
  assign n24689 = ~n24711;
  assign n24703 = ~n24717;
  assign n24712 = n24718 & n22689;
  assign n24710 = ~n24708;
  assign n24719 = n24733 ^ n24734;
  assign n24735 = ~n24733;
  assign n24736 = ~n24739;
  assign n24737 = n312 ^ n24746;
  assign n24707 = ~n24712;
  assign n24709 = n313 ^ n24719;
  assign n24725 = n24735 & n24736;
  assign n24699 = n24737 ^ n24738;
  assign n24706 = n24707 & n24701;
  assign n24700 = n24707 & n24703;
  assign n24686 = n24708 ^ n24709;
  assign n24705 = n24709 & n24710;
  assign n24720 = ~n24725;
  assign n21753 = n24700 ^ n24701;
  assign n24702 = ~n24706;
  assign n24704 = n24720 & n24721;
  assign n24683 = n24694 ^ n21753;
  assign n21819 = ~n21753;
  assign n24695 = n24702 & n24703;
  assign n24698 = n24704 ^ n24705;
  assign n24674 = n24682 ^ n24683;
  assign n24684 = n24683 & n24689;
  assign n24685 = n24695 ^ n22628;
  assign n24658 = n24698 ^ n24699;
  assign n24697 = n24695 & n22628;
  assign n24696 = ~n24695;
  assign n24663 = n24674 ^ n24675;
  assign n24678 = ~n24684;
  assign n21738 = n24685 ^ n24686;
  assign n24690 = n24658 & n22488;
  assign n24691 = ~n24658;
  assign n24693 = n24696 & n22589;
  assign n24692 = ~n24697;
  assign n24650 = n24662 ^ n24663;
  assign n24664 = n24663 & n24669;
  assign n24652 = n24676 ^ n21738;
  assign n24677 = n24678 & n24679;
  assign n21736 = ~n21738;
  assign n24660 = ~n24690;
  assign n24687 = n24691 & n22577;
  assign n24688 = n24692 & n24686;
  assign n24681 = ~n24693;
  assign n24637 = n390 ^ n24650;
  assign n24655 = ~n24664;
  assign n24667 = n24652 & n24670;
  assign n24665 = ~n24652;
  assign n24654 = ~n24677;
  assign n24673 = ~n24687;
  assign n24680 = ~n24688;
  assign n23189 = n24637 ^ n23241;
  assign n24609 = n24637 & n23241;
  assign n24638 = n24655 & n24656;
  assign n24661 = n24665 & n24666;
  assign n24643 = ~n24667;
  assign n24651 = n24654 ^ n24666;
  assign n24671 = n24680 & n24681;
  assign n24340 = ~n23189;
  assign n24612 = ~n24609;
  assign n24628 = ~n24638;
  assign n24639 = n24651 ^ n24652;
  assign n24653 = ~n24661;
  assign n24657 = n24671 ^ n22577;
  assign n24672 = ~n24671;
  assign n24623 = n24638 ^ n24639;
  assign n24640 = n24639 & n16551;
  assign n24641 = ~n24639;
  assign n24648 = n24653 & n24654;
  assign n21591 = n24657 ^ n24658;
  assign n24668 = n24672 & n24673;
  assign n24610 = n389 ^ n24623;
  assign n24627 = ~n24640;
  assign n24634 = n24641 & n389;
  assign n24604 = n24645 ^ n21591;
  assign n24642 = ~n24648;
  assign n21577 = ~n21591;
  assign n24659 = ~n24668;
  assign n24301 = n24609 ^ n24610;
  assign n24611 = ~n24610;
  assign n24624 = n24627 & n24628;
  assign n24631 = n24604 & n24620;
  assign n24617 = ~n24634;
  assign n24635 = n24642 & n24643;
  assign n24629 = ~n24604;
  assign n24649 = n24659 & n24660;
  assign n24317 = ~n24301;
  assign n24558 = n24611 & n24612;
  assign n24616 = ~n24624;
  assign n24625 = n24629 & n24630;
  assign n24602 = ~n24631;
  assign n24619 = ~n24635;
  assign n24647 = n24649 & n22493;
  assign n24646 = ~n24649;
  assign n24561 = ~n24558;
  assign n24592 = n24616 & n24617;
  assign n24605 = n24619 ^ n24620;
  assign n24618 = ~n24625;
  assign n24644 = n24646 & n22455;
  assign n24633 = ~n24647;
  assign n24593 = n24604 ^ n24605;
  assign n24580 = ~n24592;
  assign n24613 = n24618 & n24619;
  assign n24632 = n24633 & n24636;
  assign n24622 = ~n24644;
  assign n24578 = n24592 ^ n24593;
  assign n24595 = n24593 & n388;
  assign n24594 = ~n24593;
  assign n24601 = ~n24613;
  assign n24621 = ~n24632;
  assign n24626 = n24622 & n24633;
  assign n24559 = n388 ^ n24578;
  assign n24589 = n24594 & n16413;
  assign n24563 = ~n24595;
  assign n24590 = n24601 & n24602;
  assign n24606 = n24621 & n24622;
  assign n24614 = ~n24626;
  assign n24275 = n24558 ^ n24559;
  assign n24560 = ~n24559;
  assign n24579 = ~n24589;
  assign n24574 = n24590 ^ n24588;
  assign n24573 = ~n24590;
  assign n24596 = n24606 ^ n22403;
  assign n21533 = n24614 ^ n24615;
  assign n24607 = ~n24606;
  assign n24259 = ~n24275;
  assign n24514 = n24560 & n24561;
  assign n24576 = n24579 & n24580;
  assign n21471 = n24596 ^ n24597;
  assign n24575 = n24600 ^ n21533;
  assign n24603 = n24607 & n24608;
  assign n21486 = ~n21533;
  assign n24546 = n24574 ^ n24575;
  assign n24562 = ~n24576;
  assign n24520 = n24581 ^ n21471;
  assign n24586 = n24575 & n24591;
  assign n21453 = ~n21471;
  assign n24587 = ~n24575;
  assign n24598 = ~n24603;
  assign n24556 = n24546 & n387;
  assign n24545 = n24562 & n24563;
  assign n24555 = ~n24546;
  assign n24564 = n24520 & n24536;
  assign n24565 = ~n24520;
  assign n24554 = ~n24586;
  assign n24582 = n24587 & n24588;
  assign n24583 = n24598 & n24599;
  assign n24529 = n24545 ^ n24546;
  assign n24552 = n24555 & n16311;
  assign n24527 = ~n24556;
  assign n24543 = ~n24545;
  assign n24525 = ~n24564;
  assign n24557 = n24565 & n24566;
  assign n24572 = ~n24582;
  assign n24567 = n24583 ^ n22285;
  assign n24584 = ~n24583;
  assign n24515 = n387 ^ n24529;
  assign n24542 = ~n24552;
  assign n24541 = ~n24557;
  assign n21318 = n24567 ^ n24568;
  assign n24569 = n24572 & n24573;
  assign n24577 = n24584 & n24585;
  assign n23102 = n24514 ^ n24515;
  assign n24516 = ~n24515;
  assign n24539 = n24542 & n24543;
  assign n24491 = n24547 ^ n21318;
  assign n21390 = ~n21318;
  assign n24553 = ~n24569;
  assign n24570 = ~n24577;
  assign n24234 = ~n23102;
  assign n24463 = n24516 & n24514;
  assign n24526 = ~n24539;
  assign n24530 = n24491 & n24540;
  assign n24531 = ~n24491;
  assign n24548 = n24553 & n24554;
  assign n24549 = n24570 & n24571;
  assign n24466 = ~n24463;
  assign n24517 = n24526 & n24527;
  assign n24493 = ~n24530;
  assign n24528 = n24531 & n24509;
  assign n24535 = ~n24548;
  assign n24534 = n24549 ^ n22209;
  assign n24550 = ~n24549;
  assign n24512 = n24517 & n16246;
  assign n24498 = ~n24517;
  assign n24511 = ~n24528;
  assign n21210 = n24533 ^ n24534;
  assign n24519 = n24535 ^ n24536;
  assign n24532 = n24541 & n24535;
  assign n24544 = n24550 & n24551;
  assign n24506 = n24498 & n386;
  assign n24496 = ~n24512;
  assign n24457 = n24518 ^ n21210;
  assign n24497 = n24519 ^ n24520;
  assign n21341 = ~n21210;
  assign n24524 = ~n24532;
  assign n24537 = ~n24544;
  assign n24494 = n24496 & n24497;
  assign n24484 = n24498 ^ n24497;
  assign n24486 = ~n24506;
  assign n24500 = n24457 & n24507;
  assign n24499 = ~n24457;
  assign n24508 = n24524 & n24525;
  assign n24521 = n24537 & n24538;
  assign n24464 = n386 ^ n24484;
  assign n24485 = ~n24494;
  assign n24495 = n24499 & n24479;
  assign n24459 = ~n24500;
  assign n24490 = n24508 ^ n24509;
  assign n24510 = ~n24508;
  assign n24502 = n24521 ^ n22196;
  assign n24522 = ~n24521;
  assign n24194 = n24463 ^ n24464;
  assign n24465 = ~n24464;
  assign n24467 = n24485 & n24486;
  assign n24468 = n24490 ^ n24491;
  assign n24480 = ~n24495;
  assign n21171 = n24502 ^ n24503;
  assign n24501 = n24510 & n24511;
  assign n24513 = n24522 & n24523;
  assign n24179 = ~n24194;
  assign n24428 = n24465 & n24466;
  assign n24448 = n24467 ^ n24468;
  assign n24455 = ~n24467;
  assign n24477 = n24468 & n385;
  assign n24476 = ~n24468;
  assign n21226 = ~n21171;
  assign n24492 = ~n24501;
  assign n24504 = ~n24513;
  assign n24429 = n385 ^ n24448;
  assign n24469 = n24476 & n16138;
  assign n24439 = ~n24477;
  assign n24424 = n24482 ^ n21226;
  assign n24478 = n24492 & n24493;
  assign n24487 = n24504 & n24505;
  assign n24154 = n24428 ^ n24429;
  assign n24383 = n24429 & n24428;
  assign n24454 = ~n24469;
  assign n24462 = n24424 & n24470;
  assign n24456 = n24478 ^ n24479;
  assign n24461 = ~n24424;
  assign n24481 = ~n24478;
  assign n24473 = n24487 ^ n22127;
  assign n24488 = ~n24487;
  assign n23006 = ~n24154;
  assign n24449 = n24454 & n24455;
  assign n24420 = n24456 ^ n24457;
  assign n24460 = n24461 & n24444;
  assign n24426 = ~n24462;
  assign n21089 = n24472 ^ n24473;
  assign n24471 = n24480 & n24481;
  assign n24483 = n24488 & n24489;
  assign n24441 = n24420 & n384;
  assign n24438 = ~n24449;
  assign n24440 = ~n24420;
  assign n24390 = n24450 ^ n21089;
  assign n24446 = ~n24460;
  assign n21176 = ~n21089;
  assign n24458 = ~n24471;
  assign n24474 = ~n24483;
  assign n24419 = n24438 & n24439;
  assign n24430 = n24440 & n16072;
  assign n24405 = ~n24441;
  assign n24432 = n24390 & n24442;
  assign n24431 = ~n24390;
  assign n24443 = n24458 & n24459;
  assign n24451 = n24474 & n24475;
  assign n24403 = n24419 ^ n24420;
  assign n24422 = ~n24419;
  assign n24421 = ~n24430;
  assign n24427 = n24431 & n24410;
  assign n24392 = ~n24432;
  assign n24423 = n24443 ^ n24444;
  assign n24445 = ~n24443;
  assign n24434 = n24451 ^ n22054;
  assign n24452 = ~n24451;
  assign n24384 = n384 ^ n24403;
  assign n24414 = n24421 & n24422;
  assign n24386 = n24423 ^ n24424;
  assign n24412 = ~n24427;
  assign n21074 = n24434 ^ n24435;
  assign n24433 = n24445 & n24446;
  assign n24447 = n24452 & n24453;
  assign n24114 = n24383 ^ n24384;
  assign n24346 = n24384 & n24383;
  assign n24407 = n24386 & n399;
  assign n24404 = ~n24414;
  assign n24406 = ~n24386;
  assign n24353 = n24415 ^ n21074;
  assign n21004 = ~n21074;
  assign n24425 = ~n24433;
  assign n24436 = ~n24447;
  assign n24099 = ~n24114;
  assign n24385 = n24404 & n24405;
  assign n24395 = n24406 & n15958;
  assign n24368 = ~n24407;
  assign n24397 = n24353 & n24408;
  assign n24396 = ~n24353;
  assign n24409 = n24425 & n24426;
  assign n24416 = n24436 & n24437;
  assign n24366 = n24385 ^ n24386;
  assign n24388 = ~n24385;
  assign n24387 = ~n24395;
  assign n24394 = n24396 & n24372;
  assign n24355 = ~n24397;
  assign n24389 = n24409 ^ n24410;
  assign n24411 = ~n24409;
  assign n24399 = n24416 ^ n21971;
  assign n24417 = ~n24416;
  assign n24347 = n399 ^ n24366;
  assign n24377 = n24387 & n24388;
  assign n24349 = n24389 ^ n24390;
  assign n24374 = ~n24394;
  assign n20878 = n24399 ^ n24400;
  assign n24398 = n24411 & n24412;
  assign n24413 = n24417 & n24418;
  assign n24059 = n24346 ^ n24347;
  assign n24305 = n24347 & n24346;
  assign n24370 = n24349 & n398;
  assign n24367 = ~n24377;
  assign n24369 = ~n24349;
  assign n24314 = n24378 ^ n20878;
  assign n24379 = n20878 & n24393;
  assign n21015 = ~n20878;
  assign n24391 = ~n24398;
  assign n24401 = ~n24413;
  assign n24074 = ~n24059;
  assign n24308 = ~n24305;
  assign n24348 = n24367 & n24368;
  assign n24357 = n24369 & n15897;
  assign n24328 = ~n24370;
  assign n24360 = n24314 & n24333;
  assign n24358 = ~n24314;
  assign n24375 = n21015 & n23241;
  assign n23223 = ~n24379;
  assign n24371 = n24391 & n24392;
  assign n24380 = n24401 & n24402;
  assign n24326 = n24348 ^ n24349;
  assign n24351 = ~n24348;
  assign n24350 = ~n24357;
  assign n24356 = n24358 & n24359;
  assign n24316 = ~n24360;
  assign n24352 = n24371 ^ n24372;
  assign n23243 = ~n24375;
  assign n24373 = ~n24371;
  assign n24362 = n24380 ^ n21938;
  assign n24381 = ~n24380;
  assign n24306 = n398 ^ n24326;
  assign n24338 = n24350 & n24351;
  assign n24310 = n24352 ^ n24353;
  assign n24335 = ~n24356;
  assign n20938 = n24362 ^ n24363;
  assign n24361 = n24373 & n24374;
  assign n24376 = n24381 & n24382;
  assign n24032 = n24305 ^ n24306;
  assign n24307 = ~n24306;
  assign n24330 = n24310 & n397;
  assign n24327 = ~n24338;
  assign n24329 = ~n24310;
  assign n24272 = n24339 ^ n20938;
  assign n24341 = n20938 & n23189;
  assign n20928 = ~n20938;
  assign n24354 = ~n24361;
  assign n24364 = ~n24376;
  assign n24018 = ~n24032;
  assign n24264 = n24307 & n24308;
  assign n24309 = n24327 & n24328;
  assign n24319 = n24329 & n15813;
  assign n24288 = ~n24330;
  assign n24320 = n24272 & n24331;
  assign n24321 = ~n24272;
  assign n24336 = n20928 & n24340;
  assign n23191 = ~n24341;
  assign n24332 = n24354 & n24355;
  assign n24342 = n24364 & n24365;
  assign n24286 = n24309 ^ n24310;
  assign n24311 = ~n24309;
  assign n24312 = ~n24319;
  assign n24274 = ~n24320;
  assign n24318 = n24321 & n24293;
  assign n24313 = n24332 ^ n24333;
  assign n23206 = ~n24336;
  assign n24334 = ~n24332;
  assign n24323 = n24342 ^ n24343;
  assign n24344 = ~n24342;
  assign n24265 = n397 ^ n24286;
  assign n24298 = n24311 & n24312;
  assign n24268 = n24313 ^ n24314;
  assign n24295 = ~n24318;
  assign n20825 = n24323 ^ n21910;
  assign n24322 = n24334 & n24335;
  assign n24337 = n24344 & n24345;
  assign n22876 = n24264 ^ n24265;
  assign n24266 = ~n24265;
  assign n24289 = n24268 & n15732;
  assign n24287 = ~n24298;
  assign n24290 = ~n24268;
  assign n24231 = n24299 ^ n20825;
  assign n24300 = n20825 & n24317;
  assign n20812 = ~n20825;
  assign n24315 = ~n24322;
  assign n24324 = ~n24337;
  assign n23992 = ~n22876;
  assign n24222 = n24266 & n24264;
  assign n24267 = n24287 & n24288;
  assign n24270 = ~n24289;
  assign n24278 = n24290 & n396;
  assign n24279 = n24231 & n24291;
  assign n24280 = ~n24231;
  assign n23157 = ~n24300;
  assign n24296 = n20812 & n24301;
  assign n24292 = n24315 & n24316;
  assign n24302 = n24324 & n24325;
  assign n24225 = ~n24222;
  assign n24245 = n24267 ^ n24268;
  assign n24269 = ~n24267;
  assign n24247 = ~n24278;
  assign n24233 = ~n24279;
  assign n24276 = n24280 & n24251;
  assign n24271 = n24292 ^ n24293;
  assign n23173 = ~n24296;
  assign n24294 = ~n24292;
  assign n24282 = n24302 ^ n21860;
  assign n24303 = ~n24302;
  assign n24223 = n396 ^ n24245;
  assign n24256 = n24269 & n24270;
  assign n24227 = n24271 ^ n24272;
  assign n24253 = ~n24276;
  assign n24277 = n23173 & n23157;
  assign n20749 = n24282 ^ n24283;
  assign n24281 = n24294 & n24295;
  assign n24297 = n24303 & n24304;
  assign n22839 = n24222 ^ n24223;
  assign n24224 = ~n24223;
  assign n24249 = n24227 & n395;
  assign n24246 = ~n24256;
  assign n24248 = ~n24227;
  assign n24191 = n24257 ^ n20749;
  assign n24258 = n20749 & n24275;
  assign n23171 = ~n24277;
  assign n20730 = ~n20749;
  assign n24273 = ~n24281;
  assign n24284 = ~n24297;
  assign n23959 = ~n22839;
  assign n24184 = n24224 & n24225;
  assign n24226 = n24246 & n24247;
  assign n24237 = n24248 & n15662;
  assign n24207 = ~n24249;
  assign n24240 = n24191 & n24211;
  assign n24238 = ~n24191;
  assign n23122 = ~n24258;
  assign n24254 = n20730 & n24259;
  assign n24250 = n24273 & n24274;
  assign n24260 = n24284 & n24285;
  assign n24205 = n24226 ^ n24227;
  assign n24228 = ~n24226;
  assign n24229 = ~n24237;
  assign n24235 = n24238 & n24239;
  assign n24193 = ~n24240;
  assign n24230 = n24250 ^ n24251;
  assign n23140 = ~n24254;
  assign n24252 = ~n24250;
  assign n24242 = n24260 ^ n24261;
  assign n24262 = ~n24260;
  assign n24185 = n395 ^ n24205;
  assign n24216 = n24228 & n24229;
  assign n24187 = n24230 ^ n24231;
  assign n24213 = ~n24235;
  assign n24236 = n23140 & n23122;
  assign n20562 = n24242 ^ n21803;
  assign n24241 = n24252 & n24253;
  assign n24255 = n24262 & n24263;
  assign n23914 = n24184 ^ n24185;
  assign n24142 = n24185 & n24184;
  assign n24209 = n24187 & n394;
  assign n24206 = ~n24216;
  assign n24208 = ~n24187;
  assign n24151 = n24217 ^ n20562;
  assign n24218 = n20562 & n24234;
  assign n23138 = ~n24236;
  assign n20664 = ~n20562;
  assign n24232 = ~n24241;
  assign n24243 = ~n24255;
  assign n23929 = ~n23914;
  assign n24145 = ~n24142;
  assign n24186 = n24206 & n24207;
  assign n24196 = n24208 & n15572;
  assign n24166 = ~n24209;
  assign n24199 = n24151 & n24171;
  assign n24197 = ~n24151;
  assign n24214 = n20664 & n23102;
  assign n23085 = ~n24218;
  assign n24210 = n24232 & n24233;
  assign n24219 = n24243 & n24244;
  assign n24164 = n24186 ^ n24187;
  assign n24188 = ~n24186;
  assign n24189 = ~n24196;
  assign n24195 = n24197 & n24198;
  assign n24173 = ~n24199;
  assign n24190 = n24210 ^ n24211;
  assign n23104 = ~n24214;
  assign n24212 = ~n24210;
  assign n24201 = n24219 ^ n21764;
  assign n24220 = ~n24219;
  assign n24143 = n394 ^ n24164;
  assign n24176 = n24188 & n24189;
  assign n24147 = n24190 ^ n24191;
  assign n24153 = ~n24195;
  assign n20567 = n24201 ^ n24202;
  assign n24200 = n24212 & n24213;
  assign n24215 = n24220 & n24221;
  assign n23872 = n24142 ^ n24143;
  assign n24144 = ~n24143;
  assign n24167 = n24147 & n15529;
  assign n24165 = ~n24176;
  assign n24168 = ~n24147;
  assign n24131 = n20567 ^ n24177;
  assign n24178 = n20567 & n24194;
  assign n20579 = ~n20567;
  assign n24192 = ~n24200;
  assign n24203 = ~n24215;
  assign n23859 = ~n23872;
  assign n24104 = n24144 & n24145;
  assign n24146 = n24165 & n24166;
  assign n24149 = ~n24167;
  assign n24157 = n24168 & n393;
  assign n24158 = n24131 & n24169;
  assign n24159 = ~n24131;
  assign n23065 = ~n24178;
  assign n24174 = n20579 & n24179;
  assign n24170 = n24192 & n24193;
  assign n24180 = n24203 & n24204;
  assign n24124 = n24146 ^ n24147;
  assign n24148 = ~n24146;
  assign n24126 = ~n24157;
  assign n24133 = ~n24158;
  assign n24155 = n24159 & n24111;
  assign n24150 = n24170 ^ n24171;
  assign n23045 = ~n24174;
  assign n24172 = ~n24170;
  assign n24161 = n24180 ^ n24181;
  assign n24182 = ~n24180;
  assign n24105 = n393 ^ n24124;
  assign n24136 = n24148 & n24149;
  assign n24107 = n24150 ^ n24151;
  assign n24113 = ~n24155;
  assign n24156 = n23045 & n23065;
  assign n20517 = n24161 ^ n21607;
  assign n24160 = n24172 & n24173;
  assign n24175 = n24182 & n24183;
  assign n23836 = n24104 ^ n24105;
  assign n24063 = n24105 & n24104;
  assign n24127 = n24107 & n15486;
  assign n24125 = ~n24136;
  assign n24128 = ~n24107;
  assign n24092 = n24137 ^ n20517;
  assign n24138 = n20517 & n24154;
  assign n23063 = ~n24156;
  assign n20528 = ~n20517;
  assign n24152 = ~n24160;
  assign n24162 = ~n24175;
  assign n23819 = ~n23836;
  assign n24066 = ~n24063;
  assign n24106 = n24125 & n24126;
  assign n24109 = ~n24127;
  assign n24116 = n24128 & n392;
  assign n24117 = n24092 & n24129;
  assign n24118 = ~n24092;
  assign n23026 = ~n24138;
  assign n24134 = n20528 & n23006;
  assign n24130 = n24152 & n24153;
  assign n24139 = n24162 & n24163;
  assign n24086 = n24106 ^ n24107;
  assign n24108 = ~n24106;
  assign n24088 = ~n24116;
  assign n24094 = ~n24117;
  assign n24115 = n24118 & n24071;
  assign n24110 = n24130 ^ n24131;
  assign n23009 = ~n24134;
  assign n24132 = ~n24130;
  assign n24121 = n24139 ^ n21571;
  assign n24140 = ~n24139;
  assign n24064 = n392 ^ n24086;
  assign n24097 = n24108 & n24109;
  assign n24045 = n24110 ^ n24111;
  assign n24073 = ~n24115;
  assign n20425 = n24120 ^ n24121;
  assign n24119 = n24132 & n24133;
  assign n24135 = n24140 & n24141;
  assign n22623 = n24063 ^ n24064;
  assign n24065 = ~n24064;
  assign n24090 = n24045 & n407;
  assign n24087 = ~n24097;
  assign n24089 = ~n24045;
  assign n24051 = n20425 ^ n24098;
  assign n24100 = n20425 & n24114;
  assign n20471 = ~n20425;
  assign n24112 = ~n24119;
  assign n24122 = ~n24135;
  assign n23791 = ~n22623;
  assign n24022 = n24065 & n24066;
  assign n24067 = n24087 & n24088;
  assign n24077 = n24089 & n15473;
  assign n24047 = ~n24090;
  assign n24078 = n24051 & n24029;
  assign n24079 = ~n24051;
  assign n24095 = n20471 & n24099;
  assign n22991 = ~n24100;
  assign n24091 = n24112 & n24113;
  assign n24101 = n24122 & n24123;
  assign n24044 = n407 ^ n24067;
  assign n24068 = ~n24067;
  assign n24069 = ~n24077;
  assign n24053 = ~n24078;
  assign n24075 = n24079 & n24080;
  assign n24070 = n24091 ^ n24092;
  assign n22971 = ~n24095;
  assign n24093 = ~n24091;
  assign n24082 = n24101 ^ n21595;
  assign n24102 = ~n24101;
  assign n24023 = n24044 ^ n24045;
  assign n24056 = n24068 & n24069;
  assign n24025 = n24070 ^ n24071;
  assign n24031 = ~n24075;
  assign n24076 = n22991 & n22971;
  assign n20422 = n24082 ^ n24083;
  assign n24081 = n24093 & n24094;
  assign n24096 = n24102 & n24103;
  assign n23746 = n24022 ^ n24023;
  assign n23982 = n24023 & n24022;
  assign n24049 = n24025 & n406;
  assign n24046 = ~n24056;
  assign n24048 = ~n24025;
  assign n23989 = n24057 ^ n20422;
  assign n24058 = n20422 & n24074;
  assign n22989 = ~n24076;
  assign n20415 = ~n20422;
  assign n24072 = ~n24081;
  assign n24084 = ~n24096;
  assign n23762 = ~n23746;
  assign n24024 = n24046 & n24047;
  assign n24035 = n24048 & n15399;
  assign n24005 = ~n24049;
  assign n24038 = n23989 & n24010;
  assign n24036 = ~n23989;
  assign n22935 = ~n24058;
  assign n24054 = n20415 & n24059;
  assign n24050 = n24072 & n24073;
  assign n24060 = n24084 & n24085;
  assign n24003 = n24024 ^ n24025;
  assign n24026 = ~n24024;
  assign n24027 = ~n24035;
  assign n24033 = n24036 & n24037;
  assign n24012 = ~n24038;
  assign n24028 = n24050 ^ n24051;
  assign n22955 = ~n24054;
  assign n24052 = ~n24050;
  assign n24041 = n24060 ^ n21515;
  assign n24061 = ~n24060;
  assign n23983 = n406 ^ n24003;
  assign n24015 = n24026 & n24027;
  assign n23985 = n24028 ^ n24029;
  assign n23991 = ~n24033;
  assign n24034 = n22955 & n22935;
  assign n20374 = n24040 ^ n24041;
  assign n24039 = n24052 & n24053;
  assign n24055 = n24061 & n24062;
  assign n23695 = n23982 ^ n23983;
  assign n23942 = n23983 & n23982;
  assign n24006 = n23985 & n15354;
  assign n24004 = ~n24015;
  assign n24007 = ~n23985;
  assign n23948 = n24016 ^ n20374;
  assign n24017 = n20374 & n24032;
  assign n22953 = ~n24034;
  assign n20337 = ~n20374;
  assign n24030 = ~n24039;
  assign n24042 = ~n24055;
  assign n23708 = ~n23695;
  assign n23951 = ~n23942;
  assign n23984 = n24004 & n24005;
  assign n23987 = ~n24006;
  assign n23995 = n24007 & n405;
  assign n23996 = n23948 & n24008;
  assign n23997 = ~n23948;
  assign n22899 = ~n24017;
  assign n24013 = n20337 & n24018;
  assign n24009 = n24030 & n24031;
  assign n24019 = n24042 & n24043;
  assign n23963 = n23984 ^ n23985;
  assign n23986 = ~n23984;
  assign n23965 = ~n23995;
  assign n23950 = ~n23996;
  assign n23993 = n23997 & n23970;
  assign n23988 = n24009 ^ n24010;
  assign n22918 = ~n24013;
  assign n24011 = ~n24009;
  assign n23999 = n24019 ^ n21446;
  assign n24020 = ~n24019;
  assign n23943 = n405 ^ n23963;
  assign n23975 = n23986 & n23987;
  assign n23919 = n23988 ^ n23989;
  assign n23972 = ~n23993;
  assign n23994 = n22918 & n22899;
  assign n20335 = n23999 ^ n24000;
  assign n23998 = n24011 & n24012;
  assign n24014 = n24020 & n24021;
  assign n22408 = n23942 ^ n23943;
  assign n23899 = n23943 & n23951;
  assign n23966 = n23919 & n15327;
  assign n23964 = ~n23975;
  assign n23967 = ~n23919;
  assign n23925 = n23976 ^ n20335;
  assign n23977 = n20335 & n23992;
  assign n22916 = ~n23994;
  assign n20331 = ~n20335;
  assign n23990 = ~n23998;
  assign n24001 = ~n24014;
  assign n23636 = ~n22408;
  assign n23902 = ~n23899;
  assign n23944 = n23964 & n23965;
  assign n23946 = ~n23966;
  assign n23955 = n23967 & n404;
  assign n23957 = n23925 & n23968;
  assign n23956 = ~n23925;
  assign n23973 = n20331 & n22876;
  assign n22863 = ~n23977;
  assign n23969 = n23990 & n23991;
  assign n23979 = n24001 & n24002;
  assign n23918 = n404 ^ n23944;
  assign n23945 = ~n23944;
  assign n23921 = ~n23955;
  assign n23952 = n23956 & n23906;
  assign n23927 = ~n23957;
  assign n23947 = n23969 ^ n23970;
  assign n22878 = ~n23973;
  assign n23971 = ~n23969;
  assign n20247 = n23978 ^ n23979;
  assign n23980 = ~n23979;
  assign n23900 = n23918 ^ n23919;
  assign n23935 = n23945 & n23946;
  assign n23930 = n23947 ^ n23948;
  assign n23908 = ~n23952;
  assign n23958 = n23971 & n23972;
  assign n23960 = n20247 & n22839;
  assign n20290 = ~n20247;
  assign n23974 = n23980 & n23981;
  assign n23587 = n23899 ^ n23900;
  assign n23901 = ~n23900;
  assign n23923 = n23930 & n403;
  assign n23920 = ~n23935;
  assign n23922 = ~n23930;
  assign n23936 = n23953 ^ n20290;
  assign n23949 = ~n23958;
  assign n23954 = n20290 & n23959;
  assign n22841 = ~n23960;
  assign n23961 = ~n23974;
  assign n23603 = ~n23587;
  assign n23864 = n23901 & n23902;
  assign n23879 = n23920 & n23921;
  assign n23911 = n23922 & n15296;
  assign n23881 = ~n23923;
  assign n23931 = n23936 & n23937;
  assign n23924 = n23949 & n23950;
  assign n23932 = ~n23936;
  assign n22818 = ~n23954;
  assign n23938 = n23961 & n23962;
  assign n23903 = ~n23879;
  assign n23904 = ~n23911;
  assign n23905 = n23924 ^ n23925;
  assign n23871 = ~n23931;
  assign n23928 = n23932 & n23933;
  assign n23926 = ~n23924;
  assign n20269 = n23938 ^ n23939;
  assign n23940 = ~n23938;
  assign n23892 = n23903 & n23904;
  assign n23878 = n23904 & n23881;
  assign n23888 = n23905 ^ n23906;
  assign n23833 = n20269 ^ n23913;
  assign n23912 = n23926 & n23927;
  assign n23887 = ~n23928;
  assign n23915 = n20269 & n23929;
  assign n20262 = ~n20269;
  assign n23934 = n23940 & n23941;
  assign n23865 = n23878 ^ n23879;
  assign n23883 = n23888 & n402;
  assign n23880 = ~n23892;
  assign n23882 = ~n23888;
  assign n23893 = n23833 & n23909;
  assign n23884 = n23887 & n23871;
  assign n23894 = ~n23833;
  assign n23907 = ~n23912;
  assign n23910 = n20262 & n23914;
  assign n22768 = ~n23915;
  assign n23916 = ~n23934;
  assign n23526 = n23864 ^ n23865;
  assign n23824 = n23865 & n23864;
  assign n23845 = n23880 & n23881;
  assign n23873 = n23882 & n15251;
  assign n23847 = ~n23883;
  assign n23835 = ~n23893;
  assign n23889 = n23894 & n23850;
  assign n23885 = n23907 & n23908;
  assign n22793 = ~n23910;
  assign n23895 = n23916 & n23917;
  assign n23827 = ~n23824;
  assign n23866 = ~n23845;
  assign n23867 = ~n23873;
  assign n23829 = n23884 ^ n23885;
  assign n23852 = ~n23889;
  assign n23886 = ~n23885;
  assign n23890 = n22793 & n22768;
  assign n23875 = n23895 ^ n23896;
  assign n23897 = ~n23895;
  assign n23855 = n23866 & n23867;
  assign n23844 = n23867 & n23847;
  assign n23868 = n23829 & n15210;
  assign n23869 = ~n23829;
  assign n20230 = n23875 ^ n21083;
  assign n23874 = n23886 & n23887;
  assign n22791 = ~n23890;
  assign n23891 = n23897 & n23898;
  assign n23825 = n23844 ^ n23845;
  assign n23846 = ~n23855;
  assign n23811 = n23857 ^ n20230;
  assign n23831 = ~n23868;
  assign n23856 = n23869 & n401;
  assign n23858 = n20230 & n23872;
  assign n20175 = ~n20230;
  assign n23870 = ~n23874;
  assign n23876 = ~n23891;
  assign n22842 = n23824 ^ n23825;
  assign n23826 = ~n23825;
  assign n23828 = n23846 & n23847;
  assign n23838 = n23811 & n23848;
  assign n23839 = ~n23811;
  assign n23805 = ~n23856;
  assign n22721 = ~n23858;
  assign n23853 = n20175 & n23859;
  assign n23849 = n23870 & n23871;
  assign n23860 = n23876 & n23877;
  assign n22811 = n22842 ^ n22814;
  assign n23777 = n23802 ^ n22842;
  assign n23699 = n22842 & n21843;
  assign n23779 = n23826 & n23827;
  assign n23803 = n23828 ^ n23829;
  assign n23830 = ~n23828;
  assign n23813 = ~n23838;
  assign n23837 = n23839 & n23788;
  assign n23832 = n23849 ^ n23850;
  assign n22744 = ~n23853;
  assign n23851 = ~n23849;
  assign n23841 = n23860 ^ n23861;
  assign n23862 = ~n23860;
  assign n23051 = n487 ^ n23777;
  assign n19910 = n22811 ^ n23778;
  assign n23560 = n22811 & n23792;
  assign n23763 = n23777 & n487;
  assign n23780 = n401 ^ n23803;
  assign n23782 = ~n23779;
  assign n23816 = n23830 & n23831;
  assign n23784 = n23832 ^ n23833;
  assign n23790 = ~n23837;
  assign n22741 = n22744 & n22721;
  assign n20173 = n23841 ^ n20996;
  assign n23840 = n23851 & n23852;
  assign n23854 = n23862 & n23863;
  assign n23527 = n486 ^ n23763;
  assign n23766 = n23763 & n486;
  assign n23043 = ~n23051;
  assign n23764 = ~n23763;
  assign n23765 = n23779 ^ n23780;
  assign n23781 = ~n23780;
  assign n23807 = n23784 & n400;
  assign n23804 = ~n23816;
  assign n23806 = ~n23784;
  assign n23808 = n23817 ^ n20173;
  assign n23818 = n20173 & n23836;
  assign n20166 = ~n20173;
  assign n23834 = ~n23840;
  assign n23842 = ~n23854;
  assign n23750 = n23764 & n9791;
  assign n23752 = n23765 & n21819;
  assign n23513 = ~n23766;
  assign n23751 = ~n23765;
  assign n23728 = n23781 & n23782;
  assign n23783 = n23804 & n23805;
  assign n23794 = n23806 & n15157;
  assign n23755 = ~n23807;
  assign n23797 = n23808 & n23809;
  assign n23795 = ~n23808;
  assign n22663 = ~n23818;
  assign n23814 = n20166 & n23819;
  assign n23810 = n23834 & n23835;
  assign n23820 = n23842 & n23843;
  assign n23544 = ~n23750;
  assign n23737 = n23751 & n21753;
  assign n23727 = ~n23752;
  assign n23753 = n23783 ^ n23784;
  assign n23785 = ~n23783;
  assign n23786 = ~n23794;
  assign n23793 = n23795 & n23796;
  assign n23733 = ~n23797;
  assign n23787 = n23810 ^ n23811;
  assign n22687 = ~n23814;
  assign n23812 = ~n23810;
  assign n23799 = n23820 ^ n23821;
  assign n23822 = ~n23820;
  assign n23726 = n23727 & n23699;
  assign n23710 = ~n23737;
  assign n23729 = n400 ^ n23753;
  assign n23770 = n23785 & n23786;
  assign n23767 = n23787 ^ n23788;
  assign n23761 = ~n23793;
  assign n22684 = n22687 & n22663;
  assign n20148 = n23799 ^ n20913;
  assign n23798 = n23812 & n23813;
  assign n23815 = n23822 & n23823;
  assign n23709 = ~n23726;
  assign n23698 = n23727 & n23710;
  assign n23711 = n23728 ^ n23729;
  assign n23676 = n23729 & n23728;
  assign n23757 = n23767 & n415;
  assign n23754 = ~n23770;
  assign n23756 = ~n23767;
  assign n23739 = n23761 & n23733;
  assign n23758 = n23771 ^ n20148;
  assign n23772 = n20148 & n23791;
  assign n20090 = ~n20148;
  assign n23789 = ~n23798;
  assign n23800 = ~n23815;
  assign n19890 = n23698 ^ n23699;
  assign n23640 = n23709 & n23710;
  assign n23700 = n23711 & n21736;
  assign n23701 = ~n23711;
  assign n23679 = ~n23676;
  assign n23703 = n23754 & n23755;
  assign n23738 = n23756 & n15109;
  assign n23705 = ~n23757;
  assign n23741 = n23758 & n23759;
  assign n23742 = ~n23758;
  assign n22596 = ~n23772;
  assign n23768 = n20090 & n22623;
  assign n23740 = n23789 & n23790;
  assign n23773 = n23800 & n23801;
  assign n22722 = n19890 ^ n21753;
  assign n19892 = ~n19890;
  assign n23687 = ~n23640;
  assign n23675 = ~n23700;
  assign n23691 = n23701 & n21738;
  assign n23730 = ~n23703;
  assign n23731 = ~n23738;
  assign n23651 = n23739 ^ n23740;
  assign n23684 = ~n23741;
  assign n23735 = n23742 & n23743;
  assign n22625 = ~n23768;
  assign n23760 = ~n23740;
  assign n20032 = n23773 ^ n23774;
  assign n23775 = ~n23773;
  assign n23637 = n22698 ^ n22722;
  assign n23674 = n23675 & n23687;
  assign n23660 = ~n23691;
  assign n23717 = n23730 & n23731;
  assign n23718 = n23651 & n15067;
  assign n23702 = n23731 & n23705;
  assign n23719 = ~n23651;
  assign n23707 = ~n23735;
  assign n23633 = n23745 ^ n20032;
  assign n23744 = n23760 & n23761;
  assign n23747 = n20032 & n23762;
  assign n20111 = ~n20032;
  assign n23769 = n23775 & n23776;
  assign n23619 = n23637 & n23638;
  assign n23620 = ~n23637;
  assign n23659 = ~n23674;
  assign n23666 = n23660 & n23675;
  assign n23677 = n23702 ^ n23703;
  assign n23704 = ~n23717;
  assign n23682 = ~n23718;
  assign n23712 = n23719 & n414;
  assign n23713 = n23707 & n23684;
  assign n23720 = n23633 & n23734;
  assign n23721 = ~n23633;
  assign n23732 = ~n23744;
  assign n23736 = n20111 & n23746;
  assign n22525 = ~n23747;
  assign n23748 = ~n23769;
  assign n23562 = ~n23619;
  assign n23610 = n23620 & n23621;
  assign n23639 = n23659 & n23660;
  assign n23641 = ~n23666;
  assign n23605 = n23676 ^ n23677;
  assign n23678 = ~n23677;
  assign n23680 = n23704 & n23705;
  assign n23653 = ~n23712;
  assign n23689 = ~n23713;
  assign n23635 = ~n23720;
  assign n23714 = n23721 & n23656;
  assign n23688 = n23732 & n23733;
  assign n22562 = ~n23736;
  assign n23722 = n23748 & n23749;
  assign n23590 = ~n23610;
  assign n23604 = n23639 ^ n21577;
  assign n19797 = n23640 ^ n23641;
  assign n23622 = ~n23639;
  assign n23648 = n23605 & n21591;
  assign n23649 = ~n23605;
  assign n23624 = n23678 & n23679;
  assign n23650 = n414 ^ n23680;
  assign n23629 = n23688 ^ n23689;
  assign n23681 = ~n23680;
  assign n23658 = ~n23714;
  assign n23706 = ~n23688;
  assign n23715 = n22562 & n22525;
  assign n20011 = n23722 ^ n23723;
  assign n23724 = ~n23722;
  assign n23578 = n23590 & n23560;
  assign n23559 = n23590 & n23562;
  assign n19768 = n23604 ^ n23605;
  assign n22664 = n19797 ^ n21738;
  assign n19794 = ~n19797;
  assign n23592 = ~n23648;
  assign n23642 = n23649 & n21577;
  assign n23625 = n23650 ^ n23651;
  assign n23627 = ~n23624;
  assign n23662 = n23629 & n413;
  assign n23667 = n23681 & n23682;
  assign n23661 = ~n23629;
  assign n23685 = n23693 ^ n20011;
  assign n23692 = n23706 & n23707;
  assign n23694 = n20011 & n23708;
  assign n22560 = ~n23715;
  assign n20022 = ~n20011;
  assign n23716 = n23724 & n23725;
  assign n23528 = n23559 ^ n23560;
  assign n22600 = n19768 ^ n21591;
  assign n23561 = ~n23578;
  assign n23563 = n22664 ^ n22589;
  assign n19751 = ~n19768;
  assign n23606 = n23624 ^ n23625;
  assign n23623 = ~n23642;
  assign n23626 = ~n23625;
  assign n23654 = n23661 & n15056;
  assign n23596 = ~n23662;
  assign n23652 = ~n23667;
  assign n23668 = n23685 & n23686;
  assign n23669 = ~n23685;
  assign n23683 = ~n23692;
  assign n22451 = ~n23694;
  assign n23690 = n20022 & n23695;
  assign n23696 = ~n23716;
  assign n21744 = n23527 ^ n23528;
  assign n23529 = n23528 & n23544;
  assign n23519 = n22600 ^ n22488;
  assign n23488 = n23561 & n23562;
  assign n23548 = n23563 & n23564;
  assign n23549 = ~n23563;
  assign n23593 = n23606 & n21486;
  assign n23531 = ~n23606;
  assign n23611 = n23622 & n23623;
  assign n23568 = n23626 & n23627;
  assign n23628 = n23652 & n23653;
  assign n23631 = ~n23654;
  assign n23575 = ~n23668;
  assign n23663 = n23669 & n23670;
  assign n23655 = n23683 & n23684;
  assign n22485 = ~n23690;
  assign n23671 = n23696 & n23697;
  assign n23514 = n23519 & n23520;
  assign n22987 = ~n21744;
  assign n23512 = ~n23529;
  assign n23515 = ~n23519;
  assign n23522 = ~n23488;
  assign n23492 = ~n23548;
  assign n23545 = n23549 & n23550;
  assign n23579 = n23531 & n21533;
  assign n23567 = ~n23593;
  assign n23591 = ~n23611;
  assign n23594 = n23628 ^ n23629;
  assign n23630 = ~n23628;
  assign n23632 = n23655 ^ n23656;
  assign n23602 = ~n23663;
  assign n23657 = ~n23655;
  assign n23664 = n22485 & n22451;
  assign n23645 = n23671 ^ n20692;
  assign n23672 = ~n23671;
  assign n23396 = n23512 & n23513;
  assign n23441 = ~n23514;
  assign n23496 = n23515 & n23516;
  assign n23521 = ~n23545;
  assign n23533 = ~n23579;
  assign n23565 = n23591 & n23592;
  assign n23569 = n413 ^ n23594;
  assign n23612 = n23630 & n23631;
  assign n23607 = n23632 ^ n23633;
  assign n23599 = n23602 & n23575;
  assign n20009 = n23644 ^ n23645;
  assign n23643 = n23657 & n23658;
  assign n22483 = ~n23664;
  assign n23665 = n23672 & n23673;
  assign n23439 = ~n23396;
  assign n23466 = ~n23496;
  assign n23517 = n23521 & n23522;
  assign n23518 = n23521 & n23492;
  assign n23530 = n23565 ^ n21486;
  assign n23473 = n23568 ^ n23569;
  assign n23500 = n23569 & n23568;
  assign n23566 = ~n23565;
  assign n23598 = n23607 & n412;
  assign n23595 = ~n23612;
  assign n23597 = ~n23607;
  assign n23509 = n23613 ^ n20009;
  assign n23614 = n20009 & n23636;
  assign n20000 = ~n20009;
  assign n23634 = ~n23643;
  assign n23646 = ~n23665;
  assign n23472 = n23466 & n23441;
  assign n23491 = ~n23517;
  assign n23489 = ~n23518;
  assign n19744 = n23530 ^ n23531;
  assign n23535 = n23473 & n21453;
  assign n23534 = ~n23473;
  assign n23551 = n23566 & n23567;
  assign n23503 = ~n23500;
  assign n23537 = n23595 & n23596;
  assign n23580 = n23597 & n14988;
  assign n23539 = ~n23598;
  assign n23583 = n23509 & n23541;
  assign n23581 = ~n23509;
  assign n23608 = n20000 & n22408;
  assign n22375 = ~n23614;
  assign n23600 = n23634 & n23635;
  assign n23615 = n23646 & n23647;
  assign n23447 = ~n23472;
  assign n23468 = n23488 ^ n23489;
  assign n23446 = n23491 & n23492;
  assign n22535 = n19744 ^ n21533;
  assign n19738 = ~n19744;
  assign n23523 = n23534 & n21471;
  assign n23498 = ~n23535;
  assign n23532 = ~n23551;
  assign n23570 = ~n23537;
  assign n23571 = ~n23580;
  assign n23576 = n23581 & n23582;
  assign n23542 = ~n23583;
  assign n23505 = n23599 ^ n23600;
  assign n22410 = ~n23608;
  assign n23601 = ~n23600;
  assign n19981 = n23615 ^ n23616;
  assign n23617 = ~n23615;
  assign n23374 = n23446 ^ n23447;
  assign n23465 = n23468 & n485;
  assign n23388 = n22535 ^ n22455;
  assign n23464 = ~n23468;
  assign n23467 = ~n23446;
  assign n23476 = ~n23523;
  assign n23497 = n23532 & n23533;
  assign n23552 = n23570 & n23571;
  assign n23536 = n23571 & n23539;
  assign n23572 = n23505 & n14942;
  assign n23511 = ~n23576;
  assign n23573 = ~n23505;
  assign n23460 = n19981 ^ n23585;
  assign n23584 = n23601 & n23602;
  assign n23586 = n19981 & n23603;
  assign n19926 = ~n19981;
  assign n23609 = n23617 & n23618;
  assign n23423 = n23374 & n484;
  assign n23422 = ~n23374;
  assign n23450 = n23388 & n23415;
  assign n23451 = n23464 & n9753;
  assign n23412 = ~n23465;
  assign n23463 = n23466 & n23467;
  assign n23448 = ~n23388;
  assign n23474 = n23497 ^ n21471;
  assign n23499 = ~n23497;
  assign n23501 = n23536 ^ n23537;
  assign n23538 = ~n23552;
  assign n23507 = ~n23572;
  assign n23553 = n23573 & n411;
  assign n23554 = n23460 & n23485;
  assign n23555 = ~n23460;
  assign n23574 = ~n23584;
  assign n22299 = ~n23586;
  assign n23577 = n19926 & n23587;
  assign n23588 = ~n23609;
  assign n23413 = n23422 & n9721;
  assign n23363 = ~n23423;
  assign n23442 = n23448 & n23449;
  assign n23390 = ~n23450;
  assign n23438 = ~n23451;
  assign n23440 = ~n23463;
  assign n19703 = n23473 ^ n23474;
  assign n23493 = n23498 & n23499;
  assign n23490 = n23500 ^ n23501;
  assign n23502 = ~n23501;
  assign n23504 = n23538 & n23539;
  assign n23481 = ~n23553;
  assign n23462 = ~n23554;
  assign n23546 = n23555 & n23556;
  assign n23540 = n23574 & n23575;
  assign n22311 = ~n23577;
  assign n23557 = n23588 & n23589;
  assign n23385 = ~n23413;
  assign n23424 = n23438 & n23439;
  assign n23425 = n23438 & n23412;
  assign n23414 = n23440 & n23441;
  assign n23416 = ~n23442;
  assign n22440 = n19703 ^ n21471;
  assign n19699 = ~n19703;
  assign n23478 = n23490 & n21318;
  assign n23475 = ~n23493;
  assign n23477 = ~n23490;
  assign n23454 = n23502 & n23503;
  assign n23479 = n23504 ^ n23505;
  assign n23506 = ~n23504;
  assign n23508 = n23540 ^ n23541;
  assign n23487 = ~n23546;
  assign n23543 = ~n23540;
  assign n23547 = n22311 & n22299;
  assign n19931 = n23557 ^ n23558;
  assign n23387 = n23414 ^ n23415;
  assign n23343 = n22440 ^ n22416;
  assign n23411 = ~n23424;
  assign n23397 = ~n23425;
  assign n23417 = ~n23414;
  assign n23419 = n23475 & n23476;
  assign n23469 = n23477 & n21390;
  assign n23427 = ~n23478;
  assign n23455 = n411 ^ n23479;
  assign n23494 = n23506 & n23507;
  assign n23431 = n23508 ^ n23509;
  assign n23495 = n23525 ^ n19931;
  assign n22260 = n23526 ^ n19931;
  assign n23524 = n23542 & n23543;
  assign n22339 = ~n23547;
  assign n23315 = n23387 ^ n23388;
  assign n22979 = n23396 ^ n23397;
  assign n23394 = n23343 & n23409;
  assign n23398 = n23411 & n23412;
  assign n23410 = n23416 & n23417;
  assign n23395 = ~n23343;
  assign n23376 = n23454 ^ n23455;
  assign n23402 = n23455 & n23454;
  assign n23452 = ~n23419;
  assign n23453 = ~n23469;
  assign n23482 = n23431 & n14910;
  assign n23480 = ~n23494;
  assign n23483 = ~n23431;
  assign n23437 = n408 ^ n23495;
  assign n22273 = ~n22260;
  assign n23510 = ~n23524;
  assign n23365 = n23315 & n9697;
  assign n23366 = ~n23315;
  assign n22969 = ~n22979;
  assign n23345 = ~n23394;
  assign n23391 = n23395 & n23368;
  assign n23373 = ~n23398;
  assign n23389 = ~n23410;
  assign n23428 = n23376 & n21210;
  assign n23429 = ~n23376;
  assign n23443 = n23452 & n23453;
  assign n23444 = n23453 & n23427;
  assign n23405 = ~n23402;
  assign n23456 = n23480 & n23481;
  assign n23458 = ~n23482;
  assign n23470 = n23483 & n410;
  assign n23484 = n23510 & n23511;
  assign n23337 = ~n23365;
  assign n23361 = n23366 & n483;
  assign n23351 = n23373 ^ n23374;
  assign n23372 = n23385 & n23373;
  assign n23367 = n23389 & n23390;
  assign n23370 = ~n23391;
  assign n23378 = ~n23428;
  assign n23418 = n23429 & n21341;
  assign n23426 = ~n23443;
  assign n23420 = ~n23444;
  assign n23430 = n410 ^ n23456;
  assign n23457 = ~n23456;
  assign n23433 = ~n23470;
  assign n23459 = n23484 ^ n23485;
  assign n23486 = ~n23484;
  assign n22932 = n484 ^ n23351;
  assign n23317 = ~n23361;
  assign n23342 = n23367 ^ n23368;
  assign n23362 = ~n23372;
  assign n23369 = ~n23367;
  assign n23401 = ~n23418;
  assign n19663 = n23419 ^ n23420;
  assign n23399 = n23426 & n23427;
  assign n23403 = n23430 ^ n23431;
  assign n23445 = n23457 & n23458;
  assign n23382 = n23459 ^ n23460;
  assign n23471 = n23486 & n23487;
  assign n23329 = n23342 ^ n23343;
  assign n22942 = ~n22932;
  assign n23339 = n23362 & n23363;
  assign n23364 = n23369 & n23370;
  assign n22378 = n19663 ^ n21318;
  assign n23375 = n23399 ^ n21341;
  assign n23386 = n23402 ^ n23403;
  assign n19651 = ~n19663;
  assign n23400 = ~n23399;
  assign n23404 = ~n23403;
  assign n23434 = n23382 & n14879;
  assign n23432 = ~n23445;
  assign n23435 = ~n23382;
  assign n23461 = ~n23471;
  assign n23323 = n23329 & n482;
  assign n23322 = ~n23329;
  assign n23314 = n483 ^ n23339;
  assign n23338 = ~n23339;
  assign n23344 = ~n23364;
  assign n23352 = n22378 ^ n22354;
  assign n19645 = n23375 ^ n23376;
  assign n23380 = n23386 & n21171;
  assign n23379 = ~n23386;
  assign n23392 = n23400 & n23401;
  assign n23356 = n23404 & n23405;
  assign n23406 = n23432 & n23433;
  assign n23408 = ~n23434;
  assign n23421 = n23435 & n409;
  assign n23436 = n23461 & n23462;
  assign n23296 = n23314 ^ n23315;
  assign n23318 = n23322 & n9663;
  assign n23281 = ~n23323;
  assign n23330 = n23337 & n23338;
  assign n23300 = n23344 & n23345;
  assign n22290 = n19645 ^ n21210;
  assign n23346 = n23352 & n23353;
  assign n23347 = ~n23352;
  assign n19601 = ~n19645;
  assign n23371 = n23379 & n21226;
  assign n23355 = ~n23380;
  assign n23377 = ~n23392;
  assign n23381 = n409 ^ n23406;
  assign n23407 = ~n23406;
  assign n23384 = ~n23421;
  assign n23360 = n23436 ^ n23437;
  assign n22896 = n23296 ^ n22932;
  assign n23297 = ~n23296;
  assign n23299 = ~n23318;
  assign n23316 = ~n23330;
  assign n23288 = n22290 ^ n22209;
  assign n23324 = ~n23300;
  assign n23303 = ~n23346;
  assign n23340 = n23347 & n23348;
  assign n23332 = ~n23371;
  assign n23326 = n23377 & n23378;
  assign n23357 = n23381 ^ n23382;
  assign n23393 = n23407 & n23408;
  assign n22909 = ~n22896;
  assign n23265 = n23297 & n22942;
  assign n23285 = n23299 & n23281;
  assign n23286 = n23316 & n23317;
  assign n23309 = n23288 & n23319;
  assign n23308 = ~n23288;
  assign n23325 = ~n23340;
  assign n23350 = n23355 & n23332;
  assign n23341 = n23356 ^ n23357;
  assign n23354 = ~n23326;
  assign n23358 = ~n23357;
  assign n23383 = ~n23393;
  assign n23266 = n23285 ^ n23286;
  assign n23298 = ~n23286;
  assign n23304 = n23308 & n23268;
  assign n23290 = ~n23309;
  assign n23320 = n23324 & n23325;
  assign n23321 = n23325 & n23303;
  assign n23333 = n23341 & n21089;
  assign n23327 = ~n23350;
  assign n23334 = ~n23341;
  assign n23349 = n23354 & n23355;
  assign n23335 = n23358 & n23356;
  assign n23359 = n23383 & n23384;
  assign n22837 = n23265 ^ n23266;
  assign n23224 = n23266 & n23265;
  assign n23293 = n23298 & n23299;
  assign n23270 = ~n23304;
  assign n23302 = ~n23320;
  assign n23301 = ~n23321;
  assign n19550 = n23326 ^ n23327;
  assign n23295 = ~n23333;
  assign n23328 = n23334 & n21176;
  assign n23331 = ~n23349;
  assign n23336 = n23359 ^ n23360;
  assign n22850 = ~n22837;
  assign n23280 = ~n23293;
  assign n23261 = n23300 ^ n23301;
  assign n23287 = n23302 & n23303;
  assign n22223 = n21171 ^ n19550;
  assign n19581 = ~n19550;
  assign n23311 = ~n23328;
  assign n23291 = n23331 & n23332;
  assign n23277 = n23335 ^ n23336;
  assign n23260 = n23280 & n23281;
  assign n23267 = n23287 ^ n23288;
  assign n23284 = n23261 & n481;
  assign n23253 = n22223 ^ n22098;
  assign n23283 = ~n23261;
  assign n23289 = ~n23287;
  assign n23306 = n23311 & n23295;
  assign n23313 = n23277 & n21004;
  assign n23310 = ~n23291;
  assign n23312 = ~n23277;
  assign n23244 = n23260 ^ n23261;
  assign n23256 = n23267 ^ n23268;
  assign n23262 = ~n23260;
  assign n23272 = n23253 & n23275;
  assign n23274 = n23283 & n9619;
  assign n23246 = ~n23284;
  assign n23271 = ~n23253;
  assign n23282 = n23289 & n23290;
  assign n23292 = ~n23306;
  assign n23305 = n23310 & n23311;
  assign n23307 = n23312 & n21074;
  assign n23279 = ~n23313;
  assign n23225 = n481 ^ n23244;
  assign n23251 = n23256 & n480;
  assign n23250 = ~n23256;
  assign n23264 = n23271 & n23230;
  assign n23255 = ~n23272;
  assign n23263 = ~n23274;
  assign n23269 = ~n23282;
  assign n19529 = n23291 ^ n23292;
  assign n23294 = ~n23305;
  assign n23259 = ~n23307;
  assign n21414 = n23224 ^ n23225;
  assign n23194 = n23225 & n23224;
  assign n23247 = n23250 & n9577;
  assign n23208 = ~n23251;
  assign n23257 = n23262 & n23263;
  assign n23232 = ~n23264;
  assign n23252 = n23269 & n23270;
  assign n22149 = n19529 ^ n21089;
  assign n19527 = ~n19529;
  assign n23276 = n23294 & n23295;
  assign n22789 = ~n21414;
  assign n23227 = ~n23247;
  assign n23229 = n23252 ^ n23253;
  assign n23197 = n22149 ^ n22127;
  assign n23245 = ~n23257;
  assign n23254 = ~n23252;
  assign n22084 = n23276 ^ n23277;
  assign n23278 = ~n23276;
  assign n23212 = n23227 & n23208;
  assign n23220 = n23229 ^ n23230;
  assign n23233 = n23197 & n23237;
  assign n23213 = n23245 & n23246;
  assign n23234 = ~n23197;
  assign n23248 = n23254 & n23255;
  assign n23166 = n22084 ^ n22065;
  assign n19452 = n22084 ^ n21074;
  assign n23273 = n23278 & n23279;
  assign n23195 = n23212 ^ n23213;
  assign n23215 = n23220 & n495;
  assign n23214 = ~n23220;
  assign n23199 = ~n23233;
  assign n23228 = n23234 & n23217;
  assign n23226 = ~n23213;
  assign n23231 = ~n23248;
  assign n23238 = n23166 & n23249;
  assign n23239 = ~n23166;
  assign n19511 = ~n19452;
  assign n23258 = ~n23273;
  assign n21375 = n23194 ^ n23195;
  assign n23161 = n23195 & n23194;
  assign n23209 = n23214 & n9544;
  assign n23175 = ~n23215;
  assign n23221 = n23226 & n23227;
  assign n23219 = ~n23228;
  assign n23216 = n23231 & n23232;
  assign n23168 = ~n23238;
  assign n23235 = n23239 & n23183;
  assign n23240 = n23258 & n23259;
  assign n22776 = ~n21375;
  assign n23164 = ~n23161;
  assign n23193 = ~n23209;
  assign n23196 = n23216 ^ n23217;
  assign n23207 = ~n23221;
  assign n23218 = ~n23216;
  assign n23185 = ~n23235;
  assign n22031 = n23240 ^ n23241;
  assign n23242 = ~n23240;
  assign n23178 = n23193 & n23175;
  assign n23186 = n23196 ^ n23197;
  assign n23179 = n23207 & n23208;
  assign n23210 = n23218 & n23219;
  assign n23130 = n22031 ^ n22010;
  assign n19494 = n22031 ^ n20878;
  assign n23236 = n23242 & n23243;
  assign n23162 = n23178 ^ n23179;
  assign n23181 = n23186 & n494;
  assign n23180 = ~n23186;
  assign n23192 = ~n23179;
  assign n23198 = ~n23210;
  assign n23202 = n23130 & n23211;
  assign n23203 = ~n23130;
  assign n19487 = ~n19494;
  assign n23222 = ~n23236;
  assign n22719 = n23161 ^ n23162;
  assign n23163 = ~n23162;
  assign n23176 = n23180 & n9510;
  assign n23144 = ~n23181;
  assign n23187 = n23192 & n23193;
  assign n23182 = n23198 & n23199;
  assign n23132 = ~n23202;
  assign n23200 = n23203 & n23151;
  assign n23204 = n23222 & n23223;
  assign n22730 = ~n22719;
  assign n23123 = n23163 & n23164;
  assign n23159 = ~n23176;
  assign n23165 = n23182 ^ n23183;
  assign n23174 = ~n23187;
  assign n23184 = ~n23182;
  assign n23153 = ~n23200;
  assign n23188 = n23204 ^ n20928;
  assign n23205 = ~n23204;
  assign n23160 = n23159 & n23144;
  assign n23154 = n23165 ^ n23166;
  assign n23141 = n23174 & n23175;
  assign n23177 = n23184 & n23185;
  assign n19434 = n23188 ^ n23189;
  assign n23201 = n23205 & n23206;
  assign n23149 = n23154 & n493;
  assign n23142 = ~n23160;
  assign n23148 = ~n23154;
  assign n23158 = ~n23141;
  assign n21961 = n19434 ^ n20938;
  assign n23167 = ~n23177;
  assign n19399 = ~n19434;
  assign n23190 = ~n23201;
  assign n23124 = n23141 ^ n23142;
  assign n23145 = n23148 & n9459;
  assign n23108 = ~n23149;
  assign n23097 = n21961 ^ n21953;
  assign n23155 = n23158 & n23159;
  assign n23150 = n23167 & n23168;
  assign n23170 = n23190 & n23191;
  assign n22660 = n23123 ^ n23124;
  assign n23086 = n23124 & n23123;
  assign n23126 = ~n23145;
  assign n23136 = n23097 & n23146;
  assign n23129 = n23150 ^ n23151;
  assign n23135 = ~n23097;
  assign n23143 = ~n23155;
  assign n23152 = ~n23150;
  assign n19339 = n23170 ^ n23171;
  assign n23172 = ~n23170;
  assign n22672 = ~n22660;
  assign n23089 = ~n23086;
  assign n23127 = n23126 & n23108;
  assign n23091 = n23129 ^ n23130;
  assign n23133 = n23135 & n23114;
  assign n23099 = ~n23136;
  assign n23105 = n23143 & n23144;
  assign n23147 = n23152 & n23153;
  assign n21927 = n19339 ^ n20825;
  assign n19418 = ~n19339;
  assign n23169 = n23172 & n23173;
  assign n23112 = n23091 & n492;
  assign n23106 = ~n23127;
  assign n23111 = ~n23091;
  assign n23116 = ~n23133;
  assign n23125 = ~n23105;
  assign n23053 = n21927 ^ n21910;
  assign n23131 = ~n23147;
  assign n23156 = ~n23169;
  assign n23087 = n23105 ^ n23106;
  assign n23109 = n23111 & n9421;
  assign n23068 = ~n23112;
  assign n23118 = n23125 & n23126;
  assign n23119 = n23053 & n23128;
  assign n23113 = n23131 & n23132;
  assign n23120 = ~n23053;
  assign n23137 = n23156 & n23157;
  assign n22558 = n23086 ^ n23087;
  assign n23088 = ~n23087;
  assign n23093 = ~n23109;
  assign n23096 = n23113 ^ n23114;
  assign n23107 = ~n23118;
  assign n23055 = ~n23119;
  assign n23117 = n23120 & n23076;
  assign n23115 = ~n23113;
  assign n19354 = n23137 ^ n23138;
  assign n23139 = ~n23137;
  assign n22576 = ~n22558;
  assign n23046 = n23088 & n23089;
  assign n23028 = n23096 ^ n23097;
  assign n23090 = n23107 & n23108;
  assign n23110 = n23115 & n23116;
  assign n23078 = ~n23117;
  assign n21886 = n19354 ^ n20749;
  assign n19346 = ~n19354;
  assign n23134 = n23139 & n23140;
  assign n23074 = n23028 & n491;
  assign n23066 = n23090 ^ n23091;
  assign n23073 = ~n23028;
  assign n23092 = ~n23090;
  assign n23094 = n21886 ^ n21867;
  assign n23098 = ~n23110;
  assign n23121 = ~n23134;
  assign n23047 = n492 ^ n23066;
  assign n23069 = n23073 & n9407;
  assign n23030 = ~n23074;
  assign n23080 = n23092 & n23093;
  assign n23083 = n23094 & n23095;
  assign n23075 = n23098 & n23099;
  assign n23081 = ~n23094;
  assign n23101 = n23121 & n23122;
  assign n22523 = n23046 ^ n23047;
  assign n23010 = n23047 & n23046;
  assign n23050 = ~n23069;
  assign n23052 = n23075 ^ n23076;
  assign n23067 = ~n23080;
  assign n23079 = n23081 & n23082;
  assign n23021 = ~n23083;
  assign n23077 = ~n23075;
  assign n21816 = n23101 ^ n23102;
  assign n23103 = ~n23101;
  assign n22541 = ~n22523;
  assign n22993 = n23052 ^ n23053;
  assign n23048 = n23067 & n23068;
  assign n23070 = n23077 & n23078;
  assign n23038 = ~n23079;
  assign n23071 = n21816 ^ n21803;
  assign n19331 = n21816 ^ n20562;
  assign n23100 = n23103 & n23104;
  assign n23034 = n22993 & n490;
  assign n23027 = n491 ^ n23048;
  assign n23033 = ~n22993;
  assign n23049 = ~n23048;
  assign n23056 = n23038 & n23021;
  assign n23054 = ~n23070;
  assign n23061 = n23071 & n23072;
  assign n23059 = ~n23071;
  assign n19325 = ~n19331;
  assign n23084 = ~n23100;
  assign n23011 = n23027 ^ n23028;
  assign n23031 = n23033 & n9340;
  assign n22995 = ~n23034;
  assign n23041 = n23049 & n23050;
  assign n23035 = n23054 & n23055;
  assign n23036 = ~n23056;
  assign n23057 = n23059 & n23060;
  assign n22983 = ~n23061;
  assign n23062 = n23084 & n23085;
  assign n22449 = n23010 ^ n23011;
  assign n22972 = n23011 & n23010;
  assign n23014 = ~n23031;
  assign n23023 = n23035 ^ n23036;
  assign n23029 = ~n23041;
  assign n23037 = ~n23035;
  assign n23000 = ~n23057;
  assign n19271 = n23062 ^ n23063;
  assign n23064 = ~n23062;
  assign n22470 = ~n22449;
  assign n23019 = n23023 & n489;
  assign n23012 = n23029 & n23030;
  assign n23018 = ~n23023;
  assign n23032 = n23037 & n23038;
  assign n23039 = n23000 & n22983;
  assign n21792 = n19271 ^ n20579;
  assign n23042 = n19271 & n23051;
  assign n19235 = ~n19271;
  assign n23058 = n23064 & n23065;
  assign n22992 = n490 ^ n23012;
  assign n23015 = n23018 & n9304;
  assign n22959 = ~n23019;
  assign n23013 = ~n23012;
  assign n23016 = n21792 ^ n21773;
  assign n23020 = ~n23032;
  assign n22998 = ~n23039;
  assign n21805 = ~n23042;
  assign n23040 = n19235 & n23043;
  assign n23044 = ~n23058;
  assign n22973 = n22992 ^ n22993;
  assign n23002 = n23013 & n23014;
  assign n22977 = ~n23015;
  assign n23003 = n23016 & n23017;
  assign n22997 = n23020 & n23021;
  assign n23004 = ~n23016;
  assign n21831 = ~n23040;
  assign n23024 = n23044 & n23045;
  assign n22338 = n22972 ^ n22973;
  assign n22956 = n22973 & n22972;
  assign n22974 = n22977 & n22959;
  assign n22937 = n22997 ^ n22998;
  assign n22994 = ~n23002;
  assign n22946 = ~n23003;
  assign n23001 = n23004 & n23005;
  assign n22999 = ~n22997;
  assign n21828 = n21805 & n21831;
  assign n23007 = n23024 ^ n20517;
  assign n23025 = ~n23024;
  assign n22352 = ~n22338;
  assign n22981 = n22937 & n488;
  assign n22975 = n22994 & n22995;
  assign n22980 = ~n22937;
  assign n22996 = n22999 & n23000;
  assign n22965 = ~n23001;
  assign n19260 = n23006 ^ n23007;
  assign n23022 = n23025 & n23026;
  assign n22957 = n22974 ^ n22975;
  assign n22978 = n22980 & n9262;
  assign n22921 = ~n22981;
  assign n22976 = ~n22975;
  assign n22962 = n22965 & n22946;
  assign n21708 = n20528 ^ n19260;
  assign n22982 = ~n22996;
  assign n22986 = n19260 & n21744;
  assign n19248 = ~n19260;
  assign n23008 = ~n23022;
  assign n22297 = n22956 ^ n22957;
  assign n22900 = n22957 & n22956;
  assign n22924 = n21708 ^ n21685;
  assign n22967 = n22976 & n22977;
  assign n22939 = ~n22978;
  assign n22963 = n22982 & n22983;
  assign n21747 = ~n22986;
  assign n22984 = n19248 & n22987;
  assign n22988 = n23008 & n23009;
  assign n22309 = ~n22297;
  assign n22903 = ~n22900;
  assign n22951 = n22924 & n22960;
  assign n22905 = n22962 ^ n22963;
  assign n22950 = ~n22924;
  assign n22958 = ~n22967;
  assign n22964 = ~n22963;
  assign n21776 = ~n22984;
  assign n19211 = n22988 ^ n22989;
  assign n22990 = ~n22988;
  assign n22943 = n22905 & n9219;
  assign n22947 = n22950 & n22911;
  assign n22926 = ~n22951;
  assign n22936 = n22958 & n22959;
  assign n22944 = ~n22905;
  assign n22961 = n22964 & n22965;
  assign n21676 = n19211 ^ n20471;
  assign n22968 = n19211 & n22979;
  assign n19143 = ~n19211;
  assign n22985 = n22990 & n22991;
  assign n22919 = n22936 ^ n22937;
  assign n22907 = ~n22943;
  assign n22940 = n22944 & n503;
  assign n22913 = ~n22947;
  assign n22938 = ~n22936;
  assign n22887 = n21676 ^ n21641;
  assign n22945 = ~n22961;
  assign n21678 = ~n22968;
  assign n22966 = n19143 & n22969;
  assign n22970 = ~n22985;
  assign n22901 = n488 ^ n22919;
  assign n22929 = n22938 & n22939;
  assign n22881 = ~n22940;
  assign n22931 = n22887 & n22941;
  assign n22923 = n22945 & n22946;
  assign n22930 = ~n22887;
  assign n21712 = ~n22966;
  assign n22952 = n22970 & n22971;
  assign n22186 = n22900 ^ n22901;
  assign n22902 = ~n22901;
  assign n22910 = n22923 ^ n22924;
  assign n22920 = ~n22929;
  assign n22927 = n22930 & n22871;
  assign n22889 = ~n22931;
  assign n22925 = ~n22923;
  assign n22948 = n21712 & n21678;
  assign n19170 = n22952 ^ n22953;
  assign n22954 = ~n22952;
  assign n22864 = n22902 & n22903;
  assign n22892 = n22910 ^ n22911;
  assign n22904 = n22920 & n22921;
  assign n22922 = n22925 & n22926;
  assign n22873 = ~n22927;
  assign n21613 = n19170 ^ n20422;
  assign n21643 = n22932 ^ n19170;
  assign n22933 = n19170 & n22942;
  assign n21710 = ~n22948;
  assign n19122 = ~n19170;
  assign n22949 = n22954 & n22955;
  assign n22885 = n22892 & n502;
  assign n22879 = n22904 ^ n22905;
  assign n22884 = ~n22892;
  assign n22906 = ~n22904;
  assign n22854 = n21613 ^ n21583;
  assign n22912 = ~n22922;
  assign n21615 = ~n22933;
  assign n22928 = n19122 & n22932;
  assign n22934 = ~n22949;
  assign n22865 = n503 ^ n22879;
  assign n22882 = n22884 & n9190;
  assign n22846 = ~n22885;
  assign n22893 = n22906 & n22907;
  assign n22895 = n22854 & n22908;
  assign n22886 = n22912 & n22913;
  assign n22894 = ~n22854;
  assign n21645 = ~n22928;
  assign n22915 = n22934 & n22935;
  assign n19855 = n22864 ^ n22865;
  assign n22819 = n22865 & n22864;
  assign n22867 = ~n22882;
  assign n22870 = n22886 ^ n22887;
  assign n22880 = ~n22893;
  assign n22890 = n22894 & n22827;
  assign n22856 = ~n22895;
  assign n22888 = ~n22886;
  assign n19063 = n22915 ^ n22916;
  assign n22917 = ~n22915;
  assign n21864 = n19855 ^ n22842;
  assign n22746 = n19855 & n19910;
  assign n19871 = ~n19855;
  assign n22822 = ~n22819;
  assign n22868 = n22867 & n22846;
  assign n22858 = n22870 ^ n22871;
  assign n22843 = n22880 & n22881;
  assign n22883 = n22888 & n22889;
  assign n22829 = ~n22890;
  assign n21547 = n19063 ^ n20374;
  assign n22897 = n19063 & n22909;
  assign n19146 = ~n19063;
  assign n22914 = n22917 & n22918;
  assign n22812 = n22833 ^ n19871;
  assign n22852 = n22858 & n501;
  assign n22844 = ~n22868;
  assign n22851 = ~n22858;
  assign n22866 = ~n22843;
  assign n22807 = n21547 ^ n21515;
  assign n22872 = ~n22883;
  assign n22891 = n19146 & n22896;
  assign n21553 = ~n22897;
  assign n22898 = ~n22914;
  assign n18803 = n22811 ^ n22812;
  assign n21298 = n71 ^ n22812;
  assign n22530 = n22812 & n71;
  assign n22813 = ~n22812;
  assign n22820 = n22843 ^ n22844;
  assign n22847 = n22851 & n9138;
  assign n22799 = ~n22852;
  assign n22859 = n22866 & n22867;
  assign n22861 = n22807 & n22869;
  assign n22853 = n22872 & n22873;
  assign n22860 = ~n22807;
  assign n21588 = ~n22891;
  assign n22875 = n22898 & n22899;
  assign n21863 = ~n18803;
  assign n21310 = ~n21298;
  assign n22630 = n22813 & n22814;
  assign n22803 = n22819 ^ n22820;
  assign n22821 = ~n22820;
  assign n22824 = ~n22847;
  assign n22826 = n22853 ^ n22854;
  assign n22845 = ~n22859;
  assign n22857 = n22860 & n22779;
  assign n22809 = ~n22861;
  assign n22855 = ~n22853;
  assign n21585 = n21588 & n21553;
  assign n21490 = n22875 ^ n22876;
  assign n22877 = ~n22875;
  assign n22794 = n22803 & n19892;
  assign n22795 = ~n22803;
  assign n22771 = n22821 & n22822;
  assign n22825 = n22824 & n22799;
  assign n22815 = n22826 ^ n22827;
  assign n22796 = n22845 & n22846;
  assign n22848 = n22855 & n22856;
  assign n22781 = ~n22857;
  assign n22736 = n21490 ^ n21461;
  assign n19047 = n21490 ^ n20335;
  assign n22874 = n22877 & n22878;
  assign n22770 = ~n22794;
  assign n22785 = n22795 & n19890;
  assign n22777 = ~n22771;
  assign n22805 = n22815 & n500;
  assign n22797 = ~n22825;
  assign n22804 = ~n22815;
  assign n22823 = ~n22796;
  assign n22828 = ~n22848;
  assign n22835 = n22736 & n22849;
  assign n22836 = n19047 & n22850;
  assign n22834 = ~n22736;
  assign n19051 = ~n19047;
  assign n22862 = ~n22874;
  assign n22769 = n22770 & n22746;
  assign n22756 = ~n22785;
  assign n22772 = n22796 ^ n22797;
  assign n22800 = n22804 & n9098;
  assign n22752 = ~n22805;
  assign n22816 = n22823 & n22824;
  assign n22806 = n22828 & n22829;
  assign n22830 = n22834 & n22760;
  assign n22738 = ~n22835;
  assign n21492 = ~n22836;
  assign n22831 = n19051 & n22837;
  assign n22838 = n22862 & n22863;
  assign n22755 = ~n22769;
  assign n22745 = n22756 & n22770;
  assign n22732 = n22771 ^ n22772;
  assign n22724 = n22772 & n22777;
  assign n22774 = ~n22800;
  assign n22778 = n22806 ^ n22807;
  assign n22798 = ~n22816;
  assign n22808 = ~n22806;
  assign n22762 = ~n22830;
  assign n21527 = ~n22831;
  assign n21365 = n22838 ^ n22839;
  assign n22840 = ~n22838;
  assign n18772 = n22745 ^ n22746;
  assign n22731 = n22755 & n22756;
  assign n22748 = n22732 & n19794;
  assign n22747 = ~n22732;
  assign n22775 = n22774 & n22752;
  assign n22764 = n22778 ^ n22779;
  assign n22749 = n22798 & n22799;
  assign n22801 = n22808 & n22809;
  assign n22810 = n21527 & n21492;
  assign n22708 = n21365 ^ n21289;
  assign n19036 = n21365 ^ n20247;
  assign n22832 = n22840 & n22841;
  assign n22697 = n22722 ^ n18772;
  assign n22699 = n22731 ^ n22732;
  assign n18774 = ~n18772;
  assign n22733 = ~n22731;
  assign n22740 = n22747 & n19797;
  assign n22734 = ~n22748;
  assign n22758 = n22764 & n499;
  assign n22750 = ~n22775;
  assign n22757 = ~n22764;
  assign n22773 = ~n22749;
  assign n22780 = ~n22801;
  assign n22787 = n22708 & n22802;
  assign n22788 = n19036 & n21414;
  assign n21525 = ~n22810;
  assign n22786 = ~n22708;
  assign n19045 = ~n19036;
  assign n22817 = ~n22832;
  assign n22690 = n22697 & n22698;
  assign n18628 = n22699 ^ n19794;
  assign n22688 = ~n22697;
  assign n22723 = n22733 & n22734;
  assign n22701 = ~n22740;
  assign n22725 = n22749 ^ n22750;
  assign n22753 = n22757 & n9053;
  assign n22694 = ~n22758;
  assign n22765 = n22773 & n22774;
  assign n22759 = n22780 & n22781;
  assign n22782 = n22786 & n22677;
  assign n22710 = ~n22787;
  assign n21449 = ~n22788;
  assign n22783 = n19045 & n22789;
  assign n22790 = n22817 & n22818;
  assign n22682 = n22688 & n22689;
  assign n22632 = ~n22690;
  assign n18636 = ~n18628;
  assign n22700 = ~n22723;
  assign n22702 = n22724 ^ n22725;
  assign n22673 = n22725 & n22724;
  assign n22727 = ~n22753;
  assign n22735 = n22759 ^ n22760;
  assign n22751 = ~n22765;
  assign n22761 = ~n22759;
  assign n22679 = ~n22782;
  assign n21416 = ~n22783;
  assign n18920 = n22790 ^ n22791;
  assign n22792 = ~n22790;
  assign n22553 = n22664 ^ n18636;
  assign n22665 = ~n22682;
  assign n22634 = n22700 & n22701;
  assign n22691 = n22702 & n19768;
  assign n22692 = ~n22702;
  assign n22703 = n22727 & n22694;
  assign n22713 = n22735 ^ n22736;
  assign n22704 = n22751 & n22752;
  assign n22754 = n22761 & n22762;
  assign n21297 = n20269 ^ n18920;
  assign n22766 = n18920 & n22776;
  assign n18998 = ~n18920;
  assign n22784 = n22792 & n22793;
  assign n22626 = n22553 & n22589;
  assign n22627 = ~n22553;
  assign n22654 = n22665 & n22630;
  assign n22629 = n22665 & n22632;
  assign n22666 = ~n22634;
  assign n22636 = ~n22691;
  assign n22683 = n22692 & n19751;
  assign n22674 = n22703 ^ n22704;
  assign n22706 = n22713 & n498;
  assign n22705 = ~n22713;
  assign n22726 = ~n22704;
  assign n22728 = n21297 ^ n21272;
  assign n22737 = ~n22754;
  assign n22763 = n18998 & n21375;
  assign n21340 = ~n22766;
  assign n22767 = ~n22784;
  assign n22564 = ~n22626;
  assign n22620 = n22627 & n22628;
  assign n22613 = n22629 ^ n22630;
  assign n22631 = ~n22654;
  assign n22602 = n22673 ^ n22674;
  assign n22667 = ~n22683;
  assign n22675 = ~n22674;
  assign n22695 = n22705 & n9015;
  assign n22641 = ~n22706;
  assign n22714 = n22726 & n22727;
  assign n22715 = n22728 & n22729;
  assign n22707 = n22737 & n22738;
  assign n22716 = ~n22728;
  assign n21377 = ~n22763;
  assign n22742 = n22767 & n22768;
  assign n22599 = n22613 & n70;
  assign n22597 = ~n22620;
  assign n22598 = ~n22613;
  assign n22621 = n22631 & n22632;
  assign n22644 = n22602 & n19738;
  assign n22655 = n22666 & n22667;
  assign n22633 = n22667 & n22636;
  assign n22645 = ~n22602;
  assign n22605 = n22675 & n22673;
  assign n22669 = ~n22695;
  assign n22676 = n22707 ^ n22708;
  assign n22693 = ~n22714;
  assign n22617 = ~n22715;
  assign n22711 = n22716 & n22717;
  assign n22709 = ~n22707;
  assign n18970 = n22741 ^ n22742;
  assign n22743 = ~n22742;
  assign n22587 = n22598 & n3685;
  assign n22534 = ~n22599;
  assign n22588 = ~n22621;
  assign n18582 = n22633 ^ n22634;
  assign n22604 = ~n22644;
  assign n22637 = n22645 & n19744;
  assign n22635 = ~n22655;
  assign n22608 = ~n22605;
  assign n22670 = n22669 & n22641;
  assign n22656 = n22676 ^ n22677;
  assign n22638 = n22693 & n22694;
  assign n22696 = n22709 & n22710;
  assign n22651 = ~n22711;
  assign n21264 = n18970 ^ n20230;
  assign n22718 = n18970 & n22730;
  assign n18978 = ~n18970;
  assign n22739 = n22743 & n22744;
  assign n22565 = ~n22587;
  assign n22552 = n22588 ^ n22589;
  assign n22586 = n22597 & n22588;
  assign n22528 = n22600 ^ n18582;
  assign n18520 = ~n18582;
  assign n22601 = n22635 & n22636;
  assign n22570 = ~n22637;
  assign n22647 = n22656 & n497;
  assign n22639 = ~n22670;
  assign n22646 = ~n22656;
  assign n22668 = ~n22638;
  assign n22648 = n22651 & n22617;
  assign n22582 = n21264 ^ n21083;
  assign n22678 = ~n22696;
  assign n21303 = ~n22718;
  assign n22712 = n18978 & n22719;
  assign n22720 = ~n22739;
  assign n22526 = n22552 ^ n22553;
  assign n22554 = n22565 & n22530;
  assign n22529 = n22565 & n22534;
  assign n22567 = n22528 & n22577;
  assign n22563 = ~n22586;
  assign n22566 = ~n22528;
  assign n22568 = n22601 ^ n22602;
  assign n22603 = ~n22601;
  assign n22606 = n22638 ^ n22639;
  assign n22642 = n22646 & n8981;
  assign n22574 = ~n22647;
  assign n22657 = n22668 & n22669;
  assign n22659 = n22582 & n22671;
  assign n22649 = n22678 & n22679;
  assign n22658 = ~n22582;
  assign n21268 = ~n22712;
  assign n22685 = n22720 & n22721;
  assign n22516 = n22526 & n69;
  assign n22486 = n22529 ^ n22530;
  assign n22515 = ~n22526;
  assign n22533 = ~n22554;
  assign n22527 = n22563 & n22564;
  assign n22555 = n22566 & n22488;
  assign n22532 = ~n22567;
  assign n18532 = n19744 ^ n22568;
  assign n22590 = n22603 & n22604;
  assign n22578 = n22605 ^ n22606;
  assign n22607 = ~n22606;
  assign n22610 = ~n22642;
  assign n22500 = n22648 ^ n22649;
  assign n22640 = ~n22657;
  assign n22652 = n22658 & n22547;
  assign n22584 = ~n22659;
  assign n22650 = ~n22649;
  assign n22680 = n21303 & n21268;
  assign n18912 = n22684 ^ n22685;
  assign n22686 = ~n22685;
  assign n21274 = n22486 ^ n21298;
  assign n21266 = n22486 ^ n21310;
  assign n22385 = n22486 & n21298;
  assign n22505 = n22515 & n3604;
  assign n22438 = ~n22516;
  assign n22487 = n22527 ^ n22528;
  assign n22426 = n22533 & n22534;
  assign n22412 = n22535 ^ n18532;
  assign n22531 = ~n22527;
  assign n22490 = ~n22555;
  assign n18525 = ~n18532;
  assign n22571 = n22578 & n19699;
  assign n22569 = ~n22590;
  assign n22572 = ~n22578;
  assign n22542 = n22607 & n22608;
  assign n22579 = n22610 & n22574;
  assign n22614 = n22500 & n8944;
  assign n22580 = n22640 & n22641;
  assign n22615 = ~n22500;
  assign n22643 = n22650 & n22651;
  assign n22549 = ~n22652;
  assign n21177 = n18912 ^ n20173;
  assign n22661 = n18912 & n22672;
  assign n21301 = ~n22680;
  assign n18917 = ~n18912;
  assign n22681 = n22686 & n22687;
  assign n22400 = n22487 ^ n22488;
  assign n22389 = ~n22385;
  assign n22479 = ~n22505;
  assign n22491 = n22412 & n22455;
  assign n22480 = ~n22426;
  assign n22492 = ~n22412;
  assign n22517 = n22531 & n22532;
  assign n22495 = n22569 & n22570;
  assign n22536 = ~n22571;
  assign n22556 = n22572 & n19703;
  assign n22543 = n22579 ^ n22580;
  assign n22545 = ~n22542;
  assign n22540 = ~n22614;
  assign n22611 = n22615 & n496;
  assign n22609 = ~n22580;
  assign n22511 = n21177 ^ n20996;
  assign n22616 = ~n22643;
  assign n22653 = n18917 & n22660;
  assign n21223 = ~n22661;
  assign n22662 = ~n22681;
  assign n22453 = n22400 & n68;
  assign n22452 = ~n22400;
  assign n22471 = n22479 & n22480;
  assign n22472 = n22479 & n22438;
  assign n22414 = ~n22491;
  assign n22481 = n22492 & n22493;
  assign n22489 = ~n22517;
  assign n22518 = n22542 ^ n22543;
  assign n22537 = ~n22495;
  assign n22497 = ~n22556;
  assign n22544 = ~n22543;
  assign n22591 = n22609 & n22610;
  assign n22502 = ~n22611;
  assign n22592 = n22511 & n22612;
  assign n22581 = n22616 & n22617;
  assign n22593 = ~n22511;
  assign n21180 = ~n22653;
  assign n22622 = n22662 & n22663;
  assign n22436 = n22452 & n3531;
  assign n22362 = ~n22453;
  assign n22437 = ~n22471;
  assign n22427 = ~n22472;
  assign n22457 = ~n22481;
  assign n22454 = n22489 & n22490;
  assign n22506 = n22518 & n19663;
  assign n22519 = n22536 & n22537;
  assign n22494 = n22497 & n22536;
  assign n22507 = ~n22518;
  assign n22458 = n22544 & n22545;
  assign n22546 = n22581 ^ n22582;
  assign n22573 = ~n22591;
  assign n22513 = ~n22592;
  assign n22585 = n22593 & n22474;
  assign n22583 = ~n22581;
  assign n22618 = n21223 & n21180;
  assign n22594 = n22622 ^ n22623;
  assign n22624 = ~n22622;
  assign n21092 = ~n22594;
  assign n22386 = n22426 ^ n22427;
  assign n22397 = ~n22436;
  assign n22399 = n22437 & n22438;
  assign n22411 = n22454 ^ n22455;
  assign n22456 = ~n22454;
  assign n22467 = n21092 ^ n21055;
  assign n18454 = n22494 ^ n22495;
  assign n22422 = ~n22506;
  assign n22498 = n22507 & n19651;
  assign n22496 = ~n22519;
  assign n22463 = ~n22458;
  assign n22520 = n22546 ^ n22547;
  assign n22538 = n22573 & n22574;
  assign n22575 = n22583 & n22584;
  assign n22476 = ~n22585;
  assign n18890 = n22594 ^ n20148;
  assign n21221 = ~n22618;
  assign n22619 = n22624 & n22625;
  assign n20225 = n22385 ^ n22386;
  assign n22360 = n22399 ^ n22400;
  assign n22323 = n22411 ^ n22412;
  assign n22388 = ~n22386;
  assign n22398 = ~n22399;
  assign n22439 = n22456 & n22457;
  assign n22445 = n22467 & n22468;
  assign n22443 = ~n22467;
  assign n18491 = ~n18454;
  assign n22419 = n22496 & n22497;
  assign n22461 = ~n22498;
  assign n22509 = n22520 & n511;
  assign n22499 = n496 ^ n22538;
  assign n22508 = ~n22520;
  assign n22539 = ~n22538;
  assign n22548 = ~n22575;
  assign n22557 = n18890 & n22576;
  assign n18883 = ~n18890;
  assign n22595 = ~n22619;
  assign n22319 = n68 ^ n22360;
  assign n21190 = ~n20225;
  assign n22376 = n22323 & n3431;
  assign n22318 = n22388 & n22389;
  assign n22387 = n22397 & n22398;
  assign n22377 = ~n22323;
  assign n22413 = ~n22439;
  assign n22415 = n22440 ^ n18491;
  assign n22433 = n22443 & n22444;
  assign n22370 = ~n22445;
  assign n22464 = n22461 & n22422;
  assign n22460 = ~n22419;
  assign n22459 = n22499 ^ n22500;
  assign n22503 = n22508 & n8895;
  assign n22424 = ~n22509;
  assign n22521 = n22539 & n22540;
  assign n22510 = n22548 & n22549;
  assign n21096 = ~n22557;
  assign n22550 = n18883 & n22558;
  assign n22559 = n22595 & n22596;
  assign n21093 = n22318 ^ n22319;
  assign n22320 = ~n22319;
  assign n22324 = ~n22376;
  assign n22363 = n22377 & n67;
  assign n22321 = ~n22318;
  assign n22361 = ~n22387;
  assign n22329 = n22413 & n22414;
  assign n22401 = n22415 & n22416;
  assign n22402 = ~n22415;
  assign n22405 = ~n22433;
  assign n22428 = n22458 ^ n22459;
  assign n22441 = n22460 & n22461;
  assign n22420 = ~n22464;
  assign n22462 = ~n22459;
  assign n22466 = ~n22503;
  assign n22473 = n22510 ^ n22511;
  assign n22501 = ~n22521;
  assign n22512 = ~n22510;
  assign n21140 = ~n22550;
  assign n18833 = n22559 ^ n22560;
  assign n22561 = ~n22559;
  assign n21108 = ~n21093;
  assign n22238 = n22320 & n22321;
  assign n22322 = n22361 & n22362;
  assign n22283 = ~n22363;
  assign n22364 = ~n22329;
  assign n22327 = ~n22401;
  assign n22390 = n22402 & n22403;
  assign n22394 = n22370 & n22405;
  assign n18474 = n22419 ^ n22420;
  assign n22417 = n22428 & n19601;
  assign n22418 = ~n22428;
  assign n22421 = ~n22441;
  assign n22391 = n22462 & n22463;
  assign n22429 = n22466 & n22424;
  assign n22349 = n22473 ^ n22474;
  assign n22430 = n22501 & n22502;
  assign n22504 = n22512 & n22513;
  assign n21137 = n21140 & n21096;
  assign n20999 = n18833 ^ n20032;
  assign n22522 = n18833 & n22541;
  assign n18758 = ~n18833;
  assign n22551 = n22561 & n22562;
  assign n22281 = n22322 ^ n22323;
  assign n22325 = ~n22322;
  assign n22245 = n22378 ^ n18474;
  assign n22365 = ~n22390;
  assign n22358 = ~n22394;
  assign n18464 = ~n18474;
  assign n22379 = ~n22417;
  assign n22404 = n22418 & n19645;
  assign n22331 = n22421 & n22422;
  assign n22392 = n22429 ^ n22430;
  assign n22432 = n22349 & n510;
  assign n22431 = ~n22349;
  assign n22465 = ~n22430;
  assign n22293 = n20999 ^ n20962;
  assign n22475 = ~n22504;
  assign n21012 = ~n22522;
  assign n22514 = n18758 & n22523;
  assign n22524 = ~n22551;
  assign n22239 = n67 ^ n22281;
  assign n22312 = n22324 & n22325;
  assign n22344 = n22245 & n22354;
  assign n22353 = n22364 & n22365;
  assign n22328 = n22365 & n22327;
  assign n22343 = ~n22245;
  assign n22302 = n22391 ^ n22392;
  assign n22346 = ~n22404;
  assign n22380 = ~n22331;
  assign n22305 = n22392 & n22391;
  assign n22425 = n22431 & n8851;
  assign n22351 = ~n22432;
  assign n22442 = n22465 & n22466;
  assign n22446 = n22293 & n22469;
  assign n22357 = n22475 & n22476;
  assign n22447 = ~n22293;
  assign n21060 = ~n22514;
  assign n22482 = n22524 & n22525;
  assign n21023 = n22238 ^ n22239;
  assign n22166 = n22239 & n22238;
  assign n22282 = ~n22312;
  assign n22241 = n22328 ^ n22329;
  assign n22330 = n22343 & n22285;
  assign n22247 = ~n22344;
  assign n22326 = ~n22353;
  assign n22269 = n22357 ^ n22358;
  assign n22355 = n22302 & n19581;
  assign n22366 = n22379 & n22380;
  assign n22367 = n22379 & n22346;
  assign n22356 = ~n22302;
  assign n22383 = ~n22425;
  assign n22423 = ~n22442;
  assign n22295 = ~n22446;
  assign n22434 = n22447 & n22334;
  assign n22406 = ~n22357;
  assign n22477 = n21060 & n21012;
  assign n18808 = n22482 ^ n22483;
  assign n22484 = ~n22482;
  assign n21010 = ~n21023;
  assign n22169 = ~n22166;
  assign n22240 = n22282 & n22283;
  assign n22288 = n22241 & n3384;
  assign n22289 = ~n22241;
  assign n22284 = n22326 & n22327;
  assign n22287 = ~n22330;
  assign n22314 = n22269 & n509;
  assign n22313 = ~n22269;
  assign n22304 = ~n22355;
  assign n22347 = n22356 & n19550;
  assign n22345 = ~n22366;
  assign n22332 = ~n22367;
  assign n22393 = n22405 & n22406;
  assign n22381 = n22423 & n22424;
  assign n22336 = ~n22434;
  assign n20931 = n18808 ^ n20011;
  assign n22448 = n18808 & n22470;
  assign n21058 = ~n22477;
  assign n18801 = ~n18808;
  assign n22478 = n22484 & n22485;
  assign n22203 = n22240 ^ n22241;
  assign n22242 = ~n22240;
  assign n22244 = n22284 ^ n22285;
  assign n22243 = ~n22288;
  assign n22275 = n22289 & n66;
  assign n22286 = ~n22284;
  assign n22308 = n22313 & n8797;
  assign n22232 = ~n22314;
  assign n18406 = n22331 ^ n22332;
  assign n22301 = n22345 & n22346;
  assign n22265 = ~n22347;
  assign n22348 = n510 ^ n22381;
  assign n22369 = ~n22393;
  assign n22382 = ~n22381;
  assign n22215 = n20931 ^ n20787;
  assign n20934 = ~n22448;
  assign n22435 = n18801 & n22449;
  assign n22450 = ~n22478;
  assign n22167 = n66 ^ n22203;
  assign n22229 = n22242 & n22243;
  assign n22222 = n22244 ^ n22245;
  assign n22205 = ~n22275;
  assign n22274 = n22286 & n22287;
  assign n22173 = n22290 ^ n18406;
  assign n22263 = n22301 ^ n22302;
  assign n22277 = ~n22308;
  assign n18398 = ~n18406;
  assign n22303 = ~n22301;
  assign n22306 = n22348 ^ n22349;
  assign n22333 = n22369 & n22370;
  assign n22368 = n22382 & n22383;
  assign n22371 = n22215 & n22384;
  assign n22372 = ~n22215;
  assign n20977 = ~n22435;
  assign n22407 = n22450 & n22451;
  assign n20102 = n22166 ^ n22167;
  assign n22168 = ~n22167;
  assign n22207 = n22222 & n65;
  assign n22204 = ~n22229;
  assign n22206 = ~n22222;
  assign n22248 = n22173 & n22262;
  assign n18363 = n22263 ^ n19550;
  assign n22246 = ~n22274;
  assign n22249 = ~n22173;
  assign n22291 = n22303 & n22304;
  assign n22276 = n22305 ^ n22306;
  assign n22226 = n22306 & n22305;
  assign n22292 = n22333 ^ n22334;
  assign n22335 = ~n22333;
  assign n22350 = ~n22368;
  assign n22217 = ~n22371;
  assign n22359 = n22372 & n22256;
  assign n22395 = n20977 & n20934;
  assign n22373 = n22407 ^ n22408;
  assign n22409 = ~n22407;
  assign n20948 = ~n20102;
  assign n22107 = n22168 & n22169;
  assign n22143 = n22204 & n22205;
  assign n22195 = n22206 & n3342;
  assign n22145 = ~n22207;
  assign n22135 = n22223 ^ n18363;
  assign n22208 = n22246 & n22247;
  assign n22176 = ~n22248;
  assign n22230 = n22249 & n22209;
  assign n18361 = ~n18363;
  assign n22266 = n22276 & n19527;
  assign n22264 = ~n22291;
  assign n22267 = ~n22276;
  assign n22161 = n22292 ^ n22293;
  assign n22315 = n22335 & n22336;
  assign n22307 = n22350 & n22351;
  assign n22258 = ~n22359;
  assign n18669 = n20009 ^ n22373;
  assign n20975 = ~n22395;
  assign n22396 = n22409 & n22410;
  assign n22170 = ~n22143;
  assign n22171 = ~n22195;
  assign n22187 = n22135 & n22196;
  assign n22188 = ~n22135;
  assign n22172 = n22208 ^ n22209;
  assign n22210 = ~n22208;
  assign n22211 = ~n22230;
  assign n22177 = n22264 & n22265;
  assign n22224 = ~n22266;
  assign n22250 = n22267 & n19529;
  assign n22252 = n22161 & n508;
  assign n22251 = ~n22161;
  assign n22268 = n509 ^ n22307;
  assign n22294 = ~n22315;
  assign n22278 = ~n22307;
  assign n20833 = n20009 ^ n18669;
  assign n22337 = n18669 & n22352;
  assign n18719 = ~n18669;
  assign n22374 = ~n22396;
  assign n22158 = n22170 & n22171;
  assign n22142 = n22171 & n22145;
  assign n22110 = n22172 ^ n22173;
  assign n22148 = ~n22187;
  assign n22174 = n22188 & n22098;
  assign n22197 = n22210 & n22211;
  assign n22225 = ~n22177;
  assign n22190 = ~n22250;
  assign n22233 = n22251 & n8745;
  assign n22163 = ~n22252;
  assign n22227 = n22268 ^ n22269;
  assign n22270 = n22277 & n22278;
  assign n22183 = n20833 ^ n20692;
  assign n22255 = n22294 & n22295;
  assign n20846 = ~n22337;
  assign n22316 = n18719 & n22338;
  assign n22340 = n22374 & n22375;
  assign n22108 = n22142 ^ n22143;
  assign n22147 = n22110 & n64;
  assign n22144 = ~n22158;
  assign n22146 = ~n22110;
  assign n22114 = ~n22174;
  assign n22175 = ~n22197;
  assign n22212 = n22224 & n22225;
  assign n22213 = n22224 & n22190;
  assign n22198 = n22226 ^ n22227;
  assign n22136 = n22227 & n22226;
  assign n22200 = ~n22233;
  assign n22214 = n22255 ^ n22256;
  assign n22231 = ~n22270;
  assign n22254 = n22183 & n22271;
  assign n22253 = ~n22183;
  assign n22257 = ~n22255;
  assign n20890 = ~n22316;
  assign n18619 = n22339 ^ n22340;
  assign n22342 = n22340 & n22299;
  assign n22341 = ~n22340;
  assign n20062 = n22107 ^ n22108;
  assign n22040 = n22108 & n22107;
  assign n22109 = n22144 & n22145;
  assign n22132 = n22146 & n3315;
  assign n22079 = ~n22147;
  assign n22159 = n22175 & n22176;
  assign n22192 = n22198 & n19511;
  assign n22189 = ~n22212;
  assign n22178 = ~n22213;
  assign n22191 = ~n22198;
  assign n22193 = n22214 ^ n22215;
  assign n22199 = n22231 & n22232;
  assign n22234 = n22253 & n22153;
  assign n22185 = ~n22254;
  assign n22235 = n22257 & n22258;
  assign n20887 = n20890 & n20846;
  assign n20751 = n18619 ^ n19981;
  assign n22296 = n18619 & n22309;
  assign n18617 = ~n18619;
  assign n22317 = n22341 & n22311;
  assign n22310 = ~n22342;
  assign n20844 = ~n20062;
  assign n22043 = ~n22040;
  assign n22077 = n22109 ^ n22110;
  assign n22111 = ~n22109;
  assign n22112 = ~n22132;
  assign n22134 = ~n22159;
  assign n18322 = n22177 ^ n22178;
  assign n22117 = n22189 & n22190;
  assign n22179 = n22191 & n19452;
  assign n22157 = ~n22192;
  assign n22181 = n22193 & n507;
  assign n22160 = n508 ^ n22199;
  assign n22180 = ~n22193;
  assign n22201 = ~n22199;
  assign n22155 = ~n22234;
  assign n22216 = ~n22235;
  assign n22090 = n20751 ^ n20722;
  assign n20755 = ~n22296;
  assign n22279 = n18617 & n22297;
  assign n22300 = n22310 & n22311;
  assign n22298 = ~n22317;
  assign n22041 = n64 ^ n22077;
  assign n22096 = n22111 & n22112;
  assign n22097 = n22134 ^ n22135;
  assign n22133 = n22134 & n22148;
  assign n22045 = n18322 ^ n22149;
  assign n18319 = ~n18322;
  assign n22137 = n22160 ^ n22161;
  assign n22156 = ~n22117;
  assign n22129 = ~n22179;
  assign n22164 = n22180 & n8665;
  assign n22103 = ~n22181;
  assign n22194 = n22200 & n22201;
  assign n22182 = n22216 & n22217;
  assign n22218 = n22090 & n22228;
  assign n22219 = ~n22090;
  assign n20771 = ~n22279;
  assign n22280 = n22298 & n22299;
  assign n22272 = ~n22300;
  assign n20769 = n22040 ^ n22041;
  assign n22042 = ~n22041;
  assign n22078 = ~n22096;
  assign n22047 = n22097 ^ n22098;
  assign n22115 = n22045 & n22127;
  assign n22113 = ~n22133;
  assign n22116 = ~n22045;
  assign n22094 = n22136 ^ n22137;
  assign n22087 = n22137 & n22136;
  assign n22150 = n22156 & n22157;
  assign n22151 = n22157 & n22129;
  assign n22139 = ~n22164;
  assign n22152 = n22182 ^ n22183;
  assign n22162 = ~n22194;
  assign n22184 = ~n22182;
  assign n22092 = ~n22218;
  assign n22202 = n22219 & n22124;
  assign n22236 = n20771 & n20755;
  assign n22261 = n22272 & n22273;
  assign n22259 = ~n22280;
  assign n20752 = ~n20769;
  assign n20600 = n22042 & n22043;
  assign n22046 = n22078 & n22079;
  assign n22070 = n22047 & n3280;
  assign n22071 = ~n22047;
  assign n22080 = n22113 & n22114;
  assign n22051 = ~n22115;
  assign n22099 = n22116 & n22081;
  assign n22100 = n22094 & n19487;
  assign n22101 = ~n22094;
  assign n22128 = ~n22150;
  assign n22118 = ~n22151;
  assign n22119 = n22139 & n22103;
  assign n22130 = n22152 ^ n22153;
  assign n22120 = n22162 & n22163;
  assign n22165 = n22184 & n22185;
  assign n22126 = ~n22202;
  assign n20800 = ~n22236;
  assign n22237 = n22259 & n22260;
  assign n22221 = ~n22261;
  assign n22019 = n22046 ^ n22047;
  assign n22048 = ~n22046;
  assign n22049 = ~n22070;
  assign n22063 = n22071 & n79;
  assign n22044 = n22080 ^ n22081;
  assign n22082 = ~n22080;
  assign n22083 = ~n22099;
  assign n22085 = ~n22100;
  assign n22095 = n22101 & n19494;
  assign n18233 = n22117 ^ n22118;
  assign n22088 = n22119 ^ n22120;
  assign n22093 = n22128 & n22129;
  assign n22122 = n22130 & n506;
  assign n22121 = ~n22130;
  assign n22138 = ~n22120;
  assign n22154 = ~n22165;
  assign n22220 = ~n22237;
  assign n20636 = n79 ^ n22019;
  assign n22030 = n22044 ^ n22045;
  assign n22032 = n22048 & n22049;
  assign n22023 = ~n22063;
  assign n22072 = n22082 & n22083;
  assign n22064 = n22084 ^ n18233;
  assign n22067 = n22087 ^ n22088;
  assign n22066 = n22093 ^ n22094;
  assign n22056 = ~n22095;
  assign n22014 = n22088 & n22087;
  assign n18264 = ~n18233;
  assign n22086 = ~n22093;
  assign n22104 = n22121 & n8632;
  assign n22038 = ~n22122;
  assign n22131 = n22138 & n22139;
  assign n22123 = n22154 & n22155;
  assign n18647 = n22220 & n22221;
  assign n21932 = n20636 & n20600;
  assign n22021 = n22030 & n78;
  assign n22020 = ~n22030;
  assign n22022 = ~n22032;
  assign n22052 = n22064 & n22065;
  assign n18252 = n19494 ^ n22066;
  assign n22057 = n22067 & n19399;
  assign n22050 = ~n22072;
  assign n22053 = ~n22064;
  assign n22058 = ~n22067;
  assign n22073 = n22085 & n22086;
  assign n22028 = ~n22014;
  assign n22075 = ~n22104;
  assign n22089 = n22123 ^ n22124;
  assign n22102 = ~n22131;
  assign n22125 = ~n22123;
  assign n20708 = n18647 ^ n22186;
  assign n19963 = ~n18647;
  assign n21935 = ~n21932;
  assign n22009 = n22020 & n3229;
  assign n21969 = ~n22021;
  assign n21957 = n22022 & n22023;
  assign n21948 = n22031 ^ n18252;
  assign n22001 = n22050 & n22051;
  assign n21998 = ~n22052;
  assign n22033 = n22053 & n22054;
  assign n18248 = ~n18252;
  assign n22026 = ~n22057;
  assign n22034 = n22058 & n19434;
  assign n22055 = ~n22073;
  assign n22076 = n22075 & n22038;
  assign n22068 = n22089 ^ n22090;
  assign n22035 = n22102 & n22103;
  assign n22105 = n22125 & n22126;
  assign n22140 = n19963 ^ n19931;
  assign n20724 = ~n20708;
  assign n21996 = ~n22009;
  assign n21995 = ~n21957;
  assign n22006 = n21948 & n22010;
  assign n22007 = ~n21948;
  assign n22024 = ~n22001;
  assign n22025 = ~n22033;
  assign n22003 = ~n22034;
  assign n21986 = n22055 & n22056;
  assign n22060 = n22068 & n505;
  assign n22036 = ~n22076;
  assign n22059 = ~n22068;
  assign n22074 = ~n22035;
  assign n22091 = ~n22105;
  assign n20629 = n22140 ^ n22141;
  assign n21984 = n21995 & n21996;
  assign n21985 = n21996 & n21969;
  assign n21950 = ~n22006;
  assign n21999 = n22007 & n21971;
  assign n22011 = n22024 & n22025;
  assign n22000 = n22025 & n21998;
  assign n22013 = n22003 & n22026;
  assign n22027 = ~n21986;
  assign n22015 = n22035 ^ n22036;
  assign n22039 = n22059 & n8583;
  assign n21993 = ~n22060;
  assign n22069 = n22074 & n22075;
  assign n22061 = n22091 & n22092;
  assign n22062 = n20629 ^ n22106;
  assign n21968 = ~n21984;
  assign n21958 = ~n21985;
  assign n21972 = ~n21999;
  assign n21922 = n22000 ^ n22001;
  assign n21997 = ~n22011;
  assign n21987 = ~n22013;
  assign n21977 = n22014 ^ n22015;
  assign n22012 = n22026 & n22027;
  assign n21963 = n22015 & n22028;
  assign n22005 = ~n22039;
  assign n22029 = n22061 ^ n22062;
  assign n22037 = ~n22069;
  assign n21933 = n21957 ^ n21958;
  assign n21944 = n21968 & n21969;
  assign n21974 = n21922 & n3182;
  assign n21975 = ~n21922;
  assign n18174 = n21986 ^ n21987;
  assign n21970 = n21997 & n21998;
  assign n21989 = n21977 & n19418;
  assign n21988 = ~n21977;
  assign n22002 = ~n22012;
  assign n22018 = n22005 & n21993;
  assign n21966 = n504 ^ n22029;
  assign n21991 = n22037 & n22038;
  assign n19918 = n21932 ^ n21933;
  assign n21921 = n77 ^ n21944;
  assign n21934 = ~n21933;
  assign n21945 = ~n21944;
  assign n21952 = n21961 ^ n18174;
  assign n21947 = n21970 ^ n21971;
  assign n21946 = ~n21974;
  assign n21960 = n21975 & n77;
  assign n18201 = ~n18174;
  assign n21973 = ~n21970;
  assign n21982 = n21988 & n19339;
  assign n21979 = ~n21989;
  assign n21976 = n22002 & n22003;
  assign n21990 = ~n22018;
  assign n21981 = ~n21966;
  assign n22017 = n21993 & n21991;
  assign n22016 = ~n21991;
  assign n21901 = n21921 ^ n21922;
  assign n19947 = ~n19918;
  assign n21900 = n21934 & n21935;
  assign n21936 = n21945 & n21946;
  assign n21929 = n21947 ^ n21948;
  assign n21939 = n21952 & n21953;
  assign n21937 = ~n21952;
  assign n21924 = ~n21960;
  assign n21959 = n21972 & n21973;
  assign n21951 = n21976 ^ n21977;
  assign n21955 = ~n21982;
  assign n21978 = ~n21976;
  assign n21964 = n21990 ^ n21991;
  assign n22008 = n22005 & n22016;
  assign n22004 = ~n22017;
  assign n21873 = n21900 ^ n21901;
  assign n17799 = n18803 ^ n19947;
  assign n19935 = n19947 & n18803;
  assign n21902 = ~n21901;
  assign n21926 = n21929 & n76;
  assign n21923 = ~n21936;
  assign n21925 = ~n21929;
  assign n21930 = n21937 & n21938;
  assign n21894 = ~n21939;
  assign n18186 = n21951 ^ n19339;
  assign n21949 = ~n21959;
  assign n21908 = n21963 ^ n21964;
  assign n21962 = n21978 & n21979;
  assign n21919 = n21964 & n21963;
  assign n21994 = n22004 & n22005;
  assign n21992 = ~n22008;
  assign n21853 = n19935 ^ n21873;
  assign n21854 = n21902 & n21900;
  assign n21891 = n19935 & n18772;
  assign n19916 = ~n17799;
  assign n19900 = ~n19935;
  assign n21883 = n21923 & n21924;
  assign n21914 = n21925 & n3147;
  assign n21885 = ~n21926;
  assign n21847 = n21927 ^ n18186;
  assign n21915 = ~n21930;
  assign n18179 = ~n18186;
  assign n21888 = n21949 & n21950;
  assign n21941 = n21908 & n19354;
  assign n21940 = ~n21908;
  assign n21954 = ~n21962;
  assign n21983 = n21992 & n21993;
  assign n21980 = ~n21994;
  assign n17672 = n21853 ^ n18774;
  assign n21862 = n19916 & n19910;
  assign n21887 = n19900 & n18774;
  assign n21857 = ~n21854;
  assign n21845 = ~n21891;
  assign n21906 = n21847 & n21910;
  assign n21903 = ~n21883;
  assign n21904 = ~n21914;
  assign n21905 = ~n21847;
  assign n21912 = n21915 & n21894;
  assign n21916 = ~n21888;
  assign n21931 = n21940 & n19346;
  assign n21897 = ~n21941;
  assign n21928 = n21954 & n21955;
  assign n21967 = n21980 & n21981;
  assign n21965 = ~n21983;
  assign n21810 = n17672 & n19890;
  assign n17679 = ~n17672;
  assign n21842 = n21862 ^ n21863;
  assign n21836 = n21862 ^ n21864;
  assign n21874 = ~n21887;
  assign n21892 = n21903 & n21904;
  assign n21882 = n21904 & n21885;
  assign n21895 = n21905 & n21876;
  assign n21849 = ~n21906;
  assign n21889 = ~n21912;
  assign n21911 = n21915 & n21916;
  assign n21907 = n21928 ^ n19346;
  assign n21918 = ~n21931;
  assign n21917 = ~n21928;
  assign n21956 = n21965 & n21966;
  assign n21942 = ~n21967;
  assign n21787 = n21810 ^ n18774;
  assign n19725 = n7 ^ n21836;
  assign n21786 = n21842 & n21843;
  assign n21837 = ~n21836;
  assign n21865 = n21873 & n21874;
  assign n21855 = n21882 ^ n21883;
  assign n21879 = n21888 ^ n21889;
  assign n21884 = ~n21892;
  assign n21877 = ~n21895;
  assign n18077 = n21907 ^ n21908;
  assign n21893 = ~n21911;
  assign n21913 = n21917 & n21918;
  assign n21943 = ~n21956;
  assign n21752 = n21786 ^ n21787;
  assign n21820 = n21786 & n21753;
  assign n21484 = ~n19725;
  assign n21818 = ~n21786;
  assign n21653 = n21837 & n7;
  assign n21796 = n21854 ^ n21855;
  assign n21844 = ~n21865;
  assign n21856 = ~n21855;
  assign n21870 = n21879 & n75;
  assign n21808 = n21884 & n21885;
  assign n21866 = n21886 ^ n18077;
  assign n21869 = ~n21879;
  assign n21875 = n21893 & n21894;
  assign n18151 = ~n18077;
  assign n21896 = ~n21913;
  assign n21920 = n21942 & n21943;
  assign n21734 = n21752 ^ n21753;
  assign n21811 = n21818 & n21819;
  assign n21767 = ~n21820;
  assign n21832 = n21796 & n18636;
  assign n21821 = n21844 & n21845;
  assign n21833 = ~n21796;
  assign n21779 = n21856 & n21857;
  assign n21858 = n21866 & n21867;
  assign n21861 = n21869 & n3117;
  assign n21813 = ~n21870;
  assign n21839 = ~n21808;
  assign n21846 = n21875 ^ n21876;
  assign n21859 = ~n21866;
  assign n21878 = ~n21875;
  assign n21840 = n21896 & n21897;
  assign n21909 = n21919 ^ n21920;
  assign n21722 = n21734 & n6;
  assign n21720 = ~n21734;
  assign n21795 = ~n21811;
  assign n21797 = n21821 ^ n18628;
  assign n21778 = ~n21832;
  assign n21822 = n21833 & n18628;
  assign n21806 = ~n21821;
  assign n21783 = ~n21779;
  assign n21755 = n21846 ^ n21847;
  assign n21802 = ~n21858;
  assign n21850 = n21859 & n21860;
  assign n21838 = ~n21861;
  assign n21868 = n21877 & n21878;
  assign n21880 = ~n21840;
  assign n21899 = n21909 & n19325;
  assign n21898 = ~n21909;
  assign n21713 = n21720 & n21721;
  assign n21655 = ~n21722;
  assign n21788 = n21787 & n21795;
  assign n17625 = n21796 ^ n21797;
  assign n21807 = ~n21822;
  assign n21824 = n21755 & n74;
  assign n21834 = n21838 & n21839;
  assign n21823 = ~n21755;
  assign n21835 = n21838 & n21813;
  assign n21825 = ~n21850;
  assign n21848 = ~n21868;
  assign n21890 = n21898 & n19331;
  assign n21881 = ~n21899;
  assign n21689 = ~n21713;
  assign n21766 = ~n21788;
  assign n17619 = ~n17625;
  assign n21798 = n21806 & n21807;
  assign n21814 = n21823 & n3056;
  assign n21758 = ~n21824;
  assign n21812 = ~n21834;
  assign n21827 = n21825 & n21802;
  assign n21809 = ~n21835;
  assign n21799 = n21848 & n21849;
  assign n21871 = n21880 & n21881;
  assign n21852 = ~n21890;
  assign n21680 = n21689 & n21653;
  assign n21652 = n21689 & n21655;
  assign n21735 = n21766 & n21767;
  assign n21740 = n17619 & n19797;
  assign n21777 = ~n21798;
  assign n21780 = n21808 ^ n21809;
  assign n21789 = n21812 & n21813;
  assign n21790 = ~n21814;
  assign n21800 = ~n21827;
  assign n21826 = ~n21799;
  assign n21851 = ~n21871;
  assign n21872 = n21852 & n21881;
  assign n21393 = n21652 ^ n21653;
  assign n21654 = ~n21680;
  assign n21702 = n21735 ^ n21736;
  assign n21703 = n21740 ^ n18628;
  assign n21739 = n21735 & n21736;
  assign n21737 = ~n21735;
  assign n21672 = n21777 & n21778;
  assign n21756 = n21779 ^ n21780;
  assign n21754 = n74 ^ n21789;
  assign n21784 = n21799 ^ n21800;
  assign n21782 = ~n21780;
  assign n21791 = ~n21789;
  assign n21815 = n21825 & n21826;
  assign n21829 = n21851 & n21852;
  assign n21841 = ~n21872;
  assign n21409 = ~n21393;
  assign n21596 = n21654 & n21655;
  assign n21679 = n21702 ^ n21703;
  assign n21723 = n21737 & n21738;
  assign n21714 = ~n21739;
  assign n21725 = n21754 ^ n21755;
  assign n21749 = n21756 & n18582;
  assign n21726 = ~n21672;
  assign n21748 = ~n21756;
  assign n21724 = n21782 & n21783;
  assign n21769 = n21784 & n73;
  assign n21781 = n21790 & n21791;
  assign n21768 = ~n21784;
  assign n21801 = ~n21815;
  assign n18021 = n21828 ^ n21829;
  assign n21830 = ~n21829;
  assign n18112 = n21840 ^ n21841;
  assign n21620 = ~n21596;
  assign n21671 = n21679 & n5;
  assign n21669 = ~n21679;
  assign n21704 = n21714 & n21703;
  assign n21682 = ~n21723;
  assign n21648 = n21724 ^ n21725;
  assign n21727 = ~n21725;
  assign n21741 = n21748 & n18520;
  assign n21716 = ~n21749;
  assign n21728 = ~n21724;
  assign n21759 = n21768 & n3021;
  assign n21695 = ~n21769;
  assign n21757 = ~n21781;
  assign n21770 = n21801 & n21802;
  assign n21743 = n18112 ^ n21816;
  assign n18055 = ~n18021;
  assign n21817 = n21830 & n21831;
  assign n18106 = ~n18112;
  assign n21656 = n21669 & n21670;
  assign n21599 = ~n21671;
  assign n21681 = ~n21704;
  assign n21691 = n21648 & n18532;
  assign n21690 = ~n21648;
  assign n21715 = n21716 & n21726;
  assign n21658 = n21727 & n21728;
  assign n21693 = ~n21741;
  assign n21697 = n21757 & n21758;
  assign n21729 = ~n21759;
  assign n21742 = n21770 ^ n21771;
  assign n21760 = ~n21770;
  assign n21772 = n21792 ^ n18055;
  assign n21794 = n21743 & n21803;
  assign n21793 = ~n21743;
  assign n21804 = ~n21817;
  assign n21621 = ~n21656;
  assign n21500 = n21681 & n21682;
  assign n21683 = n21690 & n18525;
  assign n21624 = ~n21691;
  assign n21692 = ~n21715;
  assign n21661 = ~n21658;
  assign n21706 = n21693 & n21716;
  assign n21717 = n21742 ^ n21743;
  assign n21731 = n21729 & n21695;
  assign n21730 = ~n21697;
  assign n21762 = n21772 & n21773;
  assign n21763 = ~n21772;
  assign n21785 = n21793 & n21771;
  assign n21733 = ~n21794;
  assign n21774 = n21804 & n21805;
  assign n21616 = n21620 & n21621;
  assign n21622 = n21621 & n21599;
  assign n21549 = ~n21500;
  assign n21657 = ~n21683;
  assign n21684 = n21692 & n21693;
  assign n21673 = ~n21706;
  assign n21707 = n21717 & n72;
  assign n21718 = n21729 & n21730;
  assign n21705 = ~n21717;
  assign n21698 = ~n21731;
  assign n21667 = ~n21762;
  assign n21751 = n21763 & n21764;
  assign n21745 = n21774 ^ n19260;
  assign n21761 = ~n21785;
  assign n21775 = ~n21774;
  assign n21598 = ~n21616;
  assign n21597 = ~n21622;
  assign n17459 = n21672 ^ n21673;
  assign n21647 = ~n21684;
  assign n21659 = n21697 ^ n21698;
  assign n21696 = n21705 & n2975;
  assign n21630 = ~n21707;
  assign n21694 = ~n21718;
  assign n18026 = n21744 ^ n21745;
  assign n21700 = ~n21751;
  assign n21750 = n21760 & n21761;
  assign n21765 = n21775 & n21776;
  assign n19617 = n21596 ^ n21597;
  assign n21560 = n21598 & n21599;
  assign n21617 = n21647 ^ n21648;
  assign n21646 = n21647 & n21657;
  assign n21637 = n21658 ^ n21659;
  assign n17562 = ~n17459;
  assign n21660 = ~n21659;
  assign n21627 = n21694 & n21695;
  assign n21662 = ~n21696;
  assign n21632 = n21708 ^ n18026;
  assign n21719 = n21700 & n21667;
  assign n18031 = ~n18026;
  assign n21732 = ~n21750;
  assign n21746 = ~n21765;
  assign n21463 = n4 ^ n21560;
  assign n19646 = ~n19617;
  assign n21427 = ~n21560;
  assign n17375 = n21617 ^ n18532;
  assign n21626 = n21637 & n18454;
  assign n21610 = n17562 & n19768;
  assign n21623 = ~n21646;
  assign n21625 = ~n21637;
  assign n21602 = n21660 & n21661;
  assign n21664 = n21662 & n21630;
  assign n21663 = ~n21627;
  assign n21675 = n21632 & n21685;
  assign n21674 = ~n21632;
  assign n21687 = ~n21719;
  assign n21686 = n21732 & n21733;
  assign n21709 = n21746 & n21747;
  assign n17462 = ~n17375;
  assign n21590 = n21610 ^ n18582;
  assign n21555 = n21623 & n21624;
  assign n21618 = n21625 & n18491;
  assign n21600 = ~n21626;
  assign n21611 = ~n21602;
  assign n21649 = n21662 & n21663;
  assign n21628 = ~n21664;
  assign n21668 = n21674 & n21607;
  assign n21634 = ~n21675;
  assign n21665 = n21686 ^ n21687;
  assign n17975 = n21709 ^ n21710;
  assign n21699 = ~n21686;
  assign n21711 = ~n21709;
  assign n21554 = n17462 & n19744;
  assign n21578 = n21590 & n21591;
  assign n21576 = ~n21590;
  assign n21601 = ~n21555;
  assign n21562 = ~n21618;
  assign n21603 = n21627 ^ n21628;
  assign n21629 = ~n21649;
  assign n21651 = n21665 & n87;
  assign n21609 = ~n21668;
  assign n21650 = ~n21665;
  assign n21543 = n21676 ^ n17975;
  assign n21688 = n21699 & n21700;
  assign n17944 = ~n17975;
  assign n21701 = n21711 & n21712;
  assign n21440 = n21554 ^ n18525;
  assign n21565 = n21576 & n21577;
  assign n21518 = ~n21578;
  assign n21589 = n21600 & n21601;
  assign n21592 = n21562 & n21600;
  assign n21536 = n21602 ^ n21603;
  assign n21550 = n21603 & n21611;
  assign n21580 = n21629 & n21630;
  assign n21638 = n21650 & n2910;
  assign n21567 = ~n21651;
  assign n21639 = n21543 & n21571;
  assign n21640 = ~n21543;
  assign n21666 = ~n21688;
  assign n21677 = ~n21701;
  assign n21528 = n21440 & n21533;
  assign n21529 = ~n21440;
  assign n21548 = ~n21565;
  assign n21563 = n21536 & n18464;
  assign n21561 = ~n21589;
  assign n21556 = ~n21592;
  assign n21564 = ~n21536;
  assign n21604 = ~n21580;
  assign n21605 = ~n21638;
  assign n21545 = ~n21639;
  assign n21635 = n21640 & n21641;
  assign n21631 = n21666 & n21667;
  assign n21642 = n21677 & n21678;
  assign n21442 = ~n21528;
  assign n21519 = n21529 & n21486;
  assign n21534 = n21548 & n21549;
  assign n21539 = n21518 & n21548;
  assign n17295 = n21555 ^ n21556;
  assign n21535 = n21561 & n21562;
  assign n21538 = ~n21563;
  assign n21557 = n21564 & n18474;
  assign n21593 = n21604 & n21605;
  assign n21612 = n21605 & n21567;
  assign n21606 = n21631 ^ n21632;
  assign n21573 = ~n21635;
  assign n17885 = n21642 ^ n21643;
  assign n21633 = ~n21631;
  assign n21644 = ~n21642;
  assign n21487 = ~n21519;
  assign n21517 = ~n21534;
  assign n21499 = n21535 ^ n21536;
  assign n21501 = ~n21539;
  assign n17405 = ~n17295;
  assign n21537 = ~n21535;
  assign n21503 = ~n21557;
  assign n21566 = ~n21593;
  assign n21579 = n21606 ^ n21607;
  assign n21581 = ~n21612;
  assign n21594 = n21613 ^ n17885;
  assign n21619 = n21633 & n21634;
  assign n17939 = ~n17885;
  assign n21636 = n21644 & n21645;
  assign n17216 = n18474 ^ n21499;
  assign n21464 = n21500 ^ n21501;
  assign n21485 = n21517 & n21518;
  assign n21493 = n17405 & n19703;
  assign n21530 = n21537 & n21538;
  assign n21494 = n21566 & n21567;
  assign n21569 = n21579 & n86;
  assign n21551 = n21580 ^ n21581;
  assign n21568 = ~n21579;
  assign n21584 = n21594 & n21595;
  assign n21582 = ~n21594;
  assign n21608 = ~n21619;
  assign n21614 = ~n21636;
  assign n21423 = n21463 ^ n21464;
  assign n21465 = n17216 & n21484;
  assign n21439 = n21485 ^ n21486;
  assign n21469 = n21464 & n4;
  assign n17280 = ~n17216;
  assign n21470 = n21493 ^ n18454;
  assign n21467 = ~n21464;
  assign n21488 = ~n21485;
  assign n21502 = ~n21530;
  assign n21473 = n21550 ^ n21551;
  assign n21456 = n21551 & n21550;
  assign n21540 = ~n21494;
  assign n21558 = n21568 & n2896;
  assign n21506 = ~n21569;
  assign n21574 = n21582 & n21583;
  assign n21483 = ~n21584;
  assign n21570 = n21608 & n21609;
  assign n21586 = n21614 & n21615;
  assign n19609 = n21423 ^ n19617;
  assign n21312 = n21439 ^ n21440;
  assign n21424 = ~n21423;
  assign n21425 = n17280 & n19663;
  assign n21450 = n17280 & n19725;
  assign n19708 = ~n21465;
  assign n21451 = n21467 & n21468;
  assign n21392 = ~n21469;
  assign n21454 = n21470 & n21471;
  assign n21466 = n21487 & n21488;
  assign n21452 = ~n21470;
  assign n21472 = n21502 & n21503;
  assign n21520 = n21473 & n18406;
  assign n21521 = ~n21473;
  assign n21541 = ~n21558;
  assign n21542 = n21570 ^ n21571;
  assign n21512 = ~n21574;
  assign n17862 = n21585 ^ n21586;
  assign n21572 = ~n21570;
  assign n21587 = ~n21586;
  assign n21240 = ~n19609;
  assign n21408 = n21312 & n3;
  assign n21275 = n21424 & n19617;
  assign n21406 = ~n21312;
  assign n21281 = n21425 ^ n18464;
  assign n19727 = ~n21450;
  assign n21426 = ~n21451;
  assign n21443 = n21452 & n21453;
  assign n21369 = ~n21454;
  assign n21441 = ~n21466;
  assign n21428 = n21472 ^ n21473;
  assign n21474 = ~n21472;
  assign n21430 = ~n21520;
  assign n21504 = n21521 & n18398;
  assign n21531 = n21540 & n21541;
  assign n21532 = n21541 & n21506;
  assign n21477 = n21542 ^ n21543;
  assign n21546 = n21512 & n21483;
  assign n21559 = n21572 & n21573;
  assign n17864 = ~n17862;
  assign n21575 = n21587 & n21588;
  assign n21387 = n21406 & n21407;
  assign n21388 = n21281 & n21318;
  assign n21314 = ~n21408;
  assign n21389 = ~n21281;
  assign n21417 = n21426 & n21427;
  assign n17131 = n18406 ^ n21428;
  assign n21381 = n21441 & n21442;
  assign n21410 = ~n21443;
  assign n21475 = ~n21504;
  assign n21507 = n21477 & n2826;
  assign n21505 = ~n21531;
  assign n21495 = ~n21532;
  assign n21508 = ~n21477;
  assign n21510 = ~n21546;
  assign n21522 = n21547 ^ n17864;
  assign n21544 = ~n21559;
  assign n21552 = ~n21575;
  assign n21350 = ~n21387;
  assign n21295 = ~n21388;
  assign n21378 = n21389 & n21390;
  assign n21367 = n17131 & n19645;
  assign n21394 = n17131 & n21409;
  assign n21391 = ~n21417;
  assign n17175 = ~n17131;
  assign n21380 = n21369 & n21410;
  assign n21411 = ~n21381;
  assign n21455 = n21474 & n21475;
  assign n21457 = n21494 ^ n21495;
  assign n21476 = n21505 & n21506;
  assign n21479 = ~n21507;
  assign n21496 = n21508 & n85;
  assign n21513 = n21522 & n21523;
  assign n21514 = ~n21522;
  assign n21509 = n21544 & n21545;
  assign n21524 = n21552 & n21553;
  assign n21258 = n21367 ^ n18406;
  assign n21333 = ~n21378;
  assign n21233 = n21380 ^ n21381;
  assign n21352 = n21391 & n21392;
  assign n21379 = n17175 & n21393;
  assign n19690 = ~n21394;
  assign n21395 = n21410 & n21411;
  assign n21429 = ~n21455;
  assign n21431 = n21456 ^ n21457;
  assign n21396 = n21457 & n21456;
  assign n21432 = n21476 ^ n21477;
  assign n21478 = ~n21476;
  assign n21434 = ~n21496;
  assign n21489 = n21509 ^ n21510;
  assign n21405 = ~n21513;
  assign n21498 = n21514 & n21515;
  assign n17772 = n21524 ^ n21525;
  assign n21511 = ~n21509;
  assign n21526 = ~n21524;
  assign n21331 = n21258 & n21341;
  assign n21311 = n3 ^ n21352;
  assign n21332 = ~n21258;
  assign n21343 = n21233 & n21353;
  assign n21345 = ~n21233;
  assign n21351 = ~n21352;
  assign n19673 = ~n21379;
  assign n21368 = ~n21395;
  assign n21335 = n21429 & n21430;
  assign n21418 = n21431 & n18363;
  assign n21397 = n85 ^ n21432;
  assign n21419 = ~n21431;
  assign n21399 = ~n21396;
  assign n21458 = n21478 & n21479;
  assign n21481 = n21489 & n84;
  assign n21460 = n21490 ^ n17772;
  assign n21480 = ~n21489;
  assign n21436 = ~n21498;
  assign n21497 = n21511 & n21512;
  assign n17877 = ~n17772;
  assign n21516 = n21526 & n21527;
  assign n21276 = n21311 ^ n21312;
  assign n21260 = ~n21331;
  assign n21315 = n21332 & n21210;
  assign n21279 = ~n21343;
  assign n21334 = n21345 & n2;
  assign n21342 = n21350 & n21351;
  assign n21344 = n19673 & n19690;
  assign n21354 = n21368 & n21369;
  assign n21370 = n21396 ^ n21397;
  assign n21382 = ~n21335;
  assign n21347 = ~n21418;
  assign n21412 = n21419 & n18361;
  assign n21398 = ~n21397;
  assign n21433 = ~n21458;
  assign n21444 = n21460 & n21461;
  assign n21459 = n21480 & n2783;
  assign n21360 = ~n21481;
  assign n21462 = n21436 & n21405;
  assign n21445 = ~n21460;
  assign n21482 = ~n21497;
  assign n21491 = ~n21516;
  assign n19576 = n21275 ^ n21276;
  assign n21277 = ~n21276;
  assign n21212 = ~n21315;
  assign n21235 = ~n21334;
  assign n21313 = ~n21342;
  assign n19688 = ~n21344;
  assign n21317 = ~n21354;
  assign n21356 = n21370 & n18319;
  assign n21355 = ~n21370;
  assign n21357 = n21398 & n21399;
  assign n21383 = ~n21412;
  assign n21401 = n21433 & n21434;
  assign n21328 = ~n21444;
  assign n21437 = n21445 & n21446;
  assign n21403 = ~n21459;
  assign n21421 = ~n21462;
  assign n21420 = n21482 & n21483;
  assign n21447 = n21491 & n21492;
  assign n21151 = ~n19576;
  assign n21191 = n21277 & n21275;
  assign n21278 = n21313 & n21314;
  assign n21282 = n21317 ^ n21318;
  assign n21316 = n21333 & n21317;
  assign n21348 = n21355 & n18322;
  assign n21304 = ~n21356;
  assign n21371 = n21382 & n21383;
  assign n21372 = n21383 & n21347;
  assign n21402 = ~n21401;
  assign n21322 = n21420 ^ n21421;
  assign n21400 = n21403 & n21360;
  assign n21364 = ~n21437;
  assign n21413 = n21447 ^ n19036;
  assign n21435 = ~n21420;
  assign n21448 = ~n21447;
  assign n21232 = n2 ^ n21278;
  assign n21256 = n21281 ^ n21282;
  assign n21280 = ~n21278;
  assign n21294 = ~n21316;
  assign n21271 = ~n21348;
  assign n21346 = ~n21371;
  assign n21336 = ~n21372;
  assign n21358 = n21400 ^ n21401;
  assign n21384 = n21402 & n21403;
  assign n21386 = n21322 & n83;
  assign n21385 = ~n21322;
  assign n21361 = n21364 & n21328;
  assign n17750 = n21413 ^ n21414;
  assign n21422 = n21435 & n21436;
  assign n21438 = n21448 & n21449;
  assign n21192 = n21232 ^ n21233;
  assign n21238 = n21256 & n1;
  assign n21236 = ~n21256;
  assign n21269 = n21279 & n21280;
  assign n21257 = n21294 & n21295;
  assign n21283 = n21304 & n21271;
  assign n17147 = n21335 ^ n21336;
  assign n21284 = n21346 & n21347;
  assign n21183 = n21357 ^ n21358;
  assign n21242 = n21358 & n21357;
  assign n21359 = ~n21384;
  assign n21373 = n21385 & n2766;
  assign n21287 = ~n21386;
  assign n17835 = ~n17750;
  assign n21404 = ~n21422;
  assign n21415 = ~n21438;
  assign n21072 = n21191 ^ n21192;
  assign n21097 = n21192 & n21191;
  assign n21224 = n21236 & n21237;
  assign n21150 = ~n21238;
  assign n21209 = n21257 ^ n21258;
  assign n21234 = ~n21269;
  assign n21259 = ~n21257;
  assign n17121 = n21283 ^ n21284;
  assign n17096 = ~n17147;
  assign n21320 = n21183 & n18264;
  assign n21305 = ~n21284;
  assign n21319 = ~n21183;
  assign n21245 = ~n21242;
  assign n21321 = n21359 & n21360;
  assign n21251 = n21365 ^ n17835;
  assign n21324 = ~n21373;
  assign n21362 = n21404 & n21405;
  assign n21374 = n21415 & n21416;
  assign n21087 = ~n21072;
  assign n21101 = ~n21097;
  assign n21069 = n21209 ^ n21210;
  assign n21193 = ~n21224;
  assign n21141 = n21234 & n21235;
  assign n21239 = n17121 & n19609;
  assign n21241 = n21259 & n21260;
  assign n21213 = n17121 & n19529;
  assign n17025 = ~n17121;
  assign n21261 = n17096 & n19550;
  assign n21296 = n21304 & n21305;
  assign n21306 = n21319 & n18233;
  assign n21229 = ~n21320;
  assign n21285 = n21321 ^ n21322;
  assign n21330 = n21251 & n21337;
  assign n21323 = ~n21321;
  assign n21329 = ~n21251;
  assign n21247 = n21361 ^ n21362;
  assign n21338 = n21374 ^ n21375;
  assign n21363 = ~n21362;
  assign n21376 = ~n21374;
  assign n21169 = n21069 & n0;
  assign n21167 = ~n21069;
  assign n21182 = n21193 & n21150;
  assign n21045 = n21213 ^ n18319;
  assign n21194 = ~n21141;
  assign n19611 = ~n21239;
  assign n21225 = n17025 & n21240;
  assign n21211 = ~n21241;
  assign n21127 = n21261 ^ n18361;
  assign n21243 = n83 ^ n21285;
  assign n21270 = ~n21296;
  assign n21186 = ~n21306;
  assign n21307 = n21323 & n21324;
  assign n21309 = n21329 & n21289;
  assign n21253 = ~n21330;
  assign n21325 = n21247 & n2673;
  assign n17784 = n18920 ^ n21338;
  assign n21326 = ~n21247;
  assign n21349 = n21363 & n21364;
  assign n21366 = n21376 & n21377;
  assign n21148 = n21167 & n21168;
  assign n21071 = ~n21169;
  assign n21142 = ~n21182;
  assign n21174 = n21045 & n21089;
  assign n21181 = n21193 & n21194;
  assign n21175 = ~n21045;
  assign n21170 = n21211 & n21212;
  assign n19594 = ~n21225;
  assign n21215 = n21127 & n21226;
  assign n21214 = n21242 ^ n21243;
  assign n21216 = ~n21127;
  assign n21227 = n21270 & n21271;
  assign n21244 = ~n21243;
  assign n21163 = n21297 ^ n17784;
  assign n20325 = n21298 ^ n17784;
  assign n21286 = ~n21307;
  assign n21290 = ~n21309;
  assign n21299 = n17784 & n21310;
  assign n21249 = ~n21325;
  assign n21308 = n21326 & n82;
  assign n17776 = ~n17784;
  assign n21327 = ~n21349;
  assign n21339 = ~n21366;
  assign n21098 = n21141 ^ n21142;
  assign n21109 = ~n21148;
  assign n21128 = n21170 ^ n21171;
  assign n21048 = ~n21174;
  assign n21153 = n21175 & n21176;
  assign n21149 = ~n21181;
  assign n21172 = ~n21170;
  assign n21196 = n21214 & n18252;
  assign n21130 = ~n21215;
  assign n21197 = n21216 & n21171;
  assign n21184 = n21227 ^ n18233;
  assign n21195 = ~n21214;
  assign n21154 = n21244 & n21245;
  assign n21228 = ~n21227;
  assign n21263 = n21163 & n21272;
  assign n21246 = n21286 & n21287;
  assign n21262 = ~n21163;
  assign n21292 = n17776 & n21298;
  assign n20306 = ~n21299;
  assign n21200 = ~n21308;
  assign n21288 = n21327 & n21328;
  assign n21300 = n21339 & n21340;
  assign n19476 = n21097 ^ n21098;
  assign n21002 = n21127 ^ n21128;
  assign n21100 = ~n21098;
  assign n21111 = n21149 & n21150;
  assign n21091 = ~n21153;
  assign n16979 = n21183 ^ n21184;
  assign n21187 = n21195 & n18248;
  assign n21104 = ~n21196;
  assign n21173 = ~n21197;
  assign n21217 = n21228 & n21229;
  assign n21157 = ~n21154;
  assign n21198 = n21246 ^ n21247;
  assign n21254 = n21262 & n21204;
  assign n21165 = ~n21263;
  assign n21248 = ~n21246;
  assign n21250 = n21288 ^ n21289;
  assign n20327 = ~n21292;
  assign n17733 = n21300 ^ n21301;
  assign n21291 = ~n21288;
  assign n21302 = ~n21300;
  assign n20989 = ~n19476;
  assign n21024 = n21100 & n21101;
  assign n21068 = n0 ^ n21111;
  assign n21110 = ~n21111;
  assign n21143 = n16979 & n21151;
  assign n21152 = n21172 & n21173;
  assign n17012 = ~n16979;
  assign n21145 = ~n21187;
  assign n21155 = n82 ^ n21198;
  assign n21185 = ~n21217;
  assign n21230 = n21248 & n21249;
  assign n21159 = n21250 ^ n21251;
  assign n21206 = ~n21254;
  assign n21122 = n21264 ^ n17733;
  assign n21265 = n17733 & n21274;
  assign n21273 = n21290 & n21291;
  assign n17641 = ~n17733;
  assign n21293 = n21302 & n21303;
  assign n21025 = n21068 ^ n21069;
  assign n21027 = ~n21024;
  assign n21099 = n21109 & n21110;
  assign n19557 = ~n21143;
  assign n21131 = n17012 & n19576;
  assign n21102 = n17012 & n19452;
  assign n21129 = ~n21152;
  assign n21112 = n21145 & n21104;
  assign n21132 = n21154 ^ n21155;
  assign n21113 = n21185 & n21186;
  assign n21156 = ~n21155;
  assign n21202 = n21159 & n81;
  assign n21199 = ~n21230;
  assign n21201 = ~n21159;
  assign n21219 = n21122 & n21231;
  assign n21218 = ~n21122;
  assign n20264 = ~n21265;
  assign n21255 = n17641 & n21266;
  assign n21252 = ~n21273;
  assign n21267 = ~n21293;
  assign n20903 = n21024 ^ n21025;
  assign n21026 = ~n21025;
  assign n21070 = ~n21099;
  assign n20968 = n21102 ^ n18264;
  assign n16948 = n21112 ^ n21113;
  assign n21088 = n21129 & n21130;
  assign n19578 = ~n21131;
  assign n21114 = n21132 & n18201;
  assign n21115 = ~n21132;
  assign n21076 = n21156 & n21157;
  assign n21144 = ~n21113;
  assign n21158 = n21199 & n21200;
  assign n21188 = n21201 & n2621;
  assign n21118 = ~n21202;
  assign n21207 = n21218 & n21083;
  assign n21124 = ~n21219;
  assign n21203 = n21252 & n21253;
  assign n20286 = ~n21255;
  assign n21220 = n21267 & n21268;
  assign n20894 = ~n20903;
  assign n20949 = n21026 & n21027;
  assign n21043 = n21070 & n21071;
  assign n21062 = n20968 & n21074;
  assign n21073 = n16948 & n21087;
  assign n21046 = n21088 ^ n21089;
  assign n21063 = ~n20968;
  assign n21050 = n16948 & n19494;
  assign n16950 = ~n16948;
  assign n21090 = ~n21088;
  assign n21064 = ~n21114;
  assign n21105 = n21115 & n18174;
  assign n21133 = n21144 & n21145;
  assign n21079 = ~n21076;
  assign n21116 = n21158 ^ n21159;
  assign n21160 = ~n21158;
  assign n21161 = ~n21188;
  assign n21162 = n21203 ^ n21204;
  assign n21085 = ~n21207;
  assign n20283 = n20286 & n20264;
  assign n17517 = n21220 ^ n21221;
  assign n21205 = ~n21203;
  assign n21222 = ~n21220;
  assign n21028 = n21043 & n21044;
  assign n20876 = n21045 ^ n21046;
  assign n20924 = n21050 ^ n18252;
  assign n21013 = ~n21043;
  assign n20970 = ~n21062;
  assign n21049 = n21063 & n21004;
  assign n21061 = n16950 & n21072;
  assign n19545 = ~n21073;
  assign n21075 = n21090 & n21091;
  assign n21017 = ~n21105;
  assign n21077 = n81 ^ n21116;
  assign n21103 = ~n21133;
  assign n21146 = n21160 & n21161;
  assign n21134 = n21162 ^ n21163;
  assign n21038 = n21177 ^ n17517;
  assign n21178 = n17517 & n21190;
  assign n21189 = n21205 & n21206;
  assign n17588 = ~n17517;
  assign n21208 = n21222 & n21223;
  assign n20978 = n21013 ^ n21002;
  assign n21008 = n20924 & n21015;
  assign n21014 = n21013 & n15;
  assign n21001 = ~n21028;
  assign n20892 = ~n20876;
  assign n21007 = ~n20924;
  assign n21006 = ~n21049;
  assign n19522 = ~n21061;
  assign n21047 = ~n21075;
  assign n21029 = n21017 & n21064;
  assign n21051 = n21076 ^ n21077;
  assign n21030 = n21103 & n21104;
  assign n21078 = ~n21077;
  assign n21120 = n21134 & n80;
  assign n21117 = ~n21146;
  assign n21119 = ~n21134;
  assign n21135 = n21038 & n21147;
  assign n21136 = ~n21038;
  assign n20227 = ~n21178;
  assign n21166 = n17588 & n20225;
  assign n21164 = ~n21189;
  assign n21179 = ~n21208;
  assign n20950 = n15 ^ n20978;
  assign n20988 = n21001 & n21002;
  assign n20992 = n21007 & n20878;
  assign n20926 = ~n21008;
  assign n20966 = ~n21014;
  assign n19542 = n19545 & n19522;
  assign n16963 = n21029 ^ n21030;
  assign n21003 = n21047 & n21048;
  assign n21032 = n21051 & n18186;
  assign n21031 = ~n21051;
  assign n20983 = n21078 & n21079;
  assign n21065 = ~n21030;
  assign n21019 = n21117 & n21118;
  assign n21106 = n21119 & n2593;
  assign n21034 = ~n21120;
  assign n21040 = ~n21135;
  assign n21125 = n21136 & n20996;
  assign n21121 = n21164 & n21165;
  assign n20242 = ~n21166;
  assign n21138 = n21179 & n21180;
  assign n19403 = n20949 ^ n20950;
  assign n20837 = n20950 & n20949;
  assign n20965 = ~n20988;
  assign n20881 = ~n20992;
  assign n20990 = n16963 & n19476;
  assign n20967 = n21003 ^ n21004;
  assign n20971 = n16963 & n19434;
  assign n16969 = ~n16963;
  assign n21005 = ~n21003;
  assign n21018 = n21031 & n18179;
  assign n20942 = ~n21032;
  assign n21052 = n21064 & n21065;
  assign n20986 = ~n20983;
  assign n21080 = ~n21019;
  assign n21081 = ~n21106;
  assign n21082 = n21121 ^ n21122;
  assign n20998 = ~n21125;
  assign n17574 = n21137 ^ n21138;
  assign n21123 = ~n21121;
  assign n21139 = ~n21138;
  assign n20820 = ~n19403;
  assign n20840 = ~n20837;
  assign n20917 = n20965 & n20966;
  assign n20936 = n20967 ^ n20968;
  assign n20937 = n20971 ^ n18201;
  assign n20979 = n16969 & n20989;
  assign n19506 = ~n20990;
  assign n20991 = n21005 & n21006;
  assign n20981 = ~n21018;
  assign n21016 = ~n21052;
  assign n21066 = n21080 & n21081;
  assign n21067 = n21081 & n21034;
  assign n21053 = n21082 ^ n21083;
  assign n20958 = n21092 ^ n17574;
  assign n21094 = n17574 & n21108;
  assign n21107 = n21123 & n21124;
  assign n17586 = ~n17574;
  assign n21126 = n21139 & n21140;
  assign n20875 = n14 ^ n20917;
  assign n20921 = n20917 & n20935;
  assign n20922 = n20936 & n13;
  assign n20929 = n20937 & n20938;
  assign n20918 = ~n20917;
  assign n20919 = ~n20936;
  assign n20927 = ~n20937;
  assign n19479 = ~n20979;
  assign n20969 = ~n20991;
  assign n20982 = n20981 & n20942;
  assign n20939 = n21016 & n21017;
  assign n21036 = n21053 & n95;
  assign n21033 = ~n21066;
  assign n21020 = ~n21067;
  assign n21035 = ~n21053;
  assign n21056 = n20958 & n20913;
  assign n21054 = ~n20958;
  assign n21086 = n17586 & n21093;
  assign n20208 = ~n21094;
  assign n21084 = ~n21107;
  assign n21095 = ~n21126;
  assign n20838 = n20875 ^ n20876;
  assign n20901 = n20918 & n14;
  assign n20902 = n20919 & n20920;
  assign n20891 = ~n20921;
  assign n20761 = ~n20922;
  assign n20905 = n20927 & n20928;
  assign n20805 = ~n20929;
  assign n20923 = n20969 & n20970;
  assign n20940 = ~n20982;
  assign n20980 = ~n20939;
  assign n20984 = n21019 ^ n21020;
  assign n20952 = n21033 & n21034;
  assign n21021 = n21035 & n2483;
  assign n20954 = ~n21036;
  assign n21041 = n21054 & n21055;
  assign n20915 = ~n21056;
  assign n21037 = n21084 & n21085;
  assign n20185 = ~n21086;
  assign n21057 = n21095 & n21096;
  assign n20747 = n20837 ^ n20838;
  assign n20839 = ~n20838;
  assign n20874 = n20891 & n20892;
  assign n20849 = ~n20901;
  assign n20809 = ~n20902;
  assign n20841 = ~n20905;
  assign n20877 = n20923 ^ n20924;
  assign n16928 = n20939 ^ n20940;
  assign n20925 = ~n20923;
  assign n20972 = n20980 & n20981;
  assign n20896 = n20983 ^ n20984;
  assign n20985 = ~n20984;
  assign n20993 = ~n20952;
  assign n20994 = ~n21021;
  assign n20995 = n21037 ^ n21038;
  assign n20960 = ~n21041;
  assign n20205 = n20208 & n20185;
  assign n17543 = n21057 ^ n21058;
  assign n21039 = ~n21037;
  assign n21059 = ~n21057;
  assign n20726 = ~n20747;
  assign n20758 = n20839 & n20840;
  assign n20848 = ~n20874;
  assign n20860 = n20809 & n20761;
  assign n20859 = n20877 ^ n20878;
  assign n20861 = n20805 & n20841;
  assign n20893 = n16928 & n20903;
  assign n20904 = n20925 & n20926;
  assign n16917 = ~n16928;
  assign n20944 = n20896 & n18151;
  assign n20941 = ~n20972;
  assign n20943 = ~n20896;
  assign n20906 = n20985 & n20986;
  assign n20987 = n20993 & n20994;
  assign n20951 = n20994 & n20954;
  assign n20973 = n20995 ^ n20996;
  assign n21009 = n17543 & n21023;
  assign n21022 = n21039 & n21040;
  assign n17533 = ~n17543;
  assign n21042 = n21059 & n21060;
  assign n20772 = ~n20758;
  assign n20806 = n20848 & n20849;
  assign n20847 = n20859 & n12;
  assign n20807 = ~n20860;
  assign n20835 = ~n20859;
  assign n20822 = ~n20861;
  assign n19444 = ~n20893;
  assign n20879 = n16917 & n20894;
  assign n20851 = n16917 & n19339;
  assign n20880 = ~n20904;
  assign n20895 = n20941 & n20942;
  assign n20930 = n20943 & n18077;
  assign n20898 = ~n20944;
  assign n20907 = n20951 ^ n20952;
  assign n20909 = ~n20906;
  assign n20956 = n20973 & n94;
  assign n20953 = ~n20987;
  assign n20955 = ~n20973;
  assign n20830 = n17533 ^ n20999;
  assign n20141 = ~n21009;
  assign n21000 = n17533 & n21010;
  assign n20997 = ~n21022;
  assign n21011 = ~n21042;
  assign n20759 = n20806 ^ n20807;
  assign n20819 = n20835 & n20836;
  assign n20808 = ~n20806;
  assign n20674 = ~n20847;
  assign n20824 = n20851 ^ n18179;
  assign n19464 = ~n20879;
  assign n20821 = n20880 & n20881;
  assign n20850 = n20895 ^ n20896;
  assign n20883 = n20906 ^ n20907;
  assign n20897 = ~n20895;
  assign n20853 = ~n20930;
  assign n20908 = ~n20907;
  assign n20855 = n20953 & n20954;
  assign n20945 = n20955 & n2398;
  assign n20865 = ~n20956;
  assign n20963 = n20830 & n20869;
  assign n20961 = ~n20830;
  assign n20957 = n20997 & n20998;
  assign n20164 = ~n21000;
  assign n20974 = n21011 & n21012;
  assign n19349 = n20758 ^ n20759;
  assign n20670 = n20759 & n20772;
  assign n20794 = n20808 & n20809;
  assign n20714 = ~n20819;
  assign n20796 = n20821 ^ n20822;
  assign n20813 = n20824 & n20825;
  assign n20811 = ~n20824;
  assign n19461 = n19464 & n19444;
  assign n16837 = n20850 ^ n18151;
  assign n20842 = ~n20821;
  assign n20863 = n20883 & n18112;
  assign n20882 = n20897 & n20898;
  assign n20862 = ~n20883;
  assign n20816 = n20908 & n20909;
  assign n20910 = ~n20855;
  assign n20911 = ~n20945;
  assign n20912 = n20957 ^ n20958;
  assign n20947 = n20961 & n20962;
  assign n20871 = ~n20963;
  assign n20161 = n20164 & n20141;
  assign n17272 = n20974 ^ n20975;
  assign n20959 = ~n20957;
  assign n20976 = ~n20974;
  assign n20642 = ~n19349;
  assign n20760 = ~n20794;
  assign n20773 = n20714 & n20674;
  assign n20776 = n20796 & n11;
  assign n20774 = ~n20796;
  assign n20797 = n20811 & n20812;
  assign n20701 = ~n20813;
  assign n20810 = n16837 & n20820;
  assign n20793 = n16837 & n19354;
  assign n20823 = n20841 & n20842;
  assign n16907 = ~n16837;
  assign n20854 = n20862 & n18106;
  assign n20763 = ~n20863;
  assign n20852 = ~n20882;
  assign n20899 = n20910 & n20911;
  assign n20900 = n20911 & n20865;
  assign n20781 = n20912 ^ n20913;
  assign n20740 = n20931 ^ n17272;
  assign n20832 = ~n20947;
  assign n20932 = n17272 & n20948;
  assign n20946 = n20959 & n20960;
  assign n17435 = ~n17272;
  assign n20964 = n20976 & n20977;
  assign n20711 = n20760 & n20761;
  assign n20712 = ~n20773;
  assign n20757 = n20774 & n20775;
  assign n20605 = ~n20776;
  assign n20748 = n20793 ^ n18151;
  assign n20746 = ~n20797;
  assign n20795 = n16907 & n19403;
  assign n19423 = ~n20810;
  assign n20804 = ~n20823;
  assign n20778 = n20852 & n20853;
  assign n20815 = ~n20854;
  assign n20866 = n20781 & n2323;
  assign n20864 = ~n20899;
  assign n20856 = ~n20900;
  assign n20867 = ~n20781;
  assign n20886 = n20740 & n20787;
  assign n20884 = ~n20740;
  assign n20104 = ~n20932;
  assign n20916 = n17435 & n20102;
  assign n20914 = ~n20946;
  assign n20933 = ~n20964;
  assign n20671 = n20711 ^ n20712;
  assign n20713 = ~n20711;
  assign n20728 = n20748 & n20749;
  assign n20641 = ~n20757;
  assign n20717 = n20701 & n20746;
  assign n20729 = ~n20748;
  assign n19406 = ~n20795;
  assign n20718 = n20804 & n20805;
  assign n20777 = n20815 & n20763;
  assign n20814 = ~n20778;
  assign n20817 = n20855 ^ n20856;
  assign n20826 = n20864 & n20865;
  assign n20827 = ~n20866;
  assign n20857 = n20867 & n93;
  assign n20872 = n20884 & n20885;
  assign n20742 = ~n20886;
  assign n20868 = n20914 & n20915;
  assign n20120 = ~n20916;
  assign n20888 = n20933 & n20934;
  assign n20586 = n20670 ^ n20671;
  assign n20602 = n20671 & n20670;
  assign n20699 = n20713 & n20714;
  assign n20573 = n20717 ^ n20718;
  assign n20715 = n20641 & n20605;
  assign n20633 = ~n20728;
  assign n20716 = n20729 & n20730;
  assign n16796 = n20777 ^ n20778;
  assign n20745 = ~n20718;
  assign n20798 = n20814 & n20815;
  assign n20779 = n20816 ^ n20817;
  assign n20731 = n20817 & n20816;
  assign n20780 = n93 ^ n20826;
  assign n20828 = ~n20826;
  assign n20783 = ~n20857;
  assign n20829 = n20868 ^ n20869;
  assign n20789 = ~n20872;
  assign n17236 = n20887 ^ n20888;
  assign n20870 = ~n20868;
  assign n20889 = ~n20888;
  assign n20577 = ~n20586;
  assign n20675 = n20573 & n20683;
  assign n20673 = ~n20699;
  assign n20677 = ~n20573;
  assign n20639 = ~n20715;
  assign n20659 = ~n20716;
  assign n20725 = n20745 & n20746;
  assign n20727 = n16796 & n20747;
  assign n20698 = n16796 & n19331;
  assign n16874 = ~n16796;
  assign n20764 = n20779 & n18055;
  assign n20732 = n20780 ^ n20781;
  assign n20762 = ~n20798;
  assign n20765 = ~n20779;
  assign n20734 = ~n20731;
  assign n20818 = n20827 & n20828;
  assign n20736 = n20829 ^ n20830;
  assign n20843 = n17236 & n20062;
  assign n20858 = n20870 & n20871;
  assign n17389 = ~n17236;
  assign n20873 = n20889 & n20890;
  assign n20638 = n20673 & n20674;
  assign n20575 = ~n20675;
  assign n20661 = n20677 & n10;
  assign n20676 = n20633 & n20659;
  assign n20596 = n20698 ^ n18106;
  assign n20700 = ~n20725;
  assign n20710 = n16874 & n20726;
  assign n19391 = ~n20727;
  assign n20702 = n20731 ^ n20732;
  assign n20666 = n20762 & n20763;
  assign n20679 = ~n20764;
  assign n20750 = n20765 & n18021;
  assign n20733 = ~n20732;
  assign n20784 = n20736 & n2217;
  assign n20782 = ~n20818;
  assign n20785 = ~n20736;
  assign n20656 = n20833 ^ n17389;
  assign n20085 = ~n20843;
  assign n20834 = n17389 & n20844;
  assign n20831 = ~n20858;
  assign n20845 = ~n20873;
  assign n20603 = n20638 ^ n20639;
  assign n20640 = ~n20638;
  assign n20541 = ~n20661;
  assign n20644 = ~n20676;
  assign n20662 = n20596 & n20562;
  assign n20663 = ~n20596;
  assign n20643 = n20700 & n20701;
  assign n20684 = n20702 & n18026;
  assign n19371 = ~n20710;
  assign n20685 = ~n20702;
  assign n20648 = n20733 & n20734;
  assign n20719 = ~n20666;
  assign n20720 = ~n20750;
  assign n20735 = n20782 & n20783;
  assign n20738 = ~n20784;
  assign n20766 = n20785 & n92;
  assign n20790 = n20656 & n20799;
  assign n20791 = ~n20656;
  assign n20786 = n20831 & n20832;
  assign n20065 = ~n20834;
  assign n20801 = n20845 & n20846;
  assign n20524 = n20602 ^ n20603;
  assign n20505 = n20603 & n20602;
  assign n20630 = n20640 & n20641;
  assign n20510 = n20643 ^ n20644;
  assign n20564 = ~n20662;
  assign n20651 = n20663 & n20664;
  assign n20672 = n19391 & n19371;
  assign n20660 = ~n20643;
  assign n20646 = ~n20684;
  assign n20680 = n20685 & n18031;
  assign n20703 = n20719 & n20720;
  assign n20665 = ~n20648;
  assign n20704 = n20720 & n20679;
  assign n20686 = n20735 ^ n20736;
  assign n20737 = ~n20735;
  assign n20688 = ~n20766;
  assign n20739 = n20786 ^ n20787;
  assign n20658 = ~n20790;
  assign n20768 = n20791 & n20692;
  assign n17277 = n20800 ^ n20801;
  assign n20788 = ~n20786;
  assign n20803 = n20801 & n20755;
  assign n20802 = ~n20801;
  assign n20513 = ~n20524;
  assign n20508 = ~n20505;
  assign n20608 = n20510 & n9;
  assign n20604 = ~n20630;
  assign n20606 = ~n20510;
  assign n20598 = ~n20651;
  assign n20650 = n20659 & n20660;
  assign n19389 = ~n20672;
  assign n20612 = ~n20680;
  assign n20649 = n92 ^ n20686;
  assign n20678 = ~n20703;
  assign n20667 = ~n20704;
  assign n20721 = n20737 & n20738;
  assign n20620 = n20739 ^ n20740;
  assign n20591 = n17277 ^ n20751;
  assign n20694 = ~n20768;
  assign n20753 = n17277 & n20769;
  assign n20767 = n20788 & n20789;
  assign n17264 = ~n17277;
  assign n20792 = n20802 & n20771;
  assign n20770 = ~n20803;
  assign n20572 = n20604 & n20605;
  assign n20594 = n20606 & n20607;
  assign n20484 = ~n20608;
  assign n20637 = n20612 & n20646;
  assign n20581 = n20648 ^ n20649;
  assign n20632 = ~n20650;
  assign n20588 = n20649 & n20665;
  assign n16825 = n20666 ^ n20667;
  assign n20609 = n20678 & n20679;
  assign n20689 = n20620 & n2139;
  assign n20687 = ~n20721;
  assign n20690 = ~n20620;
  assign n20706 = n20591 & n20722;
  assign n20705 = ~n20591;
  assign n20743 = n17264 & n20752;
  assign n20024 = ~n20753;
  assign n20741 = ~n20767;
  assign n20756 = n20770 & n20771;
  assign n20754 = ~n20792;
  assign n20539 = n20572 ^ n20573;
  assign n20574 = ~n20572;
  assign n20512 = ~n20594;
  assign n20595 = n20632 & n20633;
  assign n20618 = n20581 & n17944;
  assign n20610 = ~n20637;
  assign n20631 = n16825 & n20642;
  assign n20617 = ~n20581;
  assign n16822 = ~n16825;
  assign n20647 = ~n20609;
  assign n20652 = n20687 & n20688;
  assign n20654 = ~n20689;
  assign n20681 = n20690 & n91;
  assign n20695 = n20705 & n20626;
  assign n20593 = ~n20706;
  assign n20691 = n20741 & n20742;
  assign n20029 = ~n20743;
  assign n20744 = n20754 & n20755;
  assign n20723 = ~n20756;
  assign n20506 = n10 ^ n20539;
  assign n20559 = n20574 & n20575;
  assign n20561 = n20595 ^ n20596;
  assign n16668 = n20609 ^ n20610;
  assign n20597 = ~n20595;
  assign n20613 = n20617 & n17975;
  assign n20583 = ~n20618;
  assign n20616 = n16822 & n19349;
  assign n19328 = ~n20631;
  assign n20599 = n16822 & n19271;
  assign n20634 = n20646 & n20647;
  assign n20619 = n91 ^ n20652;
  assign n20653 = ~n20652;
  assign n20622 = ~n20681;
  assign n20655 = n20691 ^ n20692;
  assign n20628 = ~n20695;
  assign n20696 = n20029 & n20024;
  assign n20693 = ~n20691;
  assign n20709 = n20723 & n20724;
  assign n20707 = ~n20744;
  assign n20459 = n20505 ^ n20506;
  assign n20507 = ~n20506;
  assign n20540 = ~n20559;
  assign n20461 = n20561 ^ n20562;
  assign n20576 = n16668 & n20586;
  assign n20587 = n20597 & n20598;
  assign n16777 = ~n16668;
  assign n20578 = n20599 ^ n18021;
  assign n20546 = ~n20613;
  assign n19351 = ~n20616;
  assign n20589 = n20619 ^ n20620;
  assign n20611 = ~n20634;
  assign n20645 = n20653 & n20654;
  assign n20635 = n20655 ^ n20656;
  assign n20682 = n20693 & n20694;
  assign n20044 = ~n20696;
  assign n20697 = n20707 & n20708;
  assign n20669 = ~n20709;
  assign n20470 = ~n20459;
  assign n20454 = n20507 & n20508;
  assign n20509 = n20540 & n20541;
  assign n20534 = n20461 & n20542;
  assign n20535 = ~n20461;
  assign n19290 = ~n20576;
  assign n20560 = n16777 & n20577;
  assign n20544 = n16777 & n19260;
  assign n20568 = n20578 & n20579;
  assign n20563 = ~n20587;
  assign n20565 = n20588 ^ n20589;
  assign n20566 = ~n20578;
  assign n20521 = n20589 & n20588;
  assign n20580 = n20611 & n20612;
  assign n20624 = n20635 & n90;
  assign n20621 = ~n20645;
  assign n20623 = ~n20635;
  assign n20657 = ~n20682;
  assign n20668 = ~n20697;
  assign n20457 = ~n20454;
  assign n20482 = n20509 ^ n20510;
  assign n20511 = ~n20509;
  assign n20463 = ~n20534;
  assign n20525 = n20535 & n8;
  assign n20527 = n20544 ^ n18026;
  assign n19309 = ~n20560;
  assign n20502 = n20563 & n20564;
  assign n20551 = n20565 & n17885;
  assign n20553 = n20566 & n20567;
  assign n20500 = ~n20568;
  assign n20543 = n20580 ^ n20581;
  assign n20552 = ~n20565;
  assign n20582 = ~n20580;
  assign n20548 = n20621 & n20622;
  assign n20614 = n20623 & n2082;
  assign n20555 = ~n20624;
  assign n20625 = n20657 & n20658;
  assign n17110 = n20668 & n20669;
  assign n20455 = n9 ^ n20482;
  assign n20497 = n20511 & n20512;
  assign n20435 = ~n20525;
  assign n20515 = n20527 & n20528;
  assign n20516 = ~n20527;
  assign n19306 = n19309 & n19290;
  assign n16723 = n20543 ^ n17975;
  assign n20536 = ~n20502;
  assign n20490 = ~n20551;
  assign n20547 = n20552 & n17939;
  assign n20537 = ~n20553;
  assign n20569 = n20582 & n20583;
  assign n20584 = ~n20548;
  assign n20585 = ~n20614;
  assign n20590 = n20625 ^ n20626;
  assign n20601 = n17110 ^ n20636;
  assign n20627 = ~n20625;
  assign n18701 = ~n17110;
  assign n20408 = n20454 ^ n20455;
  assign n20456 = ~n20455;
  assign n20483 = ~n20497;
  assign n20448 = ~n20515;
  assign n20503 = n20516 & n20517;
  assign n20514 = n16723 & n20524;
  assign n20526 = n20536 & n20537;
  assign n16636 = ~n16723;
  assign n20501 = n20500 & n20537;
  assign n20519 = ~n20547;
  assign n20545 = ~n20569;
  assign n20570 = n20584 & n20585;
  assign n20571 = n20585 & n20555;
  assign n20530 = n20590 ^ n20591;
  assign n19995 = n20600 ^ n20601;
  assign n20615 = n20627 & n20628;
  assign n20558 = n18701 ^ n20629;
  assign n20395 = ~n20408;
  assign n20406 = n20456 & n20457;
  assign n20460 = n20483 & n20484;
  assign n20410 = n20501 ^ n20502;
  assign n20476 = ~n20503;
  assign n20498 = n16636 & n20513;
  assign n19243 = ~n20514;
  assign n20486 = n16636 & n19211;
  assign n20499 = ~n20526;
  assign n20520 = n20519 & n20490;
  assign n20487 = n20545 & n20546;
  assign n20550 = n20530 & n89;
  assign n20554 = ~n20570;
  assign n20549 = ~n20571;
  assign n20556 = ~n20530;
  assign n20003 = ~n19995;
  assign n20592 = ~n20615;
  assign n20433 = n20460 ^ n20461;
  assign n20462 = ~n20460;
  assign n20478 = n20410 & n20485;
  assign n20399 = n20486 ^ n17944;
  assign n20466 = n20448 & n20476;
  assign n20479 = ~n20410;
  assign n19269 = ~n20498;
  assign n20467 = n20499 & n20500;
  assign n20488 = ~n20520;
  assign n20518 = ~n20487;
  assign n20522 = n20548 ^ n20549;
  assign n20496 = ~n20550;
  assign n20529 = n20554 & n20555;
  assign n20538 = n20556 & n2029;
  assign n20557 = n20592 & n20593;
  assign n20407 = n8 ^ n20433;
  assign n20446 = n20462 & n20463;
  assign n20345 = n20466 ^ n20467;
  assign n20465 = n20399 & n20471;
  assign n20412 = ~n20478;
  assign n20473 = n20479 & n23;
  assign n20464 = ~n20399;
  assign n19266 = n19243 & n19269;
  assign n16561 = n20487 ^ n20488;
  assign n20477 = ~n20467;
  assign n20504 = n20518 & n20519;
  assign n20493 = n20521 ^ n20522;
  assign n20474 = n20522 & n20521;
  assign n20494 = n20529 ^ n20530;
  assign n20532 = ~n20538;
  assign n20531 = ~n20529;
  assign n20533 = n20557 ^ n20558;
  assign n19127 = n20406 ^ n20407;
  assign n20365 = n20407 & n20406;
  assign n20436 = n20345 & n20442;
  assign n20434 = ~n20446;
  assign n20437 = ~n20345;
  assign n20449 = n20464 & n20425;
  assign n20401 = ~n20465;
  assign n20458 = n16561 & n20470;
  assign n20388 = ~n20473;
  assign n20472 = n20476 & n20477;
  assign n16673 = ~n16561;
  assign n20491 = n20493 & n17864;
  assign n20475 = n89 ^ n20494;
  assign n20489 = ~n20504;
  assign n20492 = ~n20493;
  assign n20480 = ~n20474;
  assign n20523 = n20531 & n20532;
  assign n20430 = n88 ^ n20533;
  assign n20375 = ~n19127;
  assign n20368 = ~n20365;
  assign n20409 = n20434 & n20435;
  assign n20372 = ~n20436;
  assign n20428 = n20437 & n22;
  assign n20426 = ~n20449;
  assign n19208 = ~n20458;
  assign n20445 = n16673 & n20459;
  assign n20438 = n16673 & n19170;
  assign n20447 = ~n20472;
  assign n20417 = n20474 ^ n20475;
  assign n20451 = n20475 & n20480;
  assign n20431 = n20489 & n20490;
  assign n20440 = ~n20491;
  assign n20481 = n20492 & n17862;
  assign n20495 = ~n20523;
  assign n20386 = n20409 ^ n20410;
  assign n20411 = ~n20409;
  assign n20347 = ~n20428;
  assign n20421 = n20438 ^ n17939;
  assign n19227 = ~n20445;
  assign n20424 = n20447 & n20448;
  assign n20443 = n20417 & n17772;
  assign n20444 = ~n20417;
  assign n20468 = ~n20431;
  assign n20469 = ~n20481;
  assign n20450 = n20495 & n20496;
  assign n20366 = n23 ^ n20386;
  assign n20397 = n20411 & n20412;
  assign n20413 = n20421 & n20422;
  assign n20398 = n20424 ^ n20425;
  assign n20414 = ~n20421;
  assign n20423 = n19227 & n19208;
  assign n20427 = ~n20424;
  assign n20392 = ~n20443;
  assign n20441 = n20444 & n17877;
  assign n20429 = n20450 ^ n20451;
  assign n20452 = n20468 & n20469;
  assign n20453 = n20469 & n20440;
  assign n19107 = n20365 ^ n20366;
  assign n20367 = ~n20366;
  assign n20387 = ~n20397;
  assign n20389 = n20398 ^ n20399;
  assign n20357 = ~n20413;
  assign n20404 = n20414 & n20415;
  assign n19225 = ~n20423;
  assign n20420 = n20426 & n20427;
  assign n20364 = n20429 ^ n20430;
  assign n20419 = ~n20441;
  assign n20439 = ~n20452;
  assign n20432 = ~n20453;
  assign n20309 = ~n19107;
  assign n20317 = n20367 & n20368;
  assign n20370 = n20387 & n20388;
  assign n20380 = n20389 & n21;
  assign n20378 = ~n20389;
  assign n20382 = ~n20404;
  assign n20403 = n20364 & n17835;
  assign n20400 = ~n20420;
  assign n20402 = ~n20364;
  assign n16641 = n20431 ^ n20432;
  assign n20416 = n20439 & n20440;
  assign n20328 = ~n20317;
  assign n20344 = n22 ^ n20370;
  assign n20371 = ~n20370;
  assign n20376 = n20378 & n20379;
  assign n20303 = ~n20380;
  assign n20383 = n20357 & n20382;
  assign n20358 = n20400 & n20401;
  assign n20394 = n20402 & n17750;
  assign n20350 = ~n20403;
  assign n20396 = n16641 & n20408;
  assign n20390 = n20416 ^ n20417;
  assign n16500 = ~n16641;
  assign n20418 = ~n20416;
  assign n20318 = n20344 ^ n20345;
  assign n20355 = n20371 & n20372;
  assign n20322 = ~n20376;
  assign n20359 = ~n20383;
  assign n16566 = n17772 ^ n20390;
  assign n20381 = ~n20358;
  assign n20373 = ~n20394;
  assign n20393 = n16500 & n20395;
  assign n19167 = ~n20396;
  assign n20384 = n16500 & n19063;
  assign n20405 = n20418 & n20419;
  assign n19072 = n20317 ^ n20318;
  assign n20300 = n20318 & n20328;
  assign n20346 = ~n20355;
  assign n20351 = n20322 & n20303;
  assign n20348 = n20358 ^ n20359;
  assign n20369 = n16566 & n20375;
  assign n20352 = n16566 & n19047;
  assign n20377 = n20381 & n20382;
  assign n16575 = ~n16566;
  assign n20313 = n20384 ^ n17862;
  assign n19189 = ~n20393;
  assign n20391 = ~n20405;
  assign n20299 = ~n19072;
  assign n20319 = n20346 & n20347;
  assign n20342 = n20348 & n20;
  assign n20320 = ~n20351;
  assign n20334 = n20352 ^ n17877;
  assign n20340 = ~n20348;
  assign n20354 = n16575 & n19127;
  assign n19150 = ~n20369;
  assign n20361 = n20313 & n20374;
  assign n20356 = ~n20377;
  assign n20362 = ~n20313;
  assign n19186 = n19189 & n19167;
  assign n20385 = n20391 & n20392;
  assign n20301 = n20319 ^ n20320;
  assign n20321 = ~n20319;
  assign n20329 = n20334 & n20335;
  assign n20333 = n20340 & n20341;
  assign n20258 = ~n20342;
  assign n20330 = ~n20334;
  assign n19130 = ~n20354;
  assign n20336 = n20356 & n20357;
  assign n20315 = ~n20361;
  assign n20353 = n20362 & n20337;
  assign n20363 = ~n20385;
  assign n20251 = n20300 ^ n20301;
  assign n20253 = n20301 & n20300;
  assign n20311 = n20321 & n20322;
  assign n20273 = ~n20329;
  assign n20323 = n20330 & n20331;
  assign n20279 = ~n20333;
  assign n20312 = n20336 ^ n20337;
  assign n20338 = ~n20336;
  assign n20339 = ~n20353;
  assign n20343 = n20363 ^ n20364;
  assign n20360 = n20363 & n20373;
  assign n20265 = ~n20251;
  assign n20256 = ~n20253;
  assign n20302 = ~n20311;
  assign n20219 = n20312 ^ n20313;
  assign n20308 = n20279 & n20258;
  assign n20298 = ~n20323;
  assign n20332 = n20338 & n20339;
  assign n16480 = n20343 ^ n17750;
  assign n20349 = ~n20360;
  assign n20276 = n20302 & n20303;
  assign n20296 = n20219 & n19;
  assign n20294 = ~n20219;
  assign n20288 = n20273 & n20298;
  assign n20277 = ~n20308;
  assign n20310 = n16480 & n19107;
  assign n20304 = n16480 & n19045;
  assign n20314 = ~n20332;
  assign n16306 = ~n16480;
  assign n20324 = n20349 & n20350;
  assign n20254 = n20276 ^ n20277;
  assign n20278 = ~n20276;
  assign n20287 = n20294 & n20295;
  assign n20221 = ~n20296;
  assign n20233 = n20304 ^ n17750;
  assign n20307 = n16306 & n20309;
  assign n19109 = ~n20310;
  assign n20289 = n20314 & n20315;
  assign n16396 = n20324 ^ n20325;
  assign n20326 = ~n20324;
  assign n18961 = n20253 ^ n20254;
  assign n20255 = ~n20254;
  assign n20270 = n20278 & n20279;
  assign n20239 = ~n20287;
  assign n20181 = n20288 ^ n20289;
  assign n20281 = n20233 & n20290;
  assign n20280 = ~n20233;
  assign n20293 = n16396 & n20299;
  assign n19092 = ~n20307;
  assign n20297 = ~n20289;
  assign n16384 = ~n16396;
  assign n20316 = n20326 & n20327;
  assign n20203 = ~n18961;
  assign n20195 = n20255 & n20256;
  assign n20257 = ~n20270;
  assign n20266 = n20181 & n20271;
  assign n20267 = ~n20181;
  assign n20274 = n20280 & n20247;
  assign n20235 = ~n20281;
  assign n19054 = ~n20293;
  assign n20291 = n20297 & n20298;
  assign n20292 = n16384 & n19072;
  assign n20282 = n16384 & n18920;
  assign n20305 = ~n20316;
  assign n20198 = ~n20195;
  assign n20237 = n20257 & n20258;
  assign n20201 = ~n20266;
  assign n20259 = n20267 & n18;
  assign n20249 = ~n20274;
  assign n20268 = n20282 ^ n17776;
  assign n20272 = ~n20291;
  assign n19074 = ~n20292;
  assign n20284 = n20305 & n20306;
  assign n20218 = n19 ^ n20237;
  assign n20238 = ~n20237;
  assign n20183 = ~n20259;
  assign n20260 = n20268 & n20269;
  assign n20246 = n20272 & n20273;
  assign n20261 = ~n20268;
  assign n16170 = n20283 ^ n20284;
  assign n20285 = ~n20284;
  assign n20196 = n20218 ^ n20219;
  assign n20231 = n20238 & n20239;
  assign n20232 = n20246 ^ n20247;
  assign n20193 = ~n20260;
  assign n20250 = n20261 & n20262;
  assign n20252 = n16170 & n20265;
  assign n20248 = ~n20246;
  assign n20243 = n16170 & n18978;
  assign n16355 = ~n16170;
  assign n20275 = n20285 & n20286;
  assign n20178 = n20195 ^ n20196;
  assign n20197 = ~n20196;
  assign n20220 = ~n20231;
  assign n20222 = n20232 ^ n20233;
  assign n20147 = n20243 ^ n17733;
  assign n20244 = n20248 & n20249;
  assign n20217 = ~n20250;
  assign n20245 = n16355 & n20251;
  assign n19030 = ~n20252;
  assign n20263 = ~n20275;
  assign n20179 = ~n20178;
  assign n20152 = n20197 & n20198;
  assign n20199 = n20220 & n20221;
  assign n20213 = n20222 & n17;
  assign n20211 = ~n20222;
  assign n20228 = n20147 & n20175;
  assign n20214 = n20217 & n20193;
  assign n20229 = ~n20147;
  assign n20234 = ~n20244;
  assign n19007 = ~n20245;
  assign n20240 = n20263 & n20264;
  assign n20155 = ~n20152;
  assign n20180 = n18 ^ n20199;
  assign n20200 = ~n20199;
  assign n20209 = n20211 & n20212;
  assign n20136 = ~n20213;
  assign n20177 = ~n20228;
  assign n20223 = n20229 & n20230;
  assign n20215 = n20234 & n20235;
  assign n19027 = n19030 & n19007;
  assign n20224 = n20240 ^ n17588;
  assign n20241 = ~n20240;
  assign n20153 = n20180 ^ n20181;
  assign n20188 = n20200 & n20201;
  assign n20159 = ~n20209;
  assign n20094 = n20214 ^ n20215;
  assign n20150 = ~n20223;
  assign n16215 = n20224 ^ n20225;
  assign n20216 = ~n20215;
  assign n20236 = n20241 & n20242;
  assign n18884 = n20152 ^ n20153;
  assign n20154 = ~n20153;
  assign n20182 = ~n20188;
  assign n20156 = n20159 & n20136;
  assign n20190 = n20094 & n20204;
  assign n20202 = n16215 & n18961;
  assign n20186 = n16215 & n18917;
  assign n20191 = ~n20094;
  assign n20210 = n20216 & n20217;
  assign n16231 = ~n16215;
  assign n20226 = ~n20236;
  assign n20129 = ~n18884;
  assign n20131 = n20154 & n20155;
  assign n20157 = n20182 & n20183;
  assign n20172 = n20186 ^ n17588;
  assign n20115 = ~n20190;
  assign n20187 = n20191 & n16;
  assign n18987 = ~n20202;
  assign n20189 = n16231 & n20203;
  assign n20192 = ~n20210;
  assign n20206 = n20226 & n20227;
  assign n20134 = ~n20131;
  assign n20132 = n20156 ^ n20157;
  assign n20158 = ~n20157;
  assign n20167 = n20172 & n20173;
  assign n20165 = ~n20172;
  assign n20096 = ~n20187;
  assign n18964 = ~n20189;
  assign n20174 = n20192 & n20193;
  assign n16174 = n20205 ^ n20206;
  assign n20207 = ~n20206;
  assign n20077 = n20131 ^ n20132;
  assign n20133 = ~n20132;
  assign n20145 = n20158 & n20159;
  assign n20160 = n20165 & n20166;
  assign n20110 = ~n20167;
  assign n20146 = n20174 ^ n20175;
  assign n20171 = n16174 & n20179;
  assign n20176 = ~n20174;
  assign n20168 = n16174 & n18890;
  assign n16186 = ~n16174;
  assign n20194 = n20207 & n20208;
  assign n20086 = ~n20077;
  assign n20075 = n20133 & n20134;
  assign n20135 = ~n20145;
  assign n20080 = n20146 ^ n20147;
  assign n20128 = ~n20160;
  assign n20069 = n20168 ^ n17574;
  assign n18949 = ~n20171;
  assign n20169 = n20176 & n20177;
  assign n20170 = n16186 & n20178;
  assign n20184 = ~n20194;
  assign n20113 = n20135 & n20136;
  assign n20125 = n20080 & n20137;
  assign n20138 = n20128 & n20110;
  assign n20126 = ~n20080;
  assign n20142 = n20069 & n20148;
  assign n20143 = ~n20069;
  assign n20149 = ~n20169;
  assign n18928 = ~n20170;
  assign n20162 = n20184 & n20185;
  assign n20093 = n16 ^ n20113;
  assign n20114 = ~n20113;
  assign n20082 = ~n20125;
  assign n20121 = n20126 & n31;
  assign n20117 = ~n20138;
  assign n20073 = ~n20142;
  assign n20139 = n20143 & n20090;
  assign n20116 = n20149 & n20150;
  assign n20144 = n18949 & n18928;
  assign n16064 = n20161 ^ n20162;
  assign n20163 = ~n20162;
  assign n20076 = n20093 ^ n20094;
  assign n20108 = n20114 & n20115;
  assign n20105 = n20116 ^ n20117;
  assign n20061 = ~n20121;
  assign n20092 = ~n20139;
  assign n20130 = n16064 & n18884;
  assign n20127 = ~n20116;
  assign n20123 = n16064 & n18833;
  assign n18947 = ~n20144;
  assign n16091 = ~n16064;
  assign n20151 = n20163 & n20164;
  assign n18793 = n20075 ^ n20076;
  assign n20037 = n20076 & n20075;
  assign n20099 = n20105 & n30;
  assign n20095 = ~n20108;
  assign n20097 = ~n20105;
  assign n20055 = n20123 ^ n17543;
  assign n20122 = n20127 & n20128;
  assign n20124 = n16091 & n20129;
  assign n18909 = ~n20130;
  assign n20140 = ~n20151;
  assign n20048 = ~n18793;
  assign n20079 = n20095 & n20096;
  assign n20088 = n20097 & n20098;
  assign n20021 = ~n20099;
  assign n20106 = n20055 & n20111;
  assign n20107 = ~n20055;
  assign n20109 = ~n20122;
  assign n18887 = ~n20124;
  assign n20118 = n20140 & n20141;
  assign n20058 = n20079 ^ n20080;
  assign n20081 = ~n20079;
  assign n20043 = ~n20088;
  assign n20057 = ~n20106;
  assign n20100 = n20107 & n20032;
  assign n20089 = n20109 & n20110;
  assign n20101 = n20118 ^ n17435;
  assign n20119 = ~n20118;
  assign n20038 = n31 ^ n20058;
  assign n20070 = n20081 & n20082;
  assign n20071 = n20043 & n20021;
  assign n20068 = n20089 ^ n20090;
  assign n20035 = ~n20100;
  assign n16004 = n20101 ^ n20102;
  assign n20091 = ~n20089;
  assign n20112 = n20119 & n20120;
  assign n18765 = n20037 ^ n20038;
  assign n20017 = n20038 & n20037;
  assign n20059 = n20068 ^ n20069;
  assign n20060 = ~n20070;
  assign n20041 = ~n20071;
  assign n20078 = n16004 & n20086;
  assign n20066 = n16004 & n18808;
  assign n20087 = n20091 & n20092;
  assign n16015 = ~n16004;
  assign n20103 = ~n20112;
  assign n20016 = ~n18765;
  assign n20053 = n20059 & n29;
  assign n20040 = n20060 & n20061;
  assign n20051 = ~n20059;
  assign n19982 = n20066 ^ n17435;
  assign n20067 = n16015 & n20077;
  assign n18867 = ~n20078;
  assign n20072 = ~n20087;
  assign n20083 = n20103 & n20104;
  assign n20018 = n20040 ^ n20041;
  assign n20049 = n20051 & n20052;
  assign n19973 = ~n20053;
  assign n20042 = ~n20040;
  assign n18846 = ~n20067;
  assign n20054 = n20072 & n20073;
  assign n20063 = n20083 ^ n17236;
  assign n20084 = ~n20083;
  assign n19950 = n20017 ^ n20018;
  assign n19967 = n20018 & n20017;
  assign n20033 = n20042 & n20043;
  assign n19990 = ~n20049;
  assign n20031 = n20054 ^ n20055;
  assign n18864 = n18867 & n18846;
  assign n15745 = n20062 ^ n20063;
  assign n20056 = ~n20054;
  assign n20074 = n20084 & n20085;
  assign n19970 = ~n19967;
  assign n20026 = n19990 & n19973;
  assign n20019 = n20031 ^ n20032;
  assign n20020 = ~n20033;
  assign n20039 = n15745 & n20048;
  assign n20027 = n15745 & n18669;
  assign n20050 = n20056 & n20057;
  assign n15913 = ~n15745;
  assign n20064 = ~n20074;
  assign n20007 = n20019 & n28;
  assign n19987 = n20020 & n20021;
  assign n19988 = ~n20026;
  assign n20005 = ~n20019;
  assign n20008 = n20027 ^ n17236;
  assign n20030 = n15913 & n18793;
  assign n18822 = ~n20039;
  assign n20034 = ~n20050;
  assign n20045 = n20064 & n20065;
  assign n19968 = n19987 ^ n19988;
  assign n19997 = n20005 & n20006;
  assign n19941 = ~n20007;
  assign n19989 = ~n19987;
  assign n19998 = n20008 & n20009;
  assign n19999 = ~n20008;
  assign n18796 = ~n20030;
  assign n20010 = n20034 & n20035;
  assign n15838 = n20044 ^ n20045;
  assign n20047 = n20045 & n20024;
  assign n20046 = ~n20045;
  assign n18873 = n19967 ^ n19968;
  assign n19969 = ~n19968;
  assign n19984 = n19989 & n19990;
  assign n19957 = ~n19997;
  assign n19946 = ~n19998;
  assign n19992 = n19999 & n20000;
  assign n19983 = n20010 ^ n20011;
  assign n20013 = n20010 & n20022;
  assign n20015 = n15838 & n18765;
  assign n20012 = ~n20010;
  assign n15826 = ~n15838;
  assign n20036 = n20046 & n20029;
  assign n20028 = ~n20047;
  assign n16779 = n18873 ^ n19916;
  assign n18825 = n18873 ^ n19947;
  assign n19953 = ~n18873;
  assign n19936 = n19969 & n19970;
  assign n19954 = n19957 & n19941;
  assign n19922 = n19982 ^ n19983;
  assign n19972 = ~n19984;
  assign n19961 = ~n19992;
  assign n20001 = n20012 & n20011;
  assign n19991 = ~n20013;
  assign n18741 = ~n20015;
  assign n20004 = n15826 & n20016;
  assign n19993 = n15826 & n18619;
  assign n20025 = n20028 & n20029;
  assign n20023 = ~n20036;
  assign n19934 = n16779 & n19947;
  assign n18824 = ~n16779;
  assign n19875 = n19953 & n17799;
  assign n19939 = ~n19936;
  assign n19964 = n19922 & n19971;
  assign n19955 = n19972 & n19973;
  assign n19965 = ~n19922;
  assign n19976 = n19961 & n19946;
  assign n19985 = n19991 & n19982;
  assign n19904 = n19993 ^ n17264;
  assign n19975 = ~n20001;
  assign n18767 = ~n20004;
  assign n20014 = n20023 & n20024;
  assign n20002 = ~n20025;
  assign n19869 = ~n19934;
  assign n19915 = n18824 & n18803;
  assign n19932 = n18824 & n19935;
  assign n19937 = n19954 ^ n19955;
  assign n19924 = ~n19964;
  assign n19962 = n19965 & n27;
  assign n19956 = ~n19955;
  assign n19959 = ~n19976;
  assign n19977 = n19904 & n19981;
  assign n19974 = ~n19985;
  assign n19978 = ~n19904;
  assign n19996 = n20002 & n20003;
  assign n19994 = ~n20014;
  assign n19909 = n19915 ^ n19916;
  assign n19917 = ~n19915;
  assign n19899 = ~n19932;
  assign n19929 = n19936 ^ n19937;
  assign n19938 = ~n19937;
  assign n19951 = n19956 & n19957;
  assign n19906 = ~n19962;
  assign n19958 = n19974 & n19975;
  assign n19908 = ~n19977;
  assign n19966 = n19978 & n19926;
  assign n19986 = n19994 & n19995;
  assign n19980 = ~n19996;
  assign n19889 = n19909 & n19910;
  assign n19911 = n19917 & n19918;
  assign n19919 = n19929 & n17679;
  assign n19920 = ~n19929;
  assign n19872 = n19938 & n19939;
  assign n19940 = ~n19951;
  assign n19948 = n19958 ^ n19959;
  assign n19960 = ~n19958;
  assign n19928 = ~n19966;
  assign n19979 = ~n19986;
  assign n19824 = n19889 ^ n19890;
  assign n19893 = n19889 & n19890;
  assign n19891 = ~n19889;
  assign n19898 = ~n19911;
  assign n19877 = ~n19919;
  assign n19912 = n19920 & n17672;
  assign n19879 = ~n19872;
  assign n19921 = n19940 & n19941;
  assign n19944 = n19948 & n26;
  assign n19942 = ~n19948;
  assign n19952 = n19960 & n19961;
  assign n15611 = n19979 & n19980;
  assign n19867 = n19891 & n19892;
  assign n19817 = ~n19893;
  assign n19895 = n19898 & n19899;
  assign n19896 = n19898 & n19900;
  assign n19901 = ~n19912;
  assign n19902 = n19921 ^ n19922;
  assign n19923 = ~n19921;
  assign n19933 = n19942 & n19943;
  assign n19860 = ~n19944;
  assign n19945 = ~n19952;
  assign n19949 = n15611 & n19963;
  assign n17227 = ~n15611;
  assign n19831 = ~n19867;
  assign n19870 = ~n19895;
  assign n19868 = ~n19896;
  assign n19897 = n19901 & n19875;
  assign n19874 = n19901 & n19877;
  assign n19873 = n27 ^ n19902;
  assign n19913 = n19923 & n19924;
  assign n19886 = ~n19933;
  assign n19925 = n19945 & n19946;
  assign n19930 = n19949 ^ n17110;
  assign n18722 = n19950 ^ n17227;
  assign n19862 = n19868 & n19869;
  assign n19863 = n19870 & n19871;
  assign n19861 = n19872 ^ n19873;
  assign n16753 = n19874 ^ n19875;
  assign n19876 = ~n19897;
  assign n19878 = ~n19873;
  assign n19905 = ~n19913;
  assign n19883 = n19886 & n19860;
  assign n19903 = n19925 ^ n19926;
  assign n19888 = n19930 ^ n19931;
  assign n19927 = ~n19925;
  assign n19856 = n19861 & n17619;
  assign n19854 = ~n19862;
  assign n19843 = ~n19863;
  assign n19834 = ~n19861;
  assign n16755 = ~n16753;
  assign n19864 = n19876 & n19877;
  assign n19857 = n19878 & n19879;
  assign n19894 = n19903 ^ n19904;
  assign n19884 = n19905 & n19906;
  assign n19914 = n19927 & n19928;
  assign n19851 = n19854 & n19855;
  assign n19852 = n19834 & n17625;
  assign n19848 = ~n19856;
  assign n19840 = n16755 & n18772;
  assign n19849 = ~n19864;
  assign n19858 = n19883 ^ n19884;
  assign n19882 = n19894 & n25;
  assign n19880 = ~n19894;
  assign n19885 = ~n19884;
  assign n19907 = ~n19914;
  assign n19825 = n19840 ^ n17672;
  assign n19841 = n19848 & n19849;
  assign n19842 = ~n19851;
  assign n19833 = ~n19852;
  assign n19835 = n19849 ^ n17625;
  assign n19850 = n19857 ^ n19858;
  assign n19821 = n19858 & n19857;
  assign n19865 = n19880 & n19881;
  assign n19830 = ~n19882;
  assign n19866 = n19885 & n19886;
  assign n19887 = n19907 & n19908;
  assign n19815 = n19824 ^ n19825;
  assign n19826 = n19831 & n19825;
  assign n16590 = n19834 ^ n19835;
  assign n19832 = ~n19841;
  assign n19827 = n19842 & n19843;
  assign n19845 = n19850 & n17562;
  assign n19844 = ~n19850;
  assign n19847 = ~n19865;
  assign n19859 = ~n19866;
  assign n19814 = n19887 ^ n19888;
  assign n19810 = n19815 & n230;
  assign n19808 = ~n19815;
  assign n19816 = ~n19826;
  assign n18304 = n231 ^ n19827;
  assign n19804 = n19832 & n19833;
  assign n16643 = ~n16590;
  assign n19828 = ~n19827;
  assign n19836 = n19844 & n17459;
  assign n19819 = ~n19845;
  assign n19853 = n19847 & n19830;
  assign n19837 = n19859 & n19860;
  assign n19802 = n19808 & n19809;
  assign n19783 = ~n19810;
  assign n19758 = n19816 & n19817;
  assign n19803 = n16643 & n18636;
  assign n19818 = ~n19804;
  assign n19775 = n19828 & n231;
  assign n19800 = ~n19836;
  assign n19838 = ~n19853;
  assign n19846 = ~n19837;
  assign n19795 = ~n19802;
  assign n19796 = n19803 ^ n17619;
  assign n19778 = ~n19758;
  assign n19811 = n19818 & n19819;
  assign n19820 = n19819 & n19800;
  assign n19822 = n19837 ^ n19838;
  assign n19839 = n19846 & n19847;
  assign n19790 = n19775 & n19795;
  assign n19791 = n19795 & n19783;
  assign n19792 = n19796 & n19797;
  assign n19793 = ~n19796;
  assign n19799 = ~n19811;
  assign n19805 = ~n19820;
  assign n19812 = n19821 ^ n19822;
  assign n19823 = ~n19822;
  assign n19829 = ~n19839;
  assign n19782 = ~n19790;
  assign n19776 = ~n19791;
  assign n19764 = ~n19792;
  assign n19787 = n19793 & n19794;
  assign n19781 = n19799 & n19800;
  assign n16539 = n19804 ^ n19805;
  assign n19807 = n19812 & n17375;
  assign n19806 = ~n19812;
  assign n19785 = n19823 & n19821;
  assign n19813 = n19829 & n19830;
  assign n19762 = n19775 ^ n19776;
  assign n19711 = n19782 & n19783;
  assign n19777 = ~n19787;
  assign n19788 = ~n19781;
  assign n16532 = ~n16539;
  assign n19801 = n19806 & n17462;
  assign n19774 = ~n19807;
  assign n19798 = n19813 ^ n19814;
  assign n19531 = n19762 ^ n18304;
  assign n19691 = n19762 & n18304;
  assign n19771 = n19777 & n19778;
  assign n19728 = ~n19711;
  assign n19772 = n19777 & n19764;
  assign n19779 = n16532 & n18520;
  assign n19786 = n24 ^ n19798;
  assign n19789 = ~n19801;
  assign n19519 = ~n19531;
  assign n19763 = ~n19771;
  assign n19759 = ~n19772;
  assign n19731 = n19779 ^ n17562;
  assign n19746 = n19785 ^ n19786;
  assign n19784 = n19788 & n19789;
  assign n19780 = n19789 & n19774;
  assign n19749 = n19758 ^ n19759;
  assign n19750 = n19763 & n19764;
  assign n19766 = n19731 & n19768;
  assign n19765 = ~n19731;
  assign n19770 = n19746 & n17295;
  assign n16441 = n19780 ^ n19781;
  assign n19769 = ~n19746;
  assign n19773 = ~n19784;
  assign n19745 = n19749 & n229;
  assign n19730 = n19750 ^ n19751;
  assign n19741 = ~n19749;
  assign n19753 = ~n19750;
  assign n19760 = n19765 & n19751;
  assign n19733 = ~n19766;
  assign n19755 = n16441 & n18532;
  assign n19767 = n19769 & n17405;
  assign n19740 = ~n19770;
  assign n19761 = n19773 & n19774;
  assign n16455 = ~n16441;
  assign n19722 = n19730 ^ n19731;
  assign n19735 = n19741 & n19742;
  assign n19713 = ~n19745;
  assign n19743 = n19755 ^ n17462;
  assign n19752 = ~n19760;
  assign n19747 = n19761 ^ n17295;
  assign n19757 = ~n19767;
  assign n19756 = ~n19761;
  assign n19717 = n19722 & n228;
  assign n19715 = ~n19722;
  assign n19729 = ~n19735;
  assign n19736 = n19743 & n19744;
  assign n16390 = n19746 ^ n19747;
  assign n19748 = n19752 & n19753;
  assign n19737 = ~n19743;
  assign n19754 = n19756 & n19757;
  assign n19709 = n19715 & n19716;
  assign n19676 = ~n19717;
  assign n19723 = n19728 & n19729;
  assign n19710 = n19729 & n19713;
  assign n19718 = n16390 & n18491;
  assign n19701 = ~n19736;
  assign n19734 = n19737 & n19738;
  assign n16402 = ~n16390;
  assign n19732 = ~n19748;
  assign n19739 = ~n19754;
  assign n19694 = ~n19709;
  assign n19692 = n19710 ^ n19711;
  assign n19702 = n19718 ^ n17405;
  assign n19712 = ~n19723;
  assign n19705 = n19732 & n19733;
  assign n19719 = ~n19734;
  assign n19724 = n19739 & n19740;
  assign n18267 = n19691 ^ n19692;
  assign n19678 = n19694 & n19676;
  assign n19665 = n19692 & n19691;
  assign n19697 = n19702 & n19703;
  assign n19698 = ~n19702;
  assign n19679 = n19712 & n19713;
  assign n19704 = n19719 & n19701;
  assign n19706 = n19724 ^ n19725;
  assign n19720 = ~n19705;
  assign n19726 = ~n19724;
  assign n19666 = n19678 ^ n19679;
  assign n19459 = ~n18267;
  assign n19668 = ~n19665;
  assign n19670 = ~n19697;
  assign n19696 = n19698 & n19699;
  assign n19657 = n19704 ^ n19705;
  assign n19693 = ~n19679;
  assign n16178 = n19706 ^ n17216;
  assign n19714 = n19719 & n19720;
  assign n19721 = n19726 & n19727;
  assign n19442 = n19665 ^ n19666;
  assign n19667 = ~n19666;
  assign n19684 = n19693 & n19694;
  assign n19685 = n19657 & n19695;
  assign n19680 = ~n19696;
  assign n19686 = ~n19657;
  assign n16281 = ~n16178;
  assign n19700 = ~n19714;
  assign n19707 = ~n19721;
  assign n19450 = ~n19442;
  assign n19619 = n19667 & n19668;
  assign n19677 = n19680 & n19670;
  assign n19675 = ~n19684;
  assign n19661 = ~n19685;
  assign n19682 = n19686 & n227;
  assign n19671 = n16281 & n18474;
  assign n19658 = n19700 & n19701;
  assign n19687 = n19707 & n19708;
  assign n19622 = ~n19619;
  assign n19662 = n19671 ^ n17280;
  assign n19656 = n19675 & n19676;
  assign n19659 = ~n19677;
  assign n19644 = ~n19682;
  assign n16236 = n19687 ^ n19688;
  assign n19681 = ~n19658;
  assign n19689 = ~n19687;
  assign n19639 = n19656 ^ n19657;
  assign n19626 = n19658 ^ n19659;
  assign n19652 = n19662 & n19663;
  assign n19650 = ~n19662;
  assign n19660 = ~n19656;
  assign n19674 = n19680 & n19681;
  assign n16224 = ~n16236;
  assign n19683 = n19689 & n19690;
  assign n19620 = n227 ^ n19639;
  assign n19642 = n19626 & n226;
  assign n19640 = ~n19626;
  assign n19647 = n19650 & n19651;
  assign n19616 = ~n19652;
  assign n19649 = n19660 & n19661;
  assign n19653 = n16224 & n18406;
  assign n19669 = ~n19674;
  assign n19672 = ~n19683;
  assign n19387 = n19619 ^ n19620;
  assign n19621 = ~n19620;
  assign n19632 = n19640 & n19641;
  assign n19607 = ~n19642;
  assign n19633 = ~n19647;
  assign n19643 = ~n19649;
  assign n19583 = n19653 ^ n17131;
  assign n19612 = n19669 & n19670;
  assign n19664 = n19672 & n19673;
  assign n19393 = ~n19387;
  assign n19586 = n19621 & n19622;
  assign n19623 = ~n19632;
  assign n19630 = n19633 & n19616;
  assign n19625 = n19643 & n19644;
  assign n19635 = n19583 & n19645;
  assign n19636 = ~n19583;
  assign n19634 = ~n19612;
  assign n19655 = n19664 & n17096;
  assign n19654 = ~n19664;
  assign n19589 = ~n19586;
  assign n19605 = n19625 ^ n19626;
  assign n19613 = ~n19630;
  assign n19629 = n19633 & n19634;
  assign n19624 = ~n19625;
  assign n19585 = ~n19635;
  assign n19631 = n19636 & n19601;
  assign n19648 = n19654 & n17147;
  assign n19638 = ~n19655;
  assign n19587 = n226 ^ n19605;
  assign n19599 = n19612 ^ n19613;
  assign n19614 = n19623 & n19624;
  assign n19615 = ~n19629;
  assign n19603 = ~n19631;
  assign n19637 = n19638 & n19646;
  assign n19628 = ~n19648;
  assign n19373 = n19586 ^ n19587;
  assign n19588 = ~n19587;
  assign n19597 = n19599 & n225;
  assign n19595 = ~n19599;
  assign n19606 = ~n19614;
  assign n19600 = n19615 & n19616;
  assign n19627 = ~n19637;
  assign n19618 = n19628 & n19638;
  assign n19369 = ~n19373;
  assign n19537 = n19588 & n19589;
  assign n19590 = n19595 & n19596;
  assign n19560 = ~n19597;
  assign n19582 = n19600 ^ n19601;
  assign n19551 = n19606 & n19607;
  assign n19602 = ~n19600;
  assign n16110 = n19617 ^ n19618;
  assign n19608 = n19627 & n19628;
  assign n19541 = n19582 ^ n19583;
  assign n19580 = ~n19590;
  assign n19579 = ~n19551;
  assign n19598 = n19602 & n19603;
  assign n19592 = n16110 & n18363;
  assign n19591 = n19608 ^ n19609;
  assign n16121 = ~n16110;
  assign n19610 = ~n19608;
  assign n19566 = n19541 & n224;
  assign n19564 = ~n19541;
  assign n19571 = n19579 & n19580;
  assign n19572 = n19580 & n19560;
  assign n16045 = n19591 ^ n17121;
  assign n19568 = n19592 ^ n17147;
  assign n19584 = ~n19598;
  assign n19604 = n19610 & n19611;
  assign n19558 = n19564 & n19565;
  assign n19524 = ~n19566;
  assign n19559 = ~n19571;
  assign n19552 = ~n19572;
  assign n19573 = n19568 & n19581;
  assign n19561 = n16045 & n18322;
  assign n19567 = n19584 & n19585;
  assign n16058 = ~n16045;
  assign n19574 = ~n19568;
  assign n19593 = ~n19604;
  assign n19538 = n19551 ^ n19552;
  assign n19546 = ~n19558;
  assign n19553 = n19559 & n19560;
  assign n19510 = n19561 ^ n17121;
  assign n19549 = n19567 ^ n19568;
  assign n19562 = ~n19573;
  assign n19569 = n19574 & n19550;
  assign n19563 = ~n19567;
  assign n19575 = n19593 & n19594;
  assign n18099 = n19537 ^ n19538;
  assign n19497 = n19538 & n19537;
  assign n19536 = n19549 ^ n19550;
  assign n19540 = ~n19553;
  assign n19554 = n19562 & n19563;
  assign n19548 = ~n19569;
  assign n19555 = n19575 ^ n19576;
  assign n19577 = ~n19575;
  assign n19305 = ~n18099;
  assign n19534 = n19536 & n239;
  assign n19500 = ~n19497;
  assign n19516 = n19540 ^ n19541;
  assign n19539 = n19546 & n19540;
  assign n19532 = ~n19536;
  assign n19547 = ~n19554;
  assign n15973 = n19555 ^ n16979;
  assign n19570 = n19577 & n19578;
  assign n19498 = n224 ^ n19516;
  assign n19525 = n19532 & n19533;
  assign n19481 = ~n19534;
  assign n19523 = ~n19539;
  assign n19526 = n19547 & n19548;
  assign n15963 = ~n15973;
  assign n19556 = ~n19570;
  assign n19292 = n19497 ^ n19498;
  assign n19499 = ~n19498;
  assign n19489 = n19523 & n19524;
  assign n19508 = ~n19525;
  assign n19509 = n19526 ^ n19527;
  assign n19530 = n19526 & n19527;
  assign n19528 = ~n19526;
  assign n19517 = n15963 & n18233;
  assign n19543 = n19556 & n19557;
  assign n19288 = ~n19292;
  assign n19468 = n19499 & n19500;
  assign n19490 = n19509 ^ n19510;
  assign n19488 = n19508 & n19481;
  assign n19507 = ~n19489;
  assign n19471 = n19517 ^ n16979;
  assign n19518 = n19528 & n19529;
  assign n19514 = ~n19530;
  assign n15756 = n19542 ^ n19543;
  assign n19544 = ~n19543;
  assign n19469 = n19488 ^ n19489;
  assign n19484 = n19490 & n238;
  assign n19482 = ~n19490;
  assign n19501 = n19507 & n19508;
  assign n19503 = n19471 & n19511;
  assign n19512 = n19514 & n19510;
  assign n19502 = ~n19471;
  assign n19492 = ~n19518;
  assign n19513 = n15756 & n18252;
  assign n19520 = n15756 & n19531;
  assign n15874 = ~n15756;
  assign n19535 = n19544 & n19545;
  assign n18044 = n19468 ^ n19469;
  assign n19424 = n19469 & n19468;
  assign n19474 = n19482 & n19483;
  assign n19448 = ~n19484;
  assign n19480 = ~n19501;
  assign n19495 = n19502 & n19452;
  assign n19473 = ~n19503;
  assign n19491 = ~n19512;
  assign n19493 = n19513 ^ n16948;
  assign n19515 = n15874 & n19519;
  assign n18301 = ~n19520;
  assign n19521 = ~n19535;
  assign n19240 = ~n18044;
  assign n19465 = ~n19474;
  assign n19446 = n19480 & n19481;
  assign n19470 = n19491 & n19492;
  assign n19485 = n19493 & n19494;
  assign n19454 = ~n19495;
  assign n19486 = ~n19493;
  assign n18284 = ~n19515;
  assign n19504 = n19521 & n19522;
  assign n19445 = n19465 & n19448;
  assign n19451 = n19470 ^ n19471;
  assign n19466 = ~n19446;
  assign n19472 = ~n19470;
  assign n19417 = ~n19485;
  assign n19475 = n19486 & n19487;
  assign n18298 = n18301 & n18284;
  assign n19477 = n19504 ^ n16963;
  assign n19505 = ~n19504;
  assign n19425 = n19445 ^ n19446;
  assign n19440 = n19451 ^ n19452;
  assign n19457 = n19465 & n19466;
  assign n19467 = n19472 & n19473;
  assign n19438 = ~n19475;
  assign n15787 = n19476 ^ n19477;
  assign n19496 = n19505 & n19506;
  assign n19205 = n19424 ^ n19425;
  assign n19374 = n19425 & n19424;
  assign n19433 = n19440 & n237;
  assign n19431 = ~n19440;
  assign n19447 = ~n19457;
  assign n19453 = ~n19467;
  assign n19458 = n19438 & n19417;
  assign n19449 = n15787 & n18174;
  assign n19460 = n15787 & n18267;
  assign n15799 = ~n15787;
  assign n19478 = ~n19496;
  assign n18011 = ~n19205;
  assign n19426 = n19431 & n19432;
  assign n19397 = ~n19433;
  assign n19395 = n19447 & n19448;
  assign n19381 = n19449 ^ n16963;
  assign n19435 = n19453 & n19454;
  assign n19436 = ~n19458;
  assign n19455 = n15799 & n19459;
  assign n18269 = ~n19460;
  assign n19462 = n19478 & n19479;
  assign n19411 = ~n19426;
  assign n19428 = n19381 & n19434;
  assign n19377 = n19435 ^ n19436;
  assign n19412 = ~n19395;
  assign n19427 = ~n19381;
  assign n19437 = ~n19435;
  assign n18246 = ~n19455;
  assign n15681 = n19461 ^ n19462;
  assign n19463 = ~n19462;
  assign n19407 = n19411 & n19412;
  assign n19394 = n19411 & n19397;
  assign n19415 = n19377 & n236;
  assign n19420 = n19427 & n19399;
  assign n19383 = ~n19428;
  assign n19413 = ~n19377;
  assign n19429 = n19437 & n19438;
  assign n19430 = n15681 & n18186;
  assign n19441 = n15681 & n19450;
  assign n15692 = ~n15681;
  assign n19456 = n19463 & n19464;
  assign n19375 = n19394 ^ n19395;
  assign n19396 = ~n19407;
  assign n19408 = n19413 & n19414;
  assign n19358 = ~n19415;
  assign n19401 = ~n19420;
  assign n19416 = ~n19429;
  assign n19363 = n19430 ^ n16928;
  assign n18230 = ~n19441;
  assign n19439 = n15692 & n19442;
  assign n19443 = ~n19456;
  assign n19171 = n19374 ^ n19375;
  assign n19332 = n19375 & n19374;
  assign n19376 = n19396 & n19397;
  assign n19379 = ~n19408;
  assign n19398 = n19416 & n19417;
  assign n19410 = n19363 & n19418;
  assign n19409 = ~n19363;
  assign n18214 = ~n19439;
  assign n19421 = n19443 & n19444;
  assign n17947 = ~n19171;
  assign n19356 = n19376 ^ n19377;
  assign n19378 = ~n19376;
  assign n19380 = n19398 ^ n19399;
  assign n19400 = ~n19398;
  assign n19402 = n19409 & n19339;
  assign n19365 = ~n19410;
  assign n18227 = n18230 & n18214;
  assign n19404 = n19421 ^ n16837;
  assign n19422 = ~n19421;
  assign n19333 = n236 ^ n19356;
  assign n19372 = n19378 & n19379;
  assign n19335 = n19380 ^ n19381;
  assign n19392 = n19400 & n19401;
  assign n19341 = ~n19402;
  assign n15656 = n19403 ^ n19404;
  assign n19419 = n19422 & n19423;
  assign n19105 = n19332 ^ n19333;
  assign n19293 = n19333 & n19332;
  assign n19361 = n19335 & n235;
  assign n19357 = ~n19372;
  assign n19359 = ~n19335;
  assign n19382 = ~n19392;
  assign n19386 = n15656 & n19393;
  assign n15591 = ~n15656;
  assign n19405 = ~n19419;
  assign n19116 = ~n19105;
  assign n19334 = n19357 & n19358;
  assign n19352 = n19359 & n19360;
  assign n19314 = ~n19361;
  assign n19362 = n19382 & n19383;
  assign n19367 = n15591 & n18077;
  assign n18177 = ~n19386;
  assign n19384 = n15591 & n19387;
  assign n19388 = n19405 & n19406;
  assign n19312 = n19334 ^ n19335;
  assign n19337 = ~n19334;
  assign n19336 = ~n19352;
  assign n19338 = n19362 ^ n19363;
  assign n19353 = n19367 ^ n16837;
  assign n19364 = ~n19362;
  assign n18197 = ~n19384;
  assign n15510 = n19388 ^ n19389;
  assign n19390 = ~n19388;
  assign n19294 = n235 ^ n19312;
  assign n19329 = n19336 & n19337;
  assign n19322 = n19338 ^ n19339;
  assign n19344 = n19353 & n19354;
  assign n19355 = n19364 & n19365;
  assign n19345 = ~n19353;
  assign n18194 = n18197 & n18177;
  assign n19368 = n15510 & n19373;
  assign n15600 = ~n15510;
  assign n19385 = n19390 & n19391;
  assign n19077 = n19293 ^ n19294;
  assign n19249 = n19294 & n19293;
  assign n19317 = n19322 & n234;
  assign n19313 = ~n19329;
  assign n19315 = ~n19322;
  assign n19300 = ~n19344;
  assign n19342 = n19345 & n19346;
  assign n19340 = ~n19355;
  assign n19347 = n15600 & n18112;
  assign n18143 = ~n19368;
  assign n19366 = n15600 & n19369;
  assign n19370 = ~n19385;
  assign n19069 = ~n19077;
  assign n19275 = n19313 & n19314;
  assign n19310 = n19315 & n19316;
  assign n19277 = ~n19317;
  assign n19297 = n19340 & n19341;
  assign n19319 = ~n19342;
  assign n19330 = n19347 ^ n16796;
  assign n18160 = ~n19366;
  assign n19348 = n19370 & n19371;
  assign n19295 = ~n19275;
  assign n19296 = ~n19310;
  assign n19320 = n19319 & n19300;
  assign n19318 = ~n19297;
  assign n19323 = n19330 & n19331;
  assign n19324 = ~n19330;
  assign n18157 = n18160 & n18143;
  assign n19326 = n19348 ^ n19349;
  assign n19350 = ~n19348;
  assign n19291 = n19295 & n19296;
  assign n19274 = n19296 & n19277;
  assign n19311 = n19318 & n19319;
  assign n19298 = ~n19320;
  assign n19258 = ~n19323;
  assign n19321 = n19324 & n19325;
  assign n15551 = n19326 ^ n16825;
  assign n19343 = n19350 & n19351;
  assign n19250 = n19274 ^ n19275;
  assign n19276 = ~n19291;
  assign n19231 = n19297 ^ n19298;
  assign n19299 = ~n19311;
  assign n19304 = n15551 & n18099;
  assign n19284 = ~n19321;
  assign n15543 = ~n15551;
  assign n19327 = ~n19343;
  assign n19038 = n19249 ^ n19250;
  assign n19213 = n19250 & n19249;
  assign n19251 = n19276 & n19277;
  assign n19280 = n19231 & n233;
  assign n19278 = ~n19231;
  assign n19281 = n19299 & n19300;
  assign n19301 = n19284 & n19258;
  assign n19286 = n15543 & n18055;
  assign n18102 = ~n19304;
  assign n19302 = n15543 & n19305;
  assign n19307 = n19327 & n19328;
  assign n19025 = ~n19038;
  assign n19230 = n233 ^ n19251;
  assign n19252 = ~n19251;
  assign n19270 = n19278 & n19279;
  assign n19233 = ~n19280;
  assign n19219 = n19286 ^ n16822;
  assign n19283 = ~n19281;
  assign n19282 = ~n19301;
  assign n18121 = ~n19302;
  assign n15440 = n19306 ^ n19307;
  assign n19308 = ~n19307;
  assign n19214 = n19230 ^ n19231;
  assign n19253 = ~n19270;
  assign n19265 = n19219 & n19271;
  assign n19193 = n19281 ^ n19282;
  assign n19272 = n19283 & n19284;
  assign n19264 = ~n19219;
  assign n19273 = n15440 & n18031;
  assign n19287 = n15440 & n19292;
  assign n15474 = ~n15440;
  assign n19303 = n19308 & n19309;
  assign n19015 = n19213 ^ n19214;
  assign n19172 = n19214 & n19213;
  assign n19244 = n19252 & n19253;
  assign n19256 = n19193 & n232;
  assign n19261 = n19264 & n19235;
  assign n19221 = ~n19265;
  assign n19254 = ~n19193;
  assign n19257 = ~n19272;
  assign n19259 = n19273 ^ n16777;
  assign n18086 = ~n19287;
  assign n19285 = n15474 & n19288;
  assign n19289 = ~n19303;
  assign n19004 = ~n19015;
  assign n19232 = ~n19244;
  assign n19245 = n19254 & n19255;
  assign n19195 = ~n19256;
  assign n19234 = n19257 & n19258;
  assign n19246 = n19259 & n19260;
  assign n19237 = ~n19261;
  assign n19247 = ~n19259;
  assign n18067 = ~n19285;
  assign n19267 = n19289 & n19290;
  assign n19215 = n19232 & n19233;
  assign n19218 = n19234 ^ n19235;
  assign n19217 = ~n19245;
  assign n19236 = ~n19234;
  assign n19182 = ~n19246;
  assign n19239 = n19247 & n19248;
  assign n19262 = n18086 & n18067;
  assign n15404 = n19266 ^ n19267;
  assign n19268 = ~n19267;
  assign n19192 = n232 ^ n19215;
  assign n19175 = n19218 ^ n19219;
  assign n19216 = ~n19215;
  assign n19228 = n19236 & n19237;
  assign n19202 = ~n19239;
  assign n19229 = n15404 & n17975;
  assign n19241 = n15404 & n18044;
  assign n18084 = ~n19262;
  assign n15452 = ~n15404;
  assign n19263 = n19268 & n19269;
  assign n19173 = n19192 ^ n19193;
  assign n19198 = n19175 & n247;
  assign n19196 = ~n19175;
  assign n19209 = n19216 & n19217;
  assign n19220 = ~n19228;
  assign n19223 = n19202 & n19182;
  assign n19158 = n19229 ^ n16723;
  assign n19238 = n15452 & n19240;
  assign n18046 = ~n19241;
  assign n19242 = ~n19263;
  assign n17716 = n19172 ^ n19173;
  assign n19136 = n19173 & n19172;
  assign n19190 = n19196 & n19197;
  assign n19156 = ~n19198;
  assign n19194 = ~n19209;
  assign n19199 = n19220 & n19221;
  assign n19212 = n19158 & n19143;
  assign n19200 = ~n19223;
  assign n19210 = ~n19158;
  assign n18029 = ~n19238;
  assign n19224 = n19242 & n19243;
  assign n18944 = ~n17716;
  assign n19139 = ~n19136;
  assign n19177 = ~n19190;
  assign n19174 = n19194 & n19195;
  assign n19184 = n19199 ^ n19200;
  assign n19201 = ~n19199;
  assign n19204 = n19210 & n19211;
  assign n19160 = ~n19212;
  assign n15392 = n19224 ^ n19225;
  assign n19226 = ~n19224;
  assign n19154 = n19174 ^ n19175;
  assign n19180 = n19184 & n246;
  assign n19176 = ~n19174;
  assign n19178 = ~n19184;
  assign n19191 = n19201 & n19202;
  assign n19145 = ~n19204;
  assign n19206 = n15392 & n18011;
  assign n15382 = ~n15392;
  assign n19222 = n19226 & n19227;
  assign n19137 = n247 ^ n19154;
  assign n19168 = n19176 & n19177;
  assign n19169 = n19178 & n19179;
  assign n19118 = ~n19180;
  assign n19181 = ~n19191;
  assign n19185 = n15382 & n17885;
  assign n19203 = n15382 & n19205;
  assign n17989 = ~n19206;
  assign n19207 = ~n19222;
  assign n17659 = n19136 ^ n19137;
  assign n19138 = ~n19137;
  assign n19155 = ~n19168;
  assign n19141 = ~n19169;
  assign n19157 = n19181 & n19182;
  assign n19099 = n19185 ^ n16673;
  assign n18013 = ~n19203;
  assign n19187 = n19207 & n19208;
  assign n18926 = ~n17659;
  assign n19110 = n19138 & n19139;
  assign n19131 = n19155 & n19156;
  assign n19151 = n19141 & n19118;
  assign n19142 = n19157 ^ n19158;
  assign n19159 = ~n19157;
  assign n19163 = n19099 & n19170;
  assign n19164 = ~n19099;
  assign n15370 = n19186 ^ n19187;
  assign n19188 = ~n19187;
  assign n19113 = ~n19110;
  assign n19095 = n19142 ^ n19143;
  assign n19140 = ~n19131;
  assign n19132 = ~n19151;
  assign n19152 = n19159 & n19160;
  assign n19101 = ~n19163;
  assign n19161 = n19164 & n19122;
  assign n19153 = n15370 & n17864;
  assign n19165 = n15370 & n19171;
  assign n15374 = ~n15370;
  assign n19183 = n19188 & n19189;
  assign n19119 = n19095 & n19125;
  assign n19111 = n19131 ^ n19132;
  assign n19120 = ~n19095;
  assign n19133 = n19140 & n19141;
  assign n19144 = ~n19152;
  assign n19085 = n19153 ^ n16641;
  assign n19124 = ~n19161;
  assign n17971 = ~n19165;
  assign n19162 = n15374 & n17947;
  assign n19166 = ~n19183;
  assign n18868 = n19110 ^ n19111;
  assign n19097 = ~n19119;
  assign n19114 = n19120 & n245;
  assign n19112 = ~n19111;
  assign n19117 = ~n19133;
  assign n19121 = n19144 & n19145;
  assign n19134 = n19085 & n19146;
  assign n19135 = ~n19085;
  assign n17950 = ~n19162;
  assign n19148 = n19166 & n19167;
  assign n18862 = ~n18868;
  assign n19058 = n19112 & n19113;
  assign n19080 = ~n19114;
  assign n19094 = n19117 & n19118;
  assign n19098 = n19121 ^ n19122;
  assign n19123 = ~n19121;
  assign n19087 = ~n19134;
  assign n19126 = n19135 & n19063;
  assign n19128 = n19148 ^ n16566;
  assign n19149 = ~n19148;
  assign n19078 = n19094 ^ n19095;
  assign n19088 = n19098 ^ n19099;
  assign n19068 = ~n19058;
  assign n19096 = ~n19094;
  assign n19115 = n19123 & n19124;
  assign n19065 = ~n19126;
  assign n15329 = n19127 ^ n19128;
  assign n19147 = n19149 & n19150;
  assign n19059 = n245 ^ n19078;
  assign n19083 = n19088 & n244;
  assign n19081 = ~n19088;
  assign n19093 = n19096 & n19097;
  assign n19100 = ~n19115;
  assign n19104 = n15329 & n19116;
  assign n15320 = ~n15329;
  assign n19129 = ~n19147;
  assign n17520 = n19058 ^ n19059;
  assign n19008 = n19059 & n19068;
  assign n19075 = n19081 & n19082;
  assign n19040 = ~n19083;
  assign n19079 = ~n19093;
  assign n19084 = n19100 & n19101;
  assign n19089 = n15320 & n17772;
  assign n17911 = ~n19104;
  assign n19102 = n15320 & n19105;
  assign n19106 = n19129 & n19130;
  assign n18843 = ~n17520;
  assign n19011 = ~n19008;
  assign n19061 = ~n19075;
  assign n19031 = n19079 & n19080;
  assign n19062 = n19084 ^ n19085;
  assign n19019 = n19089 ^ n16566;
  assign n19086 = ~n19084;
  assign n17933 = ~n19102;
  assign n19090 = n19106 ^ n19107;
  assign n19108 = ~n19106;
  assign n19056 = n19061 & n19040;
  assign n19050 = n19062 ^ n19063;
  assign n19060 = ~n19031;
  assign n19076 = n19086 & n19087;
  assign n17930 = n17933 & n17911;
  assign n15234 = n19090 ^ n16480;
  assign n19103 = n19108 & n19109;
  assign n19043 = n19050 & n243;
  assign n19032 = ~n19056;
  assign n19041 = ~n19050;
  assign n19055 = n19060 & n19061;
  assign n19064 = ~n19076;
  assign n19057 = n15234 & n17835;
  assign n19070 = n15234 & n19077;
  assign n15261 = ~n15234;
  assign n19091 = ~n19103;
  assign n19009 = n19031 ^ n19032;
  assign n19033 = n19041 & n19042;
  assign n18995 = ~n19043;
  assign n19039 = ~n19055;
  assign n19044 = n19057 ^ n16480;
  assign n19046 = n19064 & n19065;
  assign n19066 = n15261 & n19069;
  assign n17891 = ~n19070;
  assign n19071 = n19091 & n19092;
  assign n18763 = n19008 ^ n19009;
  assign n19010 = ~n19009;
  assign n19017 = ~n19033;
  assign n18988 = n19039 & n19040;
  assign n19034 = n19044 & n19045;
  assign n19018 = n19046 ^ n19047;
  assign n19049 = n19046 & n19051;
  assign n19035 = ~n19044;
  assign n19048 = ~n19046;
  assign n17870 = ~n19066;
  assign n19052 = n19071 ^ n19072;
  assign n19073 = ~n19071;
  assign n18770 = ~n18763;
  assign n18965 = n19010 & n19011;
  assign n19013 = n19017 & n18995;
  assign n18951 = n19018 ^ n19019;
  assign n19016 = ~n18988;
  assign n18959 = ~n19034;
  assign n19024 = n19035 & n19036;
  assign n19037 = n19048 & n19047;
  assign n19023 = ~n19049;
  assign n17888 = n17891 & n17870;
  assign n15195 = n19052 ^ n16384;
  assign n19067 = n19073 & n19074;
  assign n18972 = ~n18965;
  assign n18996 = n18951 & n19000;
  assign n18989 = ~n19013;
  assign n18997 = ~n18951;
  assign n19012 = n19016 & n19017;
  assign n19020 = n19023 & n19019;
  assign n18983 = ~n19024;
  assign n19002 = ~n19037;
  assign n19014 = n15195 & n17784;
  assign n19026 = n15195 & n19038;
  assign n15228 = ~n15195;
  assign n19053 = ~n19067;
  assign n18966 = n18988 ^ n18989;
  assign n18975 = ~n18996;
  assign n18990 = n18997 & n242;
  assign n18994 = ~n19012;
  assign n19003 = n18983 & n18959;
  assign n18941 = n19014 ^ n16396;
  assign n19001 = ~n19020;
  assign n19021 = n15228 & n19025;
  assign n17846 = ~n19026;
  assign n19028 = n19053 & n19054;
  assign n17365 = n18965 ^ n18966;
  assign n18931 = n18966 & n18972;
  assign n18953 = ~n18990;
  assign n18973 = n18994 & n18995;
  assign n18991 = n18941 & n18998;
  assign n18980 = n19001 & n19002;
  assign n18981 = ~n19003;
  assign n18992 = ~n18941;
  assign n17822 = ~n19021;
  assign n15160 = n19027 ^ n19028;
  assign n19029 = ~n19028;
  assign n17401 = ~n17365;
  assign n18934 = ~n18931;
  assign n18950 = n242 ^ n18973;
  assign n18968 = n18980 ^ n18981;
  assign n18974 = ~n18973;
  assign n18943 = ~n18991;
  assign n18984 = n18992 & n18920;
  assign n18982 = ~n18980;
  assign n17843 = n17846 & n17822;
  assign n18993 = n15160 & n17733;
  assign n19005 = n15160 & n19015;
  assign n15211 = ~n15160;
  assign n19022 = n19029 & n19030;
  assign n18932 = n18950 ^ n18951;
  assign n18957 = n18968 & n241;
  assign n18967 = n18974 & n18975;
  assign n18955 = ~n18968;
  assign n18976 = n18982 & n18983;
  assign n18924 = ~n18984;
  assign n18977 = n18993 ^ n16170;
  assign n18999 = n15211 & n19004;
  assign n17796 = ~n19005;
  assign n19006 = ~n19022;
  assign n18683 = n18931 ^ n18932;
  assign n18933 = ~n18932;
  assign n18954 = n18955 & n18956;
  assign n18915 = ~n18957;
  assign n18952 = ~n18967;
  assign n18958 = ~n18976;
  assign n18971 = n18977 & n18978;
  assign n18969 = ~n18977;
  assign n17768 = ~n18999;
  assign n18985 = n19006 & n19007;
  assign n18894 = n18933 & n18934;
  assign n18922 = n18952 & n18953;
  assign n18936 = ~n18954;
  assign n18940 = n18958 & n18959;
  assign n18960 = n18969 & n18970;
  assign n18879 = ~n18971;
  assign n17793 = n17796 & n17768;
  assign n18962 = n18985 ^ n16215;
  assign n18986 = ~n18985;
  assign n18897 = ~n18894;
  assign n18921 = n18936 & n18915;
  assign n18919 = n18940 ^ n18941;
  assign n18935 = ~n18922;
  assign n18942 = ~n18940;
  assign n18904 = ~n18960;
  assign n15112 = n18961 ^ n18962;
  assign n18979 = n18986 & n18987;
  assign n18910 = n18919 ^ n18920;
  assign n18895 = n18921 ^ n18922;
  assign n18929 = n18935 & n18936;
  assign n18937 = n18942 & n18943;
  assign n18901 = n18904 & n18879;
  assign n18930 = n15112 & n17517;
  assign n18945 = n15112 & n17716;
  assign n15148 = ~n15112;
  assign n18963 = ~n18979;
  assign n17854 = n18894 ^ n18895;
  assign n18900 = n18910 & n240;
  assign n18898 = ~n18910;
  assign n18896 = ~n18895;
  assign n18914 = ~n18929;
  assign n18916 = n18930 ^ n16215;
  assign n18923 = ~n18937;
  assign n18938 = n15148 & n18944;
  assign n17743 = ~n18945;
  assign n18946 = n18963 & n18964;
  assign n17824 = n17854 ^ n18873;
  assign n18745 = n17854 & n16779;
  assign n18829 = n18896 & n18897;
  assign n18891 = n18898 & n18899;
  assign n18857 = ~n18900;
  assign n18850 = n18914 & n18915;
  assign n18913 = n18916 & n18917;
  assign n18902 = n18923 & n18924;
  assign n18911 = ~n18916;
  assign n17718 = ~n18938;
  assign n15132 = n18946 ^ n18947;
  assign n18948 = ~n18946;
  assign n18847 = n17824 ^ n17799;
  assign n18874 = ~n18891;
  assign n18812 = n18901 ^ n18902;
  assign n18875 = ~n18850;
  assign n18905 = n18911 & n18912;
  assign n18842 = ~n18913;
  assign n18903 = ~n18902;
  assign n18925 = n15132 & n17659;
  assign n15130 = ~n15132;
  assign n18939 = n18948 & n18949;
  assign n18823 = n18847 & n17799;
  assign n14886 = ~n18847;
  assign n18869 = n18874 & n18875;
  assign n18870 = n18874 & n18857;
  assign n18876 = n18812 & n18888;
  assign n18877 = ~n18812;
  assign n18892 = n18903 & n18904;
  assign n18861 = ~n18905;
  assign n18906 = n15130 & n17586;
  assign n17661 = ~n18925;
  assign n18918 = n15130 & n18926;
  assign n18927 = ~n18939;
  assign n18802 = n18823 ^ n18824;
  assign n18797 = n18823 ^ n18825;
  assign n18856 = ~n18869;
  assign n18851 = ~n18870;
  assign n18837 = ~n18876;
  assign n18871 = n18877 & n255;
  assign n18880 = n18861 & n18842;
  assign n18878 = ~n18892;
  assign n18889 = n18906 ^ n16174;
  assign n17691 = ~n18918;
  assign n18907 = n18927 & n18928;
  assign n18131 = n455 ^ n18797;
  assign n18771 = n18802 & n18803;
  assign n18596 = n18797 & n455;
  assign n18830 = n18850 ^ n18851;
  assign n18835 = n18856 & n18857;
  assign n18814 = ~n18871;
  assign n18858 = n18878 & n18879;
  assign n18859 = ~n18880;
  assign n18881 = n18889 & n18890;
  assign n18882 = ~n18889;
  assign n18885 = n18907 ^ n16064;
  assign n18908 = ~n18907;
  assign n18675 = n18771 ^ n18772;
  assign n18775 = n18771 & n18772;
  assign n18140 = ~n18131;
  assign n18773 = ~n18771;
  assign n18810 = n18829 ^ n18830;
  assign n18779 = n18830 & n18829;
  assign n18811 = n255 ^ n18835;
  assign n18836 = ~n18835;
  assign n18848 = n18858 ^ n18859;
  assign n18860 = ~n18858;
  assign n18791 = ~n18881;
  assign n18872 = n18882 & n18883;
  assign n15027 = n18884 ^ n18885;
  assign n18893 = n18908 & n18909;
  assign n18768 = n18773 & n18774;
  assign n18661 = ~n18775;
  assign n18805 = n18810 & n16753;
  assign n18780 = n18811 ^ n18812;
  assign n18804 = ~n18810;
  assign n18782 = ~n18779;
  assign n18831 = n18836 & n18837;
  assign n18840 = n18848 & n254;
  assign n18838 = ~n18848;
  assign n18852 = n18860 & n18861;
  assign n18849 = n15027 & n17543;
  assign n18863 = n15027 & n18868;
  assign n18818 = ~n18872;
  assign n15088 = ~n15027;
  assign n18886 = ~n18893;
  assign n18684 = ~n18768;
  assign n18697 = n18779 ^ n18780;
  assign n18798 = n18804 & n16755;
  assign n18747 = ~n18805;
  assign n18781 = ~n18780;
  assign n18813 = ~n18831;
  assign n18832 = n18838 & n18839;
  assign n18756 = ~n18840;
  assign n18735 = n18849 ^ n16064;
  assign n18841 = ~n18852;
  assign n18853 = n18818 & n18791;
  assign n18854 = n15088 & n18862;
  assign n17634 = ~n18863;
  assign n18865 = n18886 & n18887;
  assign n18752 = n18697 & n16643;
  assign n18751 = ~n18697;
  assign n18753 = n18781 & n18782;
  assign n18776 = ~n18798;
  assign n18784 = n18813 & n18814;
  assign n18786 = ~n18832;
  assign n18827 = n18735 & n18833;
  assign n18815 = n18841 & n18842;
  assign n18826 = ~n18735;
  assign n18816 = ~n18853;
  assign n17600 = ~n18854;
  assign n14991 = n18864 ^ n18865;
  assign n18866 = ~n18865;
  assign n18743 = n18751 & n16590;
  assign n18725 = ~n18752;
  assign n18769 = n18776 & n18745;
  assign n18744 = n18776 & n18747;
  assign n18785 = ~n18784;
  assign n18783 = n18786 & n18756;
  assign n18731 = n18815 ^ n18816;
  assign n18819 = n18826 & n18758;
  assign n18737 = ~n18827;
  assign n18817 = ~n18815;
  assign n17631 = n17634 & n17600;
  assign n18828 = n14991 & n17272;
  assign n18844 = n14991 & n17520;
  assign n15044 = ~n14991;
  assign n18855 = n18866 & n18867;
  assign n18704 = ~n18743;
  assign n14864 = n18744 ^ n18745;
  assign n18746 = ~n18769;
  assign n18754 = n18783 ^ n18784;
  assign n18777 = n18785 & n18786;
  assign n18789 = n18731 & n253;
  assign n18787 = ~n18731;
  assign n18806 = n18817 & n18818;
  assign n18760 = ~n18819;
  assign n18807 = n18828 ^ n16004;
  assign n18834 = n15044 & n18843;
  assign n17560 = ~n18844;
  assign n18845 = ~n18855;
  assign n14866 = ~n14864;
  assign n18742 = n18746 & n18747;
  assign n18678 = n18753 ^ n18754;
  assign n18685 = n18754 & n18753;
  assign n18755 = ~n18777;
  assign n18778 = n18787 & n18788;
  assign n18710 = ~n18789;
  assign n18790 = ~n18806;
  assign n18799 = n18807 & n18808;
  assign n18800 = ~n18807;
  assign n17523 = ~n18834;
  assign n18820 = n18845 & n18846;
  assign n18702 = n14866 & n17679;
  assign n18729 = n18678 & n16532;
  assign n18724 = ~n18742;
  assign n18728 = ~n18678;
  assign n18688 = ~n18685;
  assign n18730 = n18755 & n18756;
  assign n18733 = ~n18778;
  assign n18757 = n18790 & n18791;
  assign n18696 = ~n18799;
  assign n18792 = n18800 & n18801;
  assign n18794 = n18820 ^ n15745;
  assign n18821 = ~n18820;
  assign n18674 = n18702 ^ n16755;
  assign n18698 = n18724 ^ n16590;
  assign n18723 = n18725 & n18724;
  assign n18726 = n18728 & n16539;
  assign n18680 = ~n18729;
  assign n18708 = n18730 ^ n18731;
  assign n18732 = ~n18730;
  assign n18734 = n18757 ^ n18758;
  assign n18759 = ~n18757;
  assign n18717 = ~n18792;
  assign n14928 = n18793 ^ n18794;
  assign n18809 = n18821 & n18822;
  assign n18659 = n18674 ^ n18675;
  assign n18676 = n18674 & n18684;
  assign n14796 = n18697 ^ n18698;
  assign n18686 = n253 ^ n18708;
  assign n18703 = ~n18723;
  assign n18655 = ~n18726;
  assign n18727 = n18732 & n18733;
  assign n18665 = n18734 ^ n18735;
  assign n18748 = n18759 & n18760;
  assign n18761 = n18717 & n18696;
  assign n18762 = n14928 & n18770;
  assign n14975 = ~n14928;
  assign n18795 = ~n18809;
  assign n18651 = n18659 & n454;
  assign n18649 = ~n18659;
  assign n18660 = ~n18676;
  assign n18653 = n14796 & n17625;
  assign n14799 = ~n14796;
  assign n18601 = n18685 ^ n18686;
  assign n18677 = n18703 & n18704;
  assign n18687 = ~n18686;
  assign n18713 = n18665 & n252;
  assign n18709 = ~n18727;
  assign n18711 = ~n18665;
  assign n18736 = ~n18748;
  assign n18715 = ~n18761;
  assign n18738 = n14975 & n17389;
  assign n17445 = ~n18762;
  assign n18749 = n14975 & n18763;
  assign n18764 = n18795 & n18796;
  assign n18646 = n18649 & n18650;
  assign n18600 = ~n18651;
  assign n18635 = n18653 ^ n16643;
  assign n18563 = n18660 & n18661;
  assign n18662 = n18601 & n16455;
  assign n18652 = n18677 ^ n18678;
  assign n18663 = ~n18601;
  assign n18637 = n18687 & n18688;
  assign n18679 = ~n18677;
  assign n18689 = n18709 & n18710;
  assign n18705 = n18711 & n18712;
  assign n18667 = ~n18713;
  assign n18714 = n18736 & n18737;
  assign n18643 = n18738 ^ n15745;
  assign n17485 = ~n18749;
  assign n18739 = n18764 ^ n18765;
  assign n18766 = ~n18764;
  assign n18626 = n18635 & n18636;
  assign n18625 = ~n18646;
  assign n18627 = ~n18635;
  assign n14766 = n18652 ^ n16539;
  assign n18598 = ~n18563;
  assign n18604 = ~n18662;
  assign n18656 = n18663 & n16441;
  assign n18672 = n18679 & n18680;
  assign n18664 = n252 ^ n18689;
  assign n18691 = ~n18689;
  assign n18690 = ~n18705;
  assign n18699 = n18714 ^ n18715;
  assign n18720 = n18643 & n18669;
  assign n18716 = ~n18714;
  assign n18718 = ~n18643;
  assign n17482 = n17485 & n17445;
  assign n14959 = n15838 ^ n18739;
  assign n18750 = n18766 & n18767;
  assign n18621 = n18625 & n18596;
  assign n18595 = n18625 & n18600;
  assign n18574 = ~n18626;
  assign n18622 = n18627 & n18628;
  assign n14762 = ~n14766;
  assign n18631 = ~n18656;
  assign n18638 = n18664 ^ n18665;
  assign n18654 = ~n18672;
  assign n18681 = n18690 & n18691;
  assign n18694 = n18699 & n251;
  assign n18692 = ~n18699;
  assign n18706 = n18716 & n18717;
  assign n18707 = n18718 & n18719;
  assign n18645 = ~n18720;
  assign n18700 = n14959 & n17277;
  assign n14913 = ~n14959;
  assign n18740 = ~n18750;
  assign n18569 = n18595 ^ n18596;
  assign n18599 = ~n18621;
  assign n18597 = ~n18622;
  assign n18594 = n14762 & n17459;
  assign n18576 = n18637 ^ n18638;
  assign n18629 = n18654 & n18655;
  assign n18639 = ~n18638;
  assign n18666 = ~n18681;
  assign n18682 = n18692 & n18693;
  assign n18613 = ~n18694;
  assign n18589 = n18700 ^ n15826;
  assign n18695 = ~n18706;
  assign n18671 = ~n18707;
  assign n18721 = n18740 & n18741;
  assign n16883 = n18569 ^ n18131;
  assign n18572 = ~n18569;
  assign n18551 = n18594 ^ n16539;
  assign n18591 = n18597 & n18598;
  assign n18493 = n18599 & n18600;
  assign n18592 = n18597 & n18574;
  assign n18611 = n18576 & n16390;
  assign n18602 = n18629 ^ n16441;
  assign n18610 = ~n18576;
  assign n18606 = n18639 & n18637;
  assign n18630 = ~n18629;
  assign n18632 = n18666 & n18667;
  assign n18641 = ~n18682;
  assign n18668 = n18695 & n18696;
  assign n14895 = n18721 ^ n18722;
  assign n18082 = ~n16883;
  assign n18466 = n18572 & n18140;
  assign n18571 = n18551 & n18582;
  assign n18570 = ~n18551;
  assign n18573 = ~n18591;
  assign n18516 = ~n18493;
  assign n18564 = ~n18592;
  assign n14694 = n18601 ^ n18602;
  assign n18605 = n18610 & n16402;
  assign n18578 = ~n18611;
  assign n18623 = n18630 & n18631;
  assign n18640 = ~n18632;
  assign n18657 = n18641 & n18613;
  assign n18642 = n18668 ^ n18669;
  assign n18670 = ~n18668;
  assign n18673 = n14895 & n18701;
  assign n15781 = ~n14895;
  assign n18548 = n18563 ^ n18564;
  assign n18562 = n18570 & n18520;
  assign n18546 = ~n18571;
  assign n18550 = n18573 & n18574;
  assign n14741 = ~n14694;
  assign n18554 = ~n18605;
  assign n18603 = ~n18623;
  assign n18634 = n18640 & n18641;
  assign n18585 = n18642 ^ n18643;
  assign n18633 = ~n18657;
  assign n18658 = n18670 & n18671;
  assign n18648 = n18673 ^ n15611;
  assign n17303 = n18683 ^ n15781;
  assign n18543 = n18548 & n453;
  assign n18519 = n18550 ^ n18551;
  assign n18541 = ~n18548;
  assign n18522 = ~n18562;
  assign n18547 = ~n18550;
  assign n18549 = n14741 & n17375;
  assign n18575 = n18603 & n18604;
  assign n18614 = n18585 & n18624;
  assign n18607 = n18632 ^ n18633;
  assign n18612 = ~n18634;
  assign n18615 = ~n18585;
  assign n18545 = n18647 ^ n18648;
  assign n18644 = ~n18658;
  assign n17289 = ~n17303;
  assign n18507 = n18519 ^ n18520;
  assign n18533 = n18541 & n18542;
  assign n18496 = ~n18543;
  assign n18540 = n18546 & n18547;
  assign n18531 = n18549 ^ n16441;
  assign n18552 = n18575 ^ n18576;
  assign n18577 = ~n18575;
  assign n18583 = n18606 ^ n18607;
  assign n18534 = n18607 & n18606;
  assign n18584 = n18612 & n18613;
  assign n18586 = ~n18614;
  assign n18608 = n18615 & n250;
  assign n18616 = n18644 & n18645;
  assign n18501 = n18507 & n452;
  assign n18499 = ~n18507;
  assign n18523 = n18531 & n18532;
  assign n18515 = ~n18533;
  assign n18521 = ~n18540;
  assign n18524 = ~n18531;
  assign n14704 = n16390 ^ n18552;
  assign n18565 = n18577 & n18578;
  assign n18580 = n18583 & n16178;
  assign n18556 = n18584 ^ n18585;
  assign n18579 = ~n18583;
  assign n18587 = ~n18584;
  assign n18558 = ~n18608;
  assign n18588 = n18616 ^ n18617;
  assign n18620 = n18616 & n18617;
  assign n18618 = ~n18616;
  assign n18490 = n18499 & n18500;
  assign n18448 = ~n18501;
  assign n18509 = n18515 & n18516;
  assign n18492 = n18515 & n18496;
  assign n18471 = n18521 & n18522;
  assign n18477 = ~n18523;
  assign n18517 = n18524 & n18525;
  assign n18508 = n14704 & n17295;
  assign n14707 = ~n14704;
  assign n18535 = n250 ^ n18556;
  assign n18553 = ~n18565;
  assign n18566 = n18579 & n16281;
  assign n18505 = ~n18580;
  assign n18581 = n18586 & n18587;
  assign n18537 = n18588 ^ n18589;
  assign n18609 = n18618 & n18619;
  assign n18593 = ~n18620;
  assign n18468 = ~n18490;
  assign n18467 = n18492 ^ n18493;
  assign n18436 = n18508 ^ n16390;
  assign n18495 = ~n18509;
  assign n18503 = ~n18471;
  assign n18502 = ~n18517;
  assign n18480 = n18534 ^ n18535;
  assign n18486 = n18535 & n18534;
  assign n18527 = n18553 & n18554;
  assign n18529 = ~n18566;
  assign n18561 = n18537 & n249;
  assign n18557 = ~n18581;
  assign n18559 = ~n18537;
  assign n18590 = n18593 & n18589;
  assign n18568 = ~n18609;
  assign n16849 = n18466 ^ n18467;
  assign n18470 = n18468 & n18448;
  assign n18425 = n18467 & n18466;
  assign n18483 = n18436 & n18491;
  assign n18445 = n18495 & n18496;
  assign n18494 = n18502 & n18503;
  assign n18497 = n18502 & n18477;
  assign n18484 = ~n18436;
  assign n18510 = n18480 & n16236;
  assign n18511 = ~n18480;
  assign n18498 = ~n18486;
  assign n18528 = ~n18527;
  assign n18526 = n18529 & n18505;
  assign n18536 = n18557 & n18558;
  assign n18555 = n18559 & n18560;
  assign n18514 = ~n18561;
  assign n18567 = ~n18590;
  assign n18073 = ~n16849;
  assign n18446 = ~n18470;
  assign n18434 = ~n18425;
  assign n18438 = ~n18483;
  assign n18478 = n18484 & n18454;
  assign n18469 = ~n18445;
  assign n18476 = ~n18494;
  assign n18472 = ~n18497;
  assign n18460 = ~n18510;
  assign n18506 = n18511 & n16224;
  assign n14666 = n18526 ^ n18527;
  assign n18518 = n18528 & n18529;
  assign n18512 = n18536 ^ n18537;
  assign n18539 = ~n18536;
  assign n18538 = ~n18555;
  assign n18544 = n18567 & n18568;
  assign n18426 = n18445 ^ n18446;
  assign n18461 = n18468 & n18469;
  assign n18428 = n18471 ^ n18472;
  assign n18453 = n18476 & n18477;
  assign n18456 = ~n18478;
  assign n18482 = ~n18506;
  assign n18485 = n14666 & n17216;
  assign n18487 = n249 ^ n18512;
  assign n14673 = ~n14666;
  assign n18504 = ~n18518;
  assign n18530 = n18538 & n18539;
  assign n18489 = n18544 ^ n18545;
  assign n16788 = n18425 ^ n18426;
  assign n18381 = n18426 & n18434;
  assign n18451 = n18428 & n451;
  assign n18435 = n18453 ^ n18454;
  assign n18447 = ~n18461;
  assign n18449 = ~n18428;
  assign n18455 = ~n18453;
  assign n18473 = n18485 ^ n16281;
  assign n18422 = n18486 ^ n18487;
  assign n18443 = n18487 & n18498;
  assign n18479 = n18504 & n18505;
  assign n18513 = ~n18530;
  assign n18008 = ~n16788;
  assign n18418 = n18435 ^ n18436;
  assign n18427 = n18447 & n18448;
  assign n18441 = n18449 & n18450;
  assign n18404 = ~n18451;
  assign n18452 = n18455 & n18456;
  assign n18462 = n18473 & n18474;
  assign n18463 = ~n18473;
  assign n18458 = n18479 ^ n18480;
  assign n18481 = ~n18479;
  assign n18488 = n18513 & n18514;
  assign n18411 = n18418 & n450;
  assign n18409 = ~n18418;
  assign n18401 = n18427 ^ n18428;
  assign n18430 = ~n18427;
  assign n18429 = ~n18441;
  assign n18437 = ~n18452;
  assign n14603 = n16236 ^ n18458;
  assign n18392 = ~n18462;
  assign n18457 = n18463 & n18464;
  assign n18475 = n18481 & n18482;
  assign n18465 = n18488 ^ n18489;
  assign n18382 = n451 ^ n18401;
  assign n18402 = n18409 & n18410;
  assign n18369 = ~n18411;
  assign n18419 = n18429 & n18430;
  assign n18412 = n18437 & n18438;
  assign n18420 = n14603 & n17175;
  assign n14654 = ~n14603;
  assign n18415 = ~n18457;
  assign n18444 = n248 ^ n18465;
  assign n18459 = ~n18475;
  assign n16730 = n18381 ^ n18382;
  assign n18383 = ~n18382;
  assign n18384 = ~n18402;
  assign n18403 = ~n18419;
  assign n18405 = n18420 ^ n16224;
  assign n18414 = ~n18412;
  assign n18439 = n18415 & n18392;
  assign n18431 = n18443 ^ n18444;
  assign n18442 = n18459 & n18460;
  assign n17968 = ~n16730;
  assign n18345 = n18383 & n18381;
  assign n18386 = n18384 & n18369;
  assign n18366 = n18403 & n18404;
  assign n18396 = n18405 & n18406;
  assign n18407 = n18414 & n18415;
  assign n18397 = ~n18405;
  assign n18424 = n18431 & n16058;
  assign n18413 = ~n18439;
  assign n18423 = ~n18431;
  assign n18440 = n18442 & n16110;
  assign n18432 = ~n18442;
  assign n18348 = ~n18345;
  assign n18367 = ~n18386;
  assign n18385 = ~n18366;
  assign n18358 = ~n18396;
  assign n18393 = n18397 & n18398;
  assign n18391 = ~n18407;
  assign n18395 = n18412 ^ n18413;
  assign n18417 = n18423 & n16045;
  assign n18365 = ~n18424;
  assign n18408 = n18432 ^ n18422;
  assign n18433 = n18432 & n16121;
  assign n18421 = ~n18440;
  assign n18346 = n18366 ^ n18367;
  assign n18378 = n18384 & n18385;
  assign n18355 = n18391 & n18392;
  assign n18372 = ~n18393;
  assign n18390 = n18395 & n449;
  assign n18388 = ~n18395;
  assign n14566 = n16110 ^ n18408;
  assign n18380 = ~n18417;
  assign n18416 = n18421 & n18422;
  assign n18400 = ~n18433;
  assign n17928 = n18345 ^ n18346;
  assign n18347 = ~n18346;
  assign n18368 = ~n18378;
  assign n18373 = n18372 & n18358;
  assign n18371 = ~n18355;
  assign n18387 = n18388 & n18389;
  assign n18330 = ~n18390;
  assign n18374 = n14566 & n17147;
  assign n14613 = ~n14566;
  assign n18394 = n18380 & n18365;
  assign n18399 = ~n18416;
  assign n17936 = ~n17928;
  assign n18325 = n18347 & n18348;
  assign n18350 = n18368 & n18369;
  assign n18370 = n18371 & n18372;
  assign n18356 = ~n18373;
  assign n18362 = n18374 ^ n16110;
  assign n18352 = ~n18387;
  assign n18376 = ~n18394;
  assign n18375 = n18399 & n18400;
  assign n18328 = ~n18325;
  assign n18342 = n18355 ^ n18356;
  assign n18351 = ~n18350;
  assign n18359 = n18362 & n18363;
  assign n18357 = ~n18370;
  assign n18360 = ~n18362;
  assign n18349 = n18352 & n18330;
  assign n14559 = n18375 ^ n18376;
  assign n18379 = ~n18375;
  assign n18336 = n18342 & n448;
  assign n18326 = n18349 ^ n18350;
  assign n18341 = n18351 & n18352;
  assign n18334 = ~n18342;
  assign n18310 = n18357 & n18358;
  assign n18316 = ~n18359;
  assign n18353 = n18360 & n18361;
  assign n14552 = ~n14559;
  assign n18377 = n18379 & n18380;
  assign n17909 = n18325 ^ n18326;
  assign n18331 = n18334 & n18335;
  assign n18290 = ~n18336;
  assign n18327 = ~n18326;
  assign n18329 = ~n18341;
  assign n18337 = ~n18310;
  assign n18338 = ~n18353;
  assign n18339 = n14552 & n17025;
  assign n18364 = ~n18377;
  assign n17915 = ~n17909;
  assign n18273 = n18327 & n18328;
  assign n18291 = n18329 & n18330;
  assign n18308 = ~n18331;
  assign n18332 = n18337 & n18338;
  assign n18333 = n18338 & n18316;
  assign n18321 = n18339 ^ n16045;
  assign n18354 = n18364 & n18365;
  assign n18309 = n18308 & n18290;
  assign n18280 = ~n18273;
  assign n18307 = ~n18291;
  assign n18317 = n18321 & n18322;
  assign n18315 = ~n18332;
  assign n18311 = ~n18333;
  assign n18318 = ~n18321;
  assign n18344 = n18354 & n15963;
  assign n18343 = ~n18354;
  assign n18306 = n18307 & n18308;
  assign n18292 = ~n18309;
  assign n18276 = n18310 ^ n18311;
  assign n18281 = n18315 & n18316;
  assign n18286 = ~n18317;
  assign n18312 = n18318 & n18319;
  assign n18340 = n18343 & n15973;
  assign n18324 = ~n18344;
  assign n18274 = n18291 ^ n18292;
  assign n18295 = n18276 & n463;
  assign n18289 = ~n18306;
  assign n18293 = ~n18276;
  assign n18302 = ~n18281;
  assign n18303 = ~n18312;
  assign n18323 = n18324 & n18304;
  assign n18314 = ~n18340;
  assign n17874 = n18273 ^ n18274;
  assign n18279 = ~n18274;
  assign n18275 = n18289 & n18290;
  assign n18287 = n18293 & n18294;
  assign n18261 = ~n18295;
  assign n18296 = n18302 & n18303;
  assign n18297 = n18303 & n18286;
  assign n18313 = ~n18323;
  assign n18320 = n18314 & n18324;
  assign n17867 = ~n17874;
  assign n18259 = n18275 ^ n18276;
  assign n18235 = n18279 & n18280;
  assign n18277 = ~n18275;
  assign n18278 = ~n18287;
  assign n18285 = ~n18296;
  assign n18282 = ~n18297;
  assign n18299 = n18313 & n18314;
  assign n18305 = ~n18320;
  assign n18236 = n463 ^ n18259;
  assign n18271 = n18277 & n18278;
  assign n18238 = n18281 ^ n18282;
  assign n18253 = n18285 & n18286;
  assign n14437 = n18298 ^ n18299;
  assign n14477 = n18304 ^ n18305;
  assign n18300 = ~n18299;
  assign n16481 = n18235 ^ n18236;
  assign n18207 = n18236 & n18235;
  assign n18265 = n18238 & n462;
  assign n18260 = ~n18271;
  assign n18262 = ~n18238;
  assign n18242 = ~n18253;
  assign n18270 = n14437 & n16950;
  assign n18272 = n14477 & n16979;
  assign n14498 = ~n14437;
  assign n18288 = n18300 & n18301;
  assign n14523 = ~n14477;
  assign n17820 = ~n16481;
  assign n18237 = n18260 & n18261;
  assign n18255 = n18262 & n18263;
  assign n18223 = ~n18265;
  assign n18251 = n18270 ^ n15756;
  assign n18254 = n18272 ^ n15973;
  assign n18283 = ~n18288;
  assign n18221 = n18237 ^ n18238;
  assign n18239 = ~n18237;
  assign n18249 = n18251 & n18252;
  assign n18232 = n18253 ^ n18254;
  assign n18240 = ~n18255;
  assign n18257 = n18254 & n18264;
  assign n18247 = ~n18251;
  assign n18256 = ~n18254;
  assign n18266 = n18283 & n18284;
  assign n18208 = n462 ^ n18221;
  assign n18224 = n18232 ^ n18233;
  assign n18231 = n18239 & n18240;
  assign n18243 = n18247 & n18248;
  assign n18193 = ~n18249;
  assign n18250 = n18256 & n18233;
  assign n18241 = ~n18257;
  assign n18244 = n18266 ^ n18267;
  assign n18268 = ~n18266;
  assign n17778 = n18207 ^ n18208;
  assign n18163 = n18208 & n18207;
  assign n18219 = n18224 & n461;
  assign n18217 = ~n18224;
  assign n18222 = ~n18231;
  assign n18234 = n18241 & n18242;
  assign n18212 = ~n18243;
  assign n14447 = n15787 ^ n18244;
  assign n18226 = ~n18250;
  assign n18258 = n18268 & n18269;
  assign n17765 = ~n17778;
  assign n18166 = ~n18163;
  assign n18215 = n18217 & n18218;
  assign n18184 = ~n18219;
  assign n18182 = n18222 & n18223;
  assign n18209 = n18212 & n18193;
  assign n18216 = n14447 & n16969;
  assign n18225 = ~n18234;
  assign n14454 = ~n14447;
  assign n18245 = ~n18258;
  assign n18204 = ~n18215;
  assign n18154 = n18216 ^ n15787;
  assign n18205 = ~n18182;
  assign n18210 = n18225 & n18226;
  assign n18228 = n18245 & n18246;
  assign n18198 = n18204 & n18205;
  assign n18181 = n18204 & n18184;
  assign n18202 = n18154 & n18174;
  assign n18200 = ~n18154;
  assign n18148 = n18209 ^ n18210;
  assign n18211 = ~n18210;
  assign n14393 = n18227 ^ n18228;
  assign n18229 = ~n18228;
  assign n18164 = n18181 ^ n18182;
  assign n18183 = ~n18198;
  assign n18189 = n18148 & n18199;
  assign n18190 = n18200 & n18201;
  assign n18156 = ~n18202;
  assign n18191 = ~n18148;
  assign n18206 = n18211 & n18212;
  assign n18203 = n14393 & n16928;
  assign n14340 = ~n14393;
  assign n18220 = n18229 & n18230;
  assign n16365 = n18163 ^ n18164;
  assign n18165 = ~n18164;
  assign n18167 = n18183 & n18184;
  assign n18168 = ~n18189;
  assign n18171 = ~n18190;
  assign n18187 = n18191 & n460;
  assign n18185 = n18203 ^ n15681;
  assign n18192 = ~n18206;
  assign n18213 = ~n18220;
  assign n17688 = ~n16365;
  assign n18126 = n18165 & n18166;
  assign n18147 = n460 ^ n18167;
  assign n18169 = ~n18167;
  assign n18180 = n18185 & n18186;
  assign n18150 = ~n18187;
  assign n18173 = n18192 & n18193;
  assign n18178 = ~n18185;
  assign n18195 = n18213 & n18214;
  assign n18127 = n18147 ^ n18148;
  assign n18161 = n18168 & n18169;
  assign n18153 = n18173 ^ n18174;
  assign n18175 = n18178 & n18179;
  assign n18118 = ~n18180;
  assign n18172 = ~n18173;
  assign n14319 = n18194 ^ n18195;
  assign n18196 = ~n18195;
  assign n17630 = n18126 ^ n18127;
  assign n18091 = n18127 & n18126;
  assign n18109 = n18153 ^ n18154;
  assign n18149 = ~n18161;
  assign n18170 = n18171 & n18172;
  assign n18138 = ~n18175;
  assign n18162 = n14319 & n16907;
  assign n14373 = ~n14319;
  assign n18188 = n18196 & n18197;
  assign n17644 = ~n17630;
  assign n18133 = n18109 & n18144;
  assign n18128 = n18149 & n18150;
  assign n18134 = ~n18109;
  assign n18135 = n18138 & n18118;
  assign n18095 = n18162 ^ n15656;
  assign n18155 = ~n18170;
  assign n18176 = ~n18188;
  assign n18108 = n459 ^ n18128;
  assign n18122 = ~n18133;
  assign n18129 = n18134 & n459;
  assign n18123 = ~n18128;
  assign n18146 = n18095 & n18151;
  assign n18136 = n18155 & n18156;
  assign n18145 = ~n18095;
  assign n18158 = n18176 & n18177;
  assign n18092 = n18108 ^ n18109;
  assign n18114 = n18122 & n18123;
  assign n18104 = ~n18129;
  assign n18088 = n18135 ^ n18136;
  assign n18139 = n18145 & n18077;
  assign n18097 = ~n18146;
  assign n18137 = ~n18136;
  assign n14282 = n18157 ^ n18158;
  assign n18159 = ~n18158;
  assign n17597 = n18091 ^ n18092;
  assign n18047 = n18092 & n18091;
  assign n18103 = ~n18114;
  assign n18115 = n18088 & n18124;
  assign n18116 = ~n18088;
  assign n18130 = n18137 & n18138;
  assign n18080 = ~n18139;
  assign n18125 = n14282 & n16874;
  assign n18141 = n14282 & n18131;
  assign n14337 = ~n14282;
  assign n18152 = n18159 & n18160;
  assign n17612 = ~n17597;
  assign n18050 = ~n18047;
  assign n18087 = n18103 & n18104;
  assign n18090 = ~n18115;
  assign n18110 = n18116 & n458;
  assign n18111 = n18125 ^ n15600;
  assign n18117 = ~n18130;
  assign n16919 = n18131 ^ n14337;
  assign n18132 = n14337 & n18140;
  assign n16921 = ~n18141;
  assign n18142 = ~n18152;
  assign n18068 = n18087 ^ n18088;
  assign n18089 = ~n18087;
  assign n18071 = ~n18110;
  assign n18107 = n18111 & n18112;
  assign n18094 = n18117 & n18118;
  assign n18105 = ~n18111;
  assign n16899 = ~n18132;
  assign n18119 = n18142 & n18143;
  assign n18048 = n458 ^ n18068;
  assign n18078 = n18089 & n18090;
  assign n18076 = n18094 ^ n18095;
  assign n18098 = n18105 & n18106;
  assign n18040 = ~n18107;
  assign n18096 = ~n18094;
  assign n18100 = n18119 ^ n15551;
  assign n18120 = ~n18119;
  assign n17495 = n18047 ^ n18048;
  assign n18049 = ~n18048;
  assign n18069 = n18076 ^ n18077;
  assign n18070 = ~n18078;
  assign n18093 = n18096 & n18097;
  assign n18064 = ~n18098;
  assign n14223 = n18099 ^ n18100;
  assign n18113 = n18120 & n18121;
  assign n17481 = ~n17495;
  assign n17996 = n18049 & n18050;
  assign n18060 = n18069 & n457;
  assign n18017 = n18070 & n18071;
  assign n18058 = ~n18069;
  assign n18061 = n18064 & n18040;
  assign n18072 = n14223 & n16825;
  assign n18081 = n14223 & n16883;
  assign n18079 = ~n18093;
  assign n14276 = ~n14223;
  assign n18101 = ~n18113;
  assign n17999 = ~n17996;
  assign n18054 = n18058 & n18059;
  assign n18019 = ~n18060;
  assign n18036 = ~n18017;
  assign n18005 = n18072 ^ n15543;
  assign n18062 = n18079 & n18080;
  assign n16885 = ~n18081;
  assign n18074 = n14276 & n18082;
  assign n18083 = n18101 & n18102;
  assign n18035 = ~n18054;
  assign n18052 = n18005 & n18055;
  assign n18001 = n18061 ^ n18062;
  assign n18053 = ~n18005;
  assign n18063 = ~n18062;
  assign n16869 = ~n18074;
  assign n14231 = n18083 ^ n18084;
  assign n18085 = ~n18083;
  assign n18032 = n18035 & n18036;
  assign n18016 = n18035 & n18019;
  assign n18037 = n18001 & n18051;
  assign n18007 = ~n18052;
  assign n18041 = n18053 & n18021;
  assign n18038 = ~n18001;
  assign n18056 = n18063 & n18064;
  assign n18065 = n14231 & n18073;
  assign n14227 = ~n14231;
  assign n18075 = n18085 & n18086;
  assign n17997 = n18016 ^ n18017;
  assign n18018 = ~n18032;
  assign n18003 = ~n18037;
  assign n18033 = n18038 & n456;
  assign n18022 = ~n18041;
  assign n18039 = ~n18056;
  assign n18042 = n14227 & n16668;
  assign n16835 = ~n18065;
  assign n18057 = n14227 & n16849;
  assign n18066 = ~n18075;
  assign n17442 = n17996 ^ n17997;
  assign n17998 = ~n17997;
  assign n18000 = n18018 & n18019;
  assign n17981 = ~n18033;
  assign n18020 = n18039 & n18040;
  assign n18030 = n18042 ^ n15440;
  assign n16851 = ~n18057;
  assign n18043 = n18066 & n18067;
  assign n17456 = ~n17442;
  assign n17960 = n17998 & n17999;
  assign n17979 = n18000 ^ n18001;
  assign n18002 = ~n18000;
  assign n18004 = n18020 ^ n18021;
  assign n18024 = n18030 & n18031;
  assign n18023 = ~n18020;
  assign n18025 = ~n18030;
  assign n18027 = n18043 ^ n18044;
  assign n18045 = ~n18043;
  assign n17961 = n456 ^ n17979;
  assign n17992 = n18002 & n18003;
  assign n17990 = n18004 ^ n18005;
  assign n18014 = n18022 & n18023;
  assign n17965 = ~n18024;
  assign n18015 = n18025 & n18026;
  assign n14153 = n15404 ^ n18027;
  assign n18034 = n18045 & n18046;
  assign n17322 = n17960 ^ n17961;
  assign n17912 = n17961 & n17960;
  assign n17984 = n17990 & n471;
  assign n17980 = ~n17992;
  assign n17982 = ~n17990;
  assign n17991 = n14153 & n16723;
  assign n18009 = n14153 & n16788;
  assign n18006 = ~n18014;
  assign n17986 = ~n18015;
  assign n14186 = ~n14153;
  assign n18028 = ~n18034;
  assign n17341 = ~n17322;
  assign n17937 = n17980 & n17981;
  assign n17974 = n17982 & n17983;
  assign n17942 = ~n17984;
  assign n17924 = n17991 ^ n15404;
  assign n17976 = n18006 & n18007;
  assign n17993 = n17986 & n17965;
  assign n17994 = n14186 & n18008;
  assign n16814 = ~n18009;
  assign n18010 = n18028 & n18029;
  assign n17962 = ~n17937;
  assign n17963 = ~n17974;
  assign n17972 = n17924 & n17975;
  assign n17973 = ~n17924;
  assign n17985 = ~n17976;
  assign n17977 = ~n17993;
  assign n16791 = ~n17994;
  assign n17987 = n18010 ^ n18011;
  assign n18012 = ~n18010;
  assign n17953 = n17962 & n17963;
  assign n17954 = n17963 & n17942;
  assign n17926 = ~n17972;
  assign n17966 = n17973 & n17944;
  assign n17897 = n17976 ^ n17977;
  assign n17978 = n17985 & n17986;
  assign n14172 = n15392 ^ n17987;
  assign n17995 = n18012 & n18013;
  assign n17941 = ~n17953;
  assign n17938 = ~n17954;
  assign n17957 = n17897 & n470;
  assign n17946 = ~n17966;
  assign n17955 = ~n17897;
  assign n17952 = n14172 & n16561;
  assign n17967 = n14172 & n16730;
  assign n17964 = ~n17978;
  assign n14095 = ~n14172;
  assign n17988 = ~n17995;
  assign n17916 = n17937 ^ n17938;
  assign n17920 = n17941 & n17942;
  assign n17904 = n17952 ^ n15392;
  assign n17951 = n17955 & n17956;
  assign n17899 = ~n17957;
  assign n17943 = n17964 & n17965;
  assign n16764 = ~n17967;
  assign n17958 = n14095 & n17968;
  assign n17969 = n17988 & n17989;
  assign n17211 = n17912 ^ n17916;
  assign n17879 = n17916 & n17912;
  assign n17896 = n470 ^ n17920;
  assign n17913 = ~n17916;
  assign n17921 = ~n17920;
  assign n17934 = n17904 & n17939;
  assign n17923 = n17943 ^ n17944;
  assign n17935 = ~n17904;
  assign n17922 = ~n17951;
  assign n17945 = ~n17943;
  assign n16733 = ~n17958;
  assign n17948 = n17969 ^ n15370;
  assign n17970 = ~n17969;
  assign n17880 = n17896 ^ n17897;
  assign n17228 = n17912 ^ n17913;
  assign n17917 = n17921 & n17922;
  assign n17914 = n17923 ^ n17924;
  assign n17906 = ~n17934;
  assign n17927 = n17935 & n17885;
  assign n17940 = n17945 & n17946;
  assign n14135 = n17947 ^ n17948;
  assign n17959 = n17970 & n17971;
  assign n16841 = n17879 ^ n17880;
  assign n17881 = ~n17880;
  assign n17902 = n17914 & n469;
  assign n17898 = ~n17917;
  assign n17900 = ~n17914;
  assign n17887 = ~n17927;
  assign n17929 = n14135 & n17936;
  assign n17925 = ~n17940;
  assign n14124 = ~n14135;
  assign n17949 = ~n17959;
  assign n16801 = n14886 ^ n16841;
  assign n16802 = n17854 ^ n16841;
  assign n17855 = ~n16841;
  assign n17830 = n17881 & n17879;
  assign n17849 = n17898 & n17899;
  assign n17893 = n17900 & n17901;
  assign n17857 = ~n17902;
  assign n17903 = n17925 & n17926;
  assign n17907 = n14124 & n16641;
  assign n17918 = n14124 & n17928;
  assign n16682 = ~n17929;
  assign n17931 = n17949 & n17950;
  assign n17823 = n16801 & n16779;
  assign n13785 = ~n16801;
  assign n17744 = n17855 & n14886;
  assign n17833 = ~n17830;
  assign n17883 = ~n17849;
  assign n17882 = ~n17893;
  assign n17884 = n17903 ^ n17904;
  assign n17841 = n17907 ^ n15370;
  assign n17905 = ~n17903;
  assign n16707 = ~n17918;
  assign n14018 = n17930 ^ n17931;
  assign n17932 = ~n17931;
  assign n17797 = n17823 ^ n17824;
  assign n17875 = n17882 & n17883;
  assign n17876 = n17882 & n17857;
  assign n17871 = n17884 ^ n17885;
  assign n17894 = n17905 & n17906;
  assign n16704 = n16707 & n16682;
  assign n17892 = n14018 & n16575;
  assign n17908 = n14018 & n17915;
  assign n14080 = ~n14018;
  assign n17919 = n17932 & n17933;
  assign n16609 = n167 ^ n17797;
  assign n17497 = n17797 & n167;
  assign n17798 = ~n17797;
  assign n17860 = n17871 & n468;
  assign n17856 = ~n17875;
  assign n17850 = ~n17876;
  assign n17858 = ~n17871;
  assign n17802 = n17892 ^ n15329;
  assign n17886 = ~n17894;
  assign n16654 = ~n17908;
  assign n17895 = n14080 & n17909;
  assign n17910 = ~n17919;
  assign n16617 = ~n16609;
  assign n17614 = n17798 & n17799;
  assign n17831 = n17849 ^ n17850;
  assign n17812 = n17856 & n17857;
  assign n17851 = n17858 & n17859;
  assign n17814 = ~n17860;
  assign n17872 = n17802 & n17877;
  assign n17861 = n17886 & n17887;
  assign n17873 = ~n17802;
  assign n16619 = ~n17895;
  assign n17889 = n17910 & n17911;
  assign n17810 = n17830 ^ n17831;
  assign n17832 = ~n17831;
  assign n17839 = ~n17812;
  assign n17838 = ~n17851;
  assign n17840 = n17861 ^ n17862;
  assign n17865 = n17861 & n17862;
  assign n17804 = ~n17872;
  assign n17866 = n17873 & n17772;
  assign n17863 = ~n17861;
  assign n16651 = n16654 & n16619;
  assign n14000 = n17888 ^ n17889;
  assign n17890 = ~n17889;
  assign n17807 = n17810 & n14866;
  assign n17806 = ~n17810;
  assign n17786 = n17832 & n17833;
  assign n17834 = n17838 & n17839;
  assign n17811 = n17838 & n17814;
  assign n17825 = n17840 ^ n17841;
  assign n17852 = n17863 & n17864;
  assign n17847 = ~n17865;
  assign n17774 = ~n17866;
  assign n17848 = n14000 & n16306;
  assign n17868 = n14000 & n17874;
  assign n14043 = ~n14000;
  assign n17878 = n17890 & n17891;
  assign n17800 = n17806 & n14864;
  assign n17780 = ~n17807;
  assign n17787 = n17811 ^ n17812;
  assign n17789 = ~n17786;
  assign n17817 = n17825 & n467;
  assign n17813 = ~n17834;
  assign n17815 = ~n17825;
  assign n17842 = n17847 & n17841;
  assign n17722 = n17848 ^ n15234;
  assign n17827 = ~n17852;
  assign n17853 = n14043 & n17867;
  assign n16588 = ~n17868;
  assign n17869 = ~n17878;
  assign n17779 = n17780 & n17744;
  assign n17769 = n17786 ^ n17787;
  assign n17759 = ~n17800;
  assign n17788 = ~n17787;
  assign n17755 = n17813 & n17814;
  assign n17808 = n17815 & n17816;
  assign n17763 = ~n17817;
  assign n17828 = n17722 & n17835;
  assign n17826 = ~n17842;
  assign n17829 = ~n17722;
  assign n16549 = ~n17853;
  assign n17844 = n17869 & n17870;
  assign n17761 = n17769 & n14799;
  assign n17758 = ~n17779;
  assign n17770 = n17759 & n17780;
  assign n17760 = ~n17769;
  assign n17729 = n17788 & n17789;
  assign n17790 = ~n17755;
  assign n17791 = ~n17808;
  assign n17801 = n17826 & n17827;
  assign n17724 = ~n17828;
  assign n17818 = n17829 & n17750;
  assign n17836 = n16588 & n16549;
  assign n13958 = n17843 ^ n17844;
  assign n17845 = ~n17844;
  assign n17703 = n17758 & n17759;
  assign n17754 = n17760 & n14796;
  assign n17709 = ~n17761;
  assign n17745 = ~n17770;
  assign n17732 = ~n17729;
  assign n17781 = n17790 & n17791;
  assign n17782 = n17791 & n17763;
  assign n17771 = n17801 ^ n17802;
  assign n17803 = ~n17801;
  assign n17752 = ~n17818;
  assign n17805 = n13958 & n16396;
  assign n17819 = n13958 & n16481;
  assign n16586 = ~n17836;
  assign n13994 = ~n13958;
  assign n17837 = n17845 & n17846;
  assign n13680 = n17744 ^ n17745;
  assign n17735 = ~n17703;
  assign n17736 = ~n17754;
  assign n17712 = n17771 ^ n17772;
  assign n17762 = ~n17781;
  assign n17756 = ~n17782;
  assign n17792 = n17803 & n17804;
  assign n17783 = n17805 ^ n15195;
  assign n16518 = ~n17819;
  assign n17809 = n13994 & n17820;
  assign n17821 = ~n17837;
  assign n17702 = n13680 & n16753;
  assign n17727 = n17735 & n17736;
  assign n17728 = n17736 & n17709;
  assign n13692 = ~n13680;
  assign n17748 = n17712 & n466;
  assign n17730 = n17755 ^ n17756;
  assign n17737 = n17762 & n17763;
  assign n17746 = ~n17712;
  assign n17777 = n17783 & n17784;
  assign n17773 = ~n17792;
  assign n17775 = ~n17783;
  assign n16484 = ~n17809;
  assign n17794 = n17821 & n17822;
  assign n17678 = n17702 ^ n14866;
  assign n17708 = ~n17727;
  assign n17704 = ~n17728;
  assign n17710 = n17729 ^ n17730;
  assign n17711 = n466 ^ n17737;
  assign n17738 = n17746 & n17747;
  assign n17694 = ~n17748;
  assign n17731 = ~n17730;
  assign n17720 = ~n17737;
  assign n17749 = n17773 & n17774;
  assign n17764 = n17775 & n17776;
  assign n17669 = ~n17777;
  assign n13946 = n17793 ^ n17794;
  assign n17795 = ~n17794;
  assign n17670 = n17678 & n17679;
  assign n17671 = ~n17678;
  assign n13626 = n17703 ^ n17704;
  assign n17649 = n17708 & n17709;
  assign n17705 = n17710 & n14762;
  assign n17681 = n17711 ^ n17712;
  assign n17706 = ~n17710;
  assign n17680 = n17731 & n17732;
  assign n17719 = ~n17738;
  assign n17721 = n17749 ^ n17750;
  assign n17751 = ~n17749;
  assign n17701 = ~n17764;
  assign n17753 = n13946 & n16355;
  assign n17766 = n13946 & n17778;
  assign n13953 = ~n13946;
  assign n17785 = n17795 & n17796;
  assign n17616 = ~n17670;
  assign n17662 = n17671 & n17672;
  assign n17582 = n17680 ^ n17681;
  assign n13619 = ~n13626;
  assign n17682 = ~n17649;
  assign n17674 = ~n17705;
  assign n17692 = n17706 & n14766;
  assign n17683 = ~n17681;
  assign n17713 = n17719 & n17720;
  assign n17684 = ~n17680;
  assign n17707 = n17721 ^ n17722;
  assign n17739 = n17751 & n17752;
  assign n17740 = n17701 & n17669;
  assign n17608 = n17753 ^ n15160;
  assign n17757 = n13953 & n17765;
  assign n16449 = ~n17766;
  assign n17767 = ~n17785;
  assign n17652 = n17582 & n14694;
  assign n17645 = ~n17662;
  assign n17646 = n13619 & n16590;
  assign n17651 = ~n17582;
  assign n17673 = n17674 & n17682;
  assign n17602 = n17683 & n17684;
  assign n17654 = ~n17692;
  assign n17697 = n17707 & n465;
  assign n17693 = ~n17713;
  assign n17695 = ~n17707;
  assign n17725 = n17608 & n17733;
  assign n17723 = ~n17739;
  assign n17699 = ~n17740;
  assign n17726 = ~n17608;
  assign n16409 = ~n17757;
  assign n17741 = n17767 & n17768;
  assign n17635 = n17645 & n17614;
  assign n17613 = n17616 & n17645;
  assign n17624 = n17646 ^ n14796;
  assign n17647 = n17651 & n14741;
  assign n17593 = ~n17652;
  assign n17653 = ~n17673;
  assign n17648 = n17654 & n17674;
  assign n17637 = n17693 & n17694;
  assign n17685 = n17695 & n17696;
  assign n17639 = ~n17697;
  assign n17698 = n17723 & n17724;
  assign n17610 = ~n17725;
  assign n17714 = n17726 & n17641;
  assign n16446 = n16449 & n16409;
  assign n17715 = n17741 ^ n15148;
  assign n17742 = ~n17741;
  assign n17590 = n17613 ^ n17614;
  assign n17617 = n17624 & n17625;
  assign n17615 = ~n17635;
  assign n17618 = ~n17624;
  assign n17626 = ~n17647;
  assign n13540 = n17648 ^ n17649;
  assign n17650 = n17653 & n17654;
  assign n17664 = ~n17637;
  assign n17663 = ~n17685;
  assign n17675 = n17698 ^ n17699;
  assign n17700 = ~n17698;
  assign n17643 = ~n17714;
  assign n13858 = n17715 ^ n17716;
  assign n17734 = n17742 & n17743;
  assign n17579 = n17590 & n166;
  assign n17577 = ~n17590;
  assign n17525 = n17615 & n17616;
  assign n17536 = ~n17617;
  assign n17601 = n17618 & n17619;
  assign n17591 = n13540 & n16539;
  assign n13571 = ~n13540;
  assign n17621 = ~n17650;
  assign n17655 = n17663 & n17664;
  assign n17636 = n17663 & n17639;
  assign n17667 = n17675 & n464;
  assign n17665 = ~n17675;
  assign n17686 = n17700 & n17701;
  assign n17687 = n13858 & n16365;
  assign n13910 = ~n13858;
  assign n17717 = ~n17734;
  assign n17561 = n17577 & n17578;
  assign n17499 = ~n17579;
  assign n17503 = n17591 ^ n14766;
  assign n17580 = ~n17525;
  assign n17581 = ~n17601;
  assign n17583 = n17621 ^ n14694;
  assign n17620 = n17621 & n17626;
  assign n17603 = n17636 ^ n17637;
  assign n17638 = ~n17655;
  assign n17656 = n17665 & n17666;
  assign n17568 = ~n17667;
  assign n17668 = ~n17686;
  assign n17657 = n13910 & n16231;
  assign n16326 = ~n17687;
  assign n17676 = n13910 & n17688;
  assign n17689 = n17717 & n17718;
  assign n17534 = ~n17561;
  assign n17546 = n17503 & n17562;
  assign n17563 = n17580 & n17581;
  assign n17564 = n17536 & n17581;
  assign n13534 = n17582 ^ n17583;
  assign n17547 = ~n17503;
  assign n17511 = n17602 ^ n17603;
  assign n17592 = ~n17620;
  assign n17604 = ~n17603;
  assign n17594 = n17638 & n17639;
  assign n17606 = ~n17656;
  assign n17541 = n17657 ^ n15112;
  assign n17640 = n17668 & n17669;
  assign n16367 = ~n17676;
  assign n17658 = n17689 ^ n15132;
  assign n17690 = ~n17689;
  assign n17524 = n17534 & n17497;
  assign n17496 = n17534 & n17499;
  assign n17504 = ~n17546;
  assign n17537 = n17547 & n17459;
  assign n17535 = ~n17563;
  assign n17526 = ~n17564;
  assign n13519 = ~n13534;
  assign n17565 = n17511 & n14704;
  assign n17548 = n17592 & n17593;
  assign n17566 = ~n17511;
  assign n17550 = n17604 & n17602;
  assign n17605 = ~n17594;
  assign n17627 = n17606 & n17568;
  assign n17607 = n17640 ^ n17641;
  assign n17642 = ~n17640;
  assign n13835 = n17658 ^ n17659;
  assign n17677 = n17690 & n17691;
  assign n17457 = n17496 ^ n17497;
  assign n17498 = ~n17524;
  assign n17500 = n17525 ^ n17526;
  assign n17502 = n17535 & n17536;
  assign n17501 = n13519 & n16455;
  assign n17464 = ~n17537;
  assign n17512 = n17548 ^ n14704;
  assign n17539 = ~n17565;
  assign n17549 = n17566 & n14707;
  assign n17538 = ~n17548;
  assign n17553 = ~n17550;
  assign n17596 = n17605 & n17606;
  assign n17584 = n17607 ^ n17608;
  assign n17595 = ~n17627;
  assign n17628 = n17642 & n17643;
  assign n17611 = n13835 & n16186;
  assign n17629 = n13835 & n17644;
  assign n13868 = ~n13835;
  assign n17660 = ~n17677;
  assign n15322 = n17457 ^ n16609;
  assign n17368 = n17457 & n16609;
  assign n17408 = n17498 & n17499;
  assign n17488 = n17500 & n165;
  assign n17413 = n17501 ^ n14741;
  assign n17458 = n17502 ^ n17503;
  assign n13486 = n17511 ^ n17512;
  assign n17486 = ~n17500;
  assign n17505 = ~n17502;
  assign n17527 = n17538 & n17539;
  assign n17507 = ~n17549;
  assign n17571 = n17584 & n479;
  assign n17551 = n17594 ^ n17595;
  assign n17567 = ~n17596;
  assign n17569 = ~n17584;
  assign n17585 = n17611 ^ n15130;
  assign n17609 = ~n17628;
  assign n16291 = ~n17629;
  assign n17622 = n13868 & n17630;
  assign n17632 = n17660 & n17661;
  assign n16547 = ~n15322;
  assign n17437 = n17458 ^ n17459;
  assign n17460 = n17413 & n17375;
  assign n17446 = n13486 & n16402;
  assign n17447 = ~n17408;
  assign n17475 = n17486 & n17487;
  assign n17411 = ~n17488;
  assign n17461 = ~n17413;
  assign n13496 = ~n13486;
  assign n17489 = n17504 & n17505;
  assign n17506 = ~n17527;
  assign n17424 = n17550 ^ n17551;
  assign n17491 = n17567 & n17568;
  assign n17554 = n17569 & n17570;
  assign n17493 = ~n17571;
  assign n17552 = ~n17551;
  assign n17572 = n17585 & n17586;
  assign n17573 = ~n17585;
  assign n17587 = n17609 & n17610;
  assign n16243 = ~n17622;
  assign n13839 = n17631 ^ n17632;
  assign n17633 = ~n17632;
  assign n17422 = n17437 & n164;
  assign n17336 = n17446 ^ n14704;
  assign n17420 = ~n17437;
  assign n17383 = ~n17460;
  assign n17449 = n17461 & n17462;
  assign n17448 = ~n17475;
  assign n17463 = ~n17489;
  assign n17465 = n17506 & n17507;
  assign n17513 = n17424 & n14666;
  assign n17514 = ~n17424;
  assign n17452 = n17552 & n17553;
  assign n17528 = ~n17491;
  assign n17529 = ~n17554;
  assign n17434 = ~n17572;
  assign n17557 = n17573 & n17574;
  assign n17575 = n17587 & n17588;
  assign n17555 = ~n17587;
  assign n16288 = n16291 & n16243;
  assign n17576 = n13839 & n16091;
  assign n17598 = n13839 & n17612;
  assign n13847 = ~n13839;
  assign n17623 = n17633 & n17634;
  assign n17403 = n17336 & n17295;
  assign n17406 = n17420 & n17421;
  assign n17331 = ~n17422;
  assign n17404 = ~n17336;
  assign n17438 = n17447 & n17448;
  assign n17407 = n17448 & n17411;
  assign n17423 = ~n17449;
  assign n17450 = n17463 & n17464;
  assign n17425 = n17465 ^ n14666;
  assign n17466 = ~n17465;
  assign n17467 = ~n17513;
  assign n17508 = n17514 & n14673;
  assign n17515 = n17528 & n17529;
  assign n17490 = n17529 & n17493;
  assign n17516 = n17555 ^ n17541;
  assign n17472 = ~n17557;
  assign n17556 = n17555 & n17517;
  assign n17540 = ~n17575;
  assign n17542 = n17576 ^ n15027;
  assign n17589 = n13847 & n17597;
  assign n16199 = ~n17598;
  assign n17599 = ~n17623;
  assign n17305 = ~n17403;
  assign n17392 = n17404 & n17405;
  assign n17370 = ~n17406;
  assign n17369 = n17407 ^ n17408;
  assign n13401 = n17424 ^ n17425;
  assign n17410 = ~n17438;
  assign n17412 = ~n17450;
  assign n17451 = n17466 & n17467;
  assign n17453 = n17490 ^ n17491;
  assign n17427 = ~n17508;
  assign n17492 = ~n17515;
  assign n17494 = n17516 ^ n17517;
  assign n17518 = n17472 & n17434;
  assign n17530 = n17540 & n17541;
  assign n17531 = n17542 & n17543;
  assign n17510 = ~n17556;
  assign n17532 = ~n17542;
  assign n16157 = ~n17589;
  assign n17558 = n17599 & n17600;
  assign n15278 = n17368 ^ n17369;
  assign n17372 = n17370 & n17331;
  assign n17344 = ~n17392;
  assign n17357 = n13401 & n16178;
  assign n17373 = ~n17369;
  assign n17327 = n17410 & n17411;
  assign n13458 = ~n13401;
  assign n17374 = n17412 ^ n17413;
  assign n17409 = n17423 & n17412;
  assign n17426 = ~n17451;
  assign n17428 = n17452 ^ n17453;
  assign n17359 = n17453 & n17452;
  assign n17395 = n17492 & n17493;
  assign n17478 = n17494 & n478;
  assign n17476 = ~n17494;
  assign n17470 = ~n17518;
  assign n17509 = ~n17530;
  assign n17355 = ~n17531;
  assign n17519 = n17532 & n17533;
  assign n17544 = n16199 & n16157;
  assign n17521 = n17558 ^ n14991;
  assign n17559 = ~n17558;
  assign n17240 = n17357 ^ n14666;
  assign n16444 = ~n15278;
  assign n17328 = ~n17372;
  assign n17290 = n17373 & n17368;
  assign n17345 = n17374 ^ n17375;
  assign n17371 = ~n17327;
  assign n17382 = ~n17409;
  assign n17338 = n17426 & n17427;
  assign n17414 = n17428 & n14603;
  assign n17415 = ~n17428;
  assign n17439 = ~n17395;
  assign n17468 = n17476 & n17477;
  assign n17397 = ~n17478;
  assign n17469 = n17509 & n17510;
  assign n17388 = ~n17519;
  assign n13792 = n17520 ^ n17521;
  assign n16197 = ~n17544;
  assign n17545 = n17559 & n17560;
  assign n17291 = n17327 ^ n17328;
  assign n17334 = n17345 & n163;
  assign n17293 = ~n17290;
  assign n17332 = ~n17345;
  assign n17358 = n17370 & n17371;
  assign n17376 = n17382 & n17383;
  assign n17384 = ~n17338;
  assign n17378 = ~n17414;
  assign n17393 = n17415 & n14654;
  assign n17440 = ~n17468;
  assign n17441 = n17469 ^ n17470;
  assign n17471 = ~n17469;
  assign n17479 = n17388 & n17355;
  assign n17455 = n13792 & n16015;
  assign n17480 = n13792 & n17495;
  assign n13803 = ~n13792;
  assign n17522 = ~n17545;
  assign n16429 = n17290 ^ n17291;
  assign n17292 = ~n17291;
  assign n17317 = n17332 & n17333;
  assign n17255 = ~n17334;
  assign n17330 = ~n17358;
  assign n17335 = ~n17376;
  assign n17377 = n17378 & n17384;
  assign n17347 = ~n17393;
  assign n17429 = n17439 & n17440;
  assign n17394 = n17440 & n17397;
  assign n17432 = n17441 & n477;
  assign n17430 = ~n17441;
  assign n17312 = n17455 ^ n15044;
  assign n17454 = n17471 & n17472;
  assign n17386 = ~n17479;
  assign n16118 = ~n17480;
  assign n17473 = n13803 & n17481;
  assign n17483 = n17522 & n17523;
  assign n16406 = ~n16429;
  assign n17213 = n17292 & n17293;
  assign n17296 = ~n17317;
  assign n17253 = n17330 & n17331;
  assign n17294 = n17335 ^ n17336;
  assign n17329 = n17335 & n17344;
  assign n17346 = ~n17377;
  assign n17337 = n17378 & n17347;
  assign n17360 = n17394 ^ n17395;
  assign n17396 = ~n17429;
  assign n17416 = n17430 & n17431;
  assign n17321 = ~n17432;
  assign n17417 = n17312 & n17435;
  assign n17418 = ~n17312;
  assign n17433 = ~n17454;
  assign n16069 = ~n17473;
  assign n13664 = n17482 ^ n17483;
  assign n17484 = ~n17483;
  assign n17265 = n17294 ^ n17295;
  assign n17252 = n17296 & n17255;
  assign n17297 = ~n17253;
  assign n17304 = ~n17329;
  assign n13391 = n17337 ^ n17338;
  assign n17230 = n17346 & n17347;
  assign n17339 = n17359 ^ n17360;
  assign n17307 = n17360 & n17359;
  assign n17349 = n17396 & n17397;
  assign n17362 = ~n17416;
  assign n17314 = ~n17417;
  assign n17398 = n17418 & n17272;
  assign n17385 = n17433 & n17434;
  assign n16115 = n16118 & n16069;
  assign n17419 = n13664 & n15913;
  assign n17443 = n13664 & n17456;
  assign n13729 = ~n13664;
  assign n17474 = n17484 & n17485;
  assign n17214 = n17252 ^ n17253;
  assign n17250 = n17265 & n162;
  assign n17248 = ~n17265;
  assign n17281 = n17296 & n17297;
  assign n17279 = n17304 & n17305;
  assign n17267 = n13391 & n16236;
  assign n13397 = ~n13391;
  assign n17298 = ~n17230;
  assign n17319 = n17339 & n14566;
  assign n17318 = ~n17339;
  assign n17310 = ~n17307;
  assign n17361 = ~n17349;
  assign n17348 = n17362 & n17321;
  assign n17363 = n17385 ^ n17386;
  assign n17275 = ~n17398;
  assign n17387 = ~n17385;
  assign n17201 = n17419 ^ n14975;
  assign n17436 = n13729 & n17442;
  assign n16025 = ~n17443;
  assign n17444 = ~n17474;
  assign n16309 = n17213 ^ n17214;
  assign n17150 = n17214 & n17213;
  assign n17241 = n17248 & n17249;
  assign n17187 = ~n17250;
  assign n17155 = n17267 ^ n14603;
  assign n17266 = n17279 & n17280;
  assign n17254 = ~n17281;
  assign n17251 = ~n17279;
  assign n17306 = n17318 & n14613;
  assign n17283 = ~n17319;
  assign n17308 = n17348 ^ n17349;
  assign n17350 = n17361 & n17362;
  assign n17353 = n17363 & n476;
  assign n17351 = ~n17363;
  assign n17379 = n17387 & n17388;
  assign n17381 = n17201 & n17389;
  assign n17380 = ~n17201;
  assign n15979 = ~n17436;
  assign n17399 = n17444 & n17445;
  assign n15200 = ~n16309;
  assign n17217 = ~n17241;
  assign n17215 = n17251 ^ n17240;
  assign n17185 = n17254 & n17255;
  assign n17256 = n17251 & n17216;
  assign n17239 = ~n17266;
  assign n17282 = n17283 & n17298;
  assign n17258 = ~n17306;
  assign n17284 = n17307 ^ n17308;
  assign n17309 = ~n17308;
  assign n17320 = ~n17350;
  assign n17340 = n17351 & n17352;
  assign n17244 = ~n17353;
  assign n17354 = ~n17379;
  assign n17364 = n17380 & n17236;
  assign n17204 = ~n17381;
  assign n17390 = n16025 & n15979;
  assign n17366 = n17399 ^ n14959;
  assign n17402 = n17399 & n17365;
  assign n17400 = ~n17399;
  assign n17195 = n17215 ^ n17216;
  assign n17184 = n17217 & n17187;
  assign n17229 = n17239 & n17240;
  assign n17218 = ~n17185;
  assign n17207 = ~n17256;
  assign n17257 = ~n17282;
  assign n17268 = n17258 & n17283;
  assign n17269 = n17284 & n14559;
  assign n17270 = ~n17284;
  assign n17221 = n17309 & n17310;
  assign n17260 = n17320 & n17321;
  assign n17286 = ~n17340;
  assign n17311 = n17354 & n17355;
  assign n17238 = ~n17364;
  assign n13677 = n17365 ^ n17366;
  assign n16023 = ~n17390;
  assign n17391 = n17400 & n17401;
  assign n17326 = ~n17402;
  assign n17151 = n17184 ^ n17185;
  assign n17183 = n17195 & n161;
  assign n17181 = ~n17195;
  assign n17208 = n17217 & n17218;
  assign n17206 = ~n17229;
  assign n17197 = n17257 & n17258;
  assign n17231 = ~n17268;
  assign n17190 = ~n17269;
  assign n17259 = n17270 & n14552;
  assign n17224 = ~n17221;
  assign n17285 = ~n17260;
  assign n17299 = n17286 & n17244;
  assign n17271 = n17311 ^ n17312;
  assign n17313 = ~n17311;
  assign n17301 = n13677 & n15838;
  assign n17323 = n13677 & n17341;
  assign n13689 = ~n13677;
  assign n17367 = n17326 & n14913;
  assign n17343 = ~n17391;
  assign n16265 = n17150 ^ n17151;
  assign n17089 = n17151 & n17150;
  assign n17174 = n17181 & n17182;
  assign n17118 = ~n17183;
  assign n17188 = n17206 & n17207;
  assign n17186 = ~n17208;
  assign n13360 = n17230 ^ n17231;
  assign n17219 = ~n17197;
  assign n17220 = ~n17259;
  assign n17242 = n17271 ^ n17272;
  assign n17273 = n17285 & n17286;
  assign n17261 = ~n17299;
  assign n17276 = n17301 ^ n14959;
  assign n17300 = n17313 & n17314;
  assign n17315 = n13689 & n17322;
  assign n15916 = ~n17323;
  assign n17356 = n17343 & n14959;
  assign n17342 = ~n17367;
  assign n16241 = ~n16265;
  assign n17092 = ~n17089;
  assign n17152 = ~n17174;
  assign n17116 = n17186 & n17187;
  assign n17176 = n17188 & n17131;
  assign n17160 = ~n17188;
  assign n17209 = n17219 & n17220;
  assign n13349 = ~n13360;
  assign n17196 = n17220 & n17190;
  assign n17234 = n17242 & n475;
  assign n17232 = ~n17242;
  assign n17222 = n17260 ^ n17261;
  assign n17243 = ~n17273;
  assign n17262 = n17276 & n17277;
  assign n17263 = ~n17276;
  assign n17274 = ~n17300;
  assign n15893 = ~n17315;
  assign n17324 = n17342 & n17343;
  assign n17325 = ~n17356;
  assign n17115 = n17152 & n17118;
  assign n17130 = n17160 ^ n17155;
  assign n17153 = ~n17116;
  assign n17161 = n17160 & n17175;
  assign n17154 = ~n17176;
  assign n17162 = n13349 & n16121;
  assign n13296 = n17196 ^ n17197;
  assign n17189 = ~n17209;
  assign n17198 = n17221 ^ n17222;
  assign n17225 = n17232 & n17233;
  assign n17166 = ~n17234;
  assign n17164 = n17243 & n17244;
  assign n17223 = ~n17222;
  assign n17144 = ~n17262;
  assign n17245 = n17263 & n17264;
  assign n17235 = n17274 & n17275;
  assign n15931 = n15916 & n15893;
  assign n17302 = ~n17324;
  assign n17316 = n17325 & n17326;
  assign n17090 = n17115 ^ n17116;
  assign n17064 = n17130 ^ n17131;
  assign n17145 = n17152 & n17153;
  assign n17146 = n17154 & n17155;
  assign n17120 = ~n17161;
  assign n17066 = n17162 ^ n14566;
  assign n17148 = n13296 & n16058;
  assign n17126 = n17189 & n17190;
  assign n13327 = ~n13296;
  assign n17192 = n17198 & n14477;
  assign n17191 = ~n17198;
  assign n17134 = n17223 & n17224;
  assign n17199 = ~n17225;
  assign n17200 = ~n17164;
  assign n17202 = n17235 ^ n17236;
  assign n17173 = ~n17245;
  assign n17237 = ~n17235;
  assign n17287 = n17302 & n17303;
  assign n17288 = ~n17316;
  assign n16176 = n17089 ^ n17090;
  assign n17102 = n17064 & n17111;
  assign n17091 = ~n17090;
  assign n17103 = ~n17064;
  assign n17117 = ~n17145;
  assign n17119 = ~n17146;
  assign n17133 = n17066 & n17147;
  assign n17047 = n17148 ^ n14559;
  assign n17132 = ~n17066;
  assign n17157 = ~n17126;
  assign n17177 = n17191 & n14523;
  assign n17156 = ~n17192;
  assign n17193 = n17199 & n17200;
  assign n17163 = n17199 & n17166;
  assign n17178 = n17201 ^ n17202;
  assign n17137 = ~n17134;
  assign n17210 = n17173 & n17144;
  assign n17226 = n17237 & n17238;
  assign n17247 = ~n17287;
  assign n17278 = n17288 & n17289;
  assign n16155 = ~n16176;
  assign n17041 = n17091 & n17092;
  assign n17086 = ~n17102;
  assign n17094 = n17103 & n160;
  assign n17093 = n17117 & n17118;
  assign n17095 = n17119 & n17120;
  assign n17112 = n17047 & n17121;
  assign n17122 = n17132 & n17096;
  assign n17068 = ~n17133;
  assign n17113 = ~n17047;
  assign n17149 = n17156 & n17157;
  assign n17135 = n17163 ^ n17164;
  assign n17124 = ~n17177;
  assign n17169 = n17178 & n474;
  assign n17165 = ~n17193;
  assign n17167 = ~n17178;
  assign n17171 = ~n17210;
  assign n17203 = ~n17226;
  assign n17246 = ~n17278;
  assign n17063 = n160 ^ n17093;
  assign n17062 = ~n17094;
  assign n17065 = n17095 ^ n17096;
  assign n17087 = ~n17093;
  assign n17097 = ~n17095;
  assign n17049 = ~n17112;
  assign n17104 = n17113 & n17025;
  assign n17098 = ~n17122;
  assign n17114 = n17134 ^ n17135;
  assign n17123 = ~n17149;
  assign n17125 = n17124 & n17156;
  assign n17136 = ~n17135;
  assign n17100 = n17165 & n17166;
  assign n17158 = n17167 & n17168;
  assign n17108 = ~n17169;
  assign n17170 = n17203 & n17204;
  assign n13557 = n17246 & n17247;
  assign n17042 = n17063 ^ n17064;
  assign n17054 = n17065 ^ n17066;
  assign n17076 = n17086 & n17087;
  assign n17088 = n17097 & n17098;
  assign n17027 = ~n17104;
  assign n17105 = n17114 & n14498;
  assign n17050 = n17123 & n17124;
  assign n13235 = n17125 ^ n17126;
  assign n17106 = ~n17114;
  assign n17071 = n17136 & n17137;
  assign n17138 = ~n17100;
  assign n17139 = ~n17158;
  assign n17081 = n17170 ^ n17171;
  assign n17172 = ~n17170;
  assign n17194 = n13557 & n17227;
  assign n17212 = n13557 & n17228;
  assign n14935 = ~n13557;
  assign n16067 = n17041 ^ n17042;
  assign n16981 = n17042 & n17041;
  assign n17045 = n17054 & n175;
  assign n17043 = ~n17054;
  assign n17061 = ~n17076;
  assign n17067 = ~n17088;
  assign n17077 = n13235 & n15973;
  assign n17056 = ~n17105;
  assign n17099 = n17106 & n14437;
  assign n17078 = ~n17050;
  assign n13303 = ~n13235;
  assign n17074 = ~n17071;
  assign n17127 = n17138 & n17139;
  assign n17128 = n17139 & n17108;
  assign n17142 = n17081 & n473;
  assign n17140 = ~n17081;
  assign n17159 = n17172 & n17173;
  assign n17085 = n17194 ^ n14895;
  assign n17205 = n14935 & n17211;
  assign n17180 = ~n17212;
  assign n16092 = ~n16067;
  assign n17038 = n17043 & n17044;
  assign n17002 = ~n17045;
  assign n17000 = n17061 & n17062;
  assign n17046 = n17067 & n17068;
  assign n16991 = n17077 ^ n14477;
  assign n17079 = ~n17099;
  assign n17107 = ~n17127;
  assign n17101 = ~n17128;
  assign n17129 = n17140 & n17141;
  assign n17060 = ~n17142;
  assign n17143 = ~n17159;
  assign n17179 = ~n17205;
  assign n17022 = ~n17038;
  assign n17024 = n17046 ^ n17047;
  assign n17023 = ~n17000;
  assign n17048 = ~n17046;
  assign n17069 = n17078 & n17079;
  assign n17070 = n17079 & n17056;
  assign n17072 = n17100 ^ n17101;
  assign n17080 = n17107 & n17108;
  assign n17083 = ~n17129;
  assign n17109 = n17143 & n17144;
  assign n15866 = n17179 & n17180;
  assign n17021 = n17022 & n17023;
  assign n16999 = n17022 & n17002;
  assign n17010 = n17024 ^ n17025;
  assign n17039 = n17048 & n17049;
  assign n17055 = ~n17069;
  assign n17051 = ~n17070;
  assign n17013 = n17071 ^ n17072;
  assign n17057 = n17080 ^ n17081;
  assign n17073 = ~n17072;
  assign n17082 = ~n17080;
  assign n17084 = n17109 ^ n17110;
  assign n15848 = ~n15866;
  assign n16982 = n16999 ^ n17000;
  assign n17005 = n17010 & n174;
  assign n17001 = ~n17021;
  assign n17003 = ~n17010;
  assign n17026 = ~n17039;
  assign n13277 = n17050 ^ n17051;
  assign n17031 = n17055 & n17056;
  assign n17053 = n17013 & n14447;
  assign n17030 = n473 ^ n17057;
  assign n17052 = ~n17013;
  assign n17029 = n17073 & n17074;
  assign n17075 = n17082 & n17083;
  assign n17058 = n17084 ^ n17085;
  assign n15051 = n16981 ^ n16982;
  assign n16983 = ~n16982;
  assign n16957 = n17001 & n17002;
  assign n16995 = n17003 & n17004;
  assign n16966 = ~n17005;
  assign n17011 = n17026 & n17027;
  assign n16970 = n17029 ^ n17030;
  assign n17014 = n17031 ^ n14447;
  assign n13268 = ~n13277;
  assign n17033 = ~n17031;
  assign n17040 = n17052 & n14454;
  assign n17032 = ~n17053;
  assign n17034 = ~n17030;
  assign n17037 = n472 ^ n17058;
  assign n17035 = ~n17029;
  assign n17059 = ~n17075;
  assign n16005 = ~n15051;
  assign n16939 = n16983 & n16981;
  assign n16984 = ~n16957;
  assign n16985 = ~n16995;
  assign n17006 = n17011 & n17012;
  assign n13233 = n17013 ^ n17014;
  assign n16996 = ~n17011;
  assign n17016 = n16970 & n14340;
  assign n17007 = n13268 & n15874;
  assign n17015 = ~n16970;
  assign n17028 = n17032 & n17033;
  assign n17017 = n17034 & n17035;
  assign n17020 = ~n17040;
  assign n17036 = n17059 & n17060;
  assign n16976 = n16984 & n16985;
  assign n16977 = n16985 & n16966;
  assign n16978 = n16996 ^ n16991;
  assign n16980 = n13233 & n15799;
  assign n16997 = n16996 & n16979;
  assign n16990 = ~n17006;
  assign n13239 = ~n13233;
  assign n16931 = n17007 ^ n14437;
  assign n17008 = n17015 & n14393;
  assign n16975 = ~n17016;
  assign n17019 = ~n17028;
  assign n17018 = n17036 ^ n17037;
  assign n16965 = ~n16976;
  assign n16958 = ~n16977;
  assign n16967 = n16978 ^ n16979;
  assign n16968 = n16980 ^ n14447;
  assign n16986 = n16990 & n16991;
  assign n16973 = ~n16997;
  assign n16992 = ~n17008;
  assign n16998 = n17017 ^ n17018;
  assign n17009 = n17019 & n17020;
  assign n16940 = n16957 ^ n16958;
  assign n16913 = n16965 & n16966;
  assign n16961 = n16967 & n173;
  assign n16964 = n16968 & n16969;
  assign n16959 = ~n16967;
  assign n16962 = ~n16968;
  assign n16972 = ~n16986;
  assign n16994 = n16998 & n14373;
  assign n16993 = ~n16998;
  assign n16989 = ~n17009;
  assign n15890 = n16939 ^ n16940;
  assign n15765 = n16940 & n16939;
  assign n16941 = ~n16913;
  assign n16946 = n16959 & n16960;
  assign n16924 = ~n16961;
  assign n16952 = n16962 & n16963;
  assign n16890 = ~n16964;
  assign n16947 = n16972 & n16973;
  assign n16971 = n16989 ^ n14393;
  assign n16987 = n16989 & n16992;
  assign n16988 = n16993 & n14319;
  assign n16938 = ~n16994;
  assign n15914 = ~n15890;
  assign n16942 = ~n16946;
  assign n16930 = n16947 ^ n16948;
  assign n16903 = ~n16952;
  assign n16951 = n16947 & n16948;
  assign n16949 = ~n16947;
  assign n13139 = n16970 ^ n16971;
  assign n16974 = ~n16987;
  assign n16956 = ~n16988;
  assign n16922 = n16930 ^ n16931;
  assign n16932 = n16941 & n16942;
  assign n16933 = n16942 & n16924;
  assign n16935 = n16890 & n16903;
  assign n16944 = n16949 & n16950;
  assign n16943 = ~n16951;
  assign n16936 = n13139 & n15692;
  assign n13178 = ~n13139;
  assign n16954 = n16974 & n16975;
  assign n16953 = n16956 & n16938;
  assign n16912 = n16922 & n172;
  assign n16910 = ~n16922;
  assign n16923 = ~n16932;
  assign n16914 = ~n16933;
  assign n16901 = ~n16935;
  assign n16927 = n16936 ^ n14393;
  assign n16934 = n16943 & n16931;
  assign n16926 = ~n16944;
  assign n13152 = n16953 ^ n16954;
  assign n16955 = ~n16954;
  assign n16906 = n16910 & n16911;
  assign n16879 = ~n16912;
  assign n15731 = n16913 ^ n16914;
  assign n16875 = n16923 & n16924;
  assign n16915 = n16927 & n16928;
  assign n16916 = ~n16927;
  assign n16925 = ~n16934;
  assign n16929 = n13152 & n15656;
  assign n13160 = ~n13152;
  assign n16945 = n16955 & n16956;
  assign n16856 = n15731 & n15765;
  assign n16894 = ~n16906;
  assign n16895 = ~n16875;
  assign n16855 = ~n16915;
  assign n16908 = n16916 & n16917;
  assign n16900 = n16925 & n16926;
  assign n16817 = n16929 ^ n14319;
  assign n16937 = ~n16945;
  assign n16891 = n16894 & n16895;
  assign n16892 = n16894 & n16879;
  assign n16893 = n16900 ^ n16901;
  assign n16905 = n16817 & n16907;
  assign n16873 = ~n16908;
  assign n16902 = ~n16900;
  assign n16904 = ~n16817;
  assign n16918 = n16937 & n16938;
  assign n16878 = ~n16891;
  assign n16876 = ~n16892;
  assign n16888 = n16893 & n171;
  assign n16886 = ~n16893;
  assign n16870 = n16855 & n16873;
  assign n16896 = n16902 & n16903;
  assign n16897 = n16904 & n16837;
  assign n16819 = ~n16905;
  assign n13094 = n16918 ^ n16919;
  assign n16920 = ~n16918;
  assign n16857 = n16875 ^ n16876;
  assign n16845 = n16878 & n16879;
  assign n16880 = n16886 & n16887;
  assign n16844 = ~n16888;
  assign n16889 = ~n16896;
  assign n16839 = ~n16897;
  assign n13087 = ~n13094;
  assign n16909 = n16920 & n16921;
  assign n14931 = n16856 ^ n16857;
  assign n16828 = n16857 & n16856;
  assign n16861 = ~n16845;
  assign n16862 = ~n16880;
  assign n16871 = n16889 & n16890;
  assign n16881 = n13087 & n15510;
  assign n16898 = ~n16909;
  assign n12791 = n14931 ^ n13785;
  assign n14898 = n14931 ^ n16841;
  assign n16748 = n14931 & n13785;
  assign n16858 = n16861 & n16862;
  assign n16863 = n16862 & n16844;
  assign n16827 = n16870 ^ n16871;
  assign n16872 = ~n16871;
  assign n16769 = n16881 ^ n14282;
  assign n16882 = n16898 & n16899;
  assign n14897 = ~n12791;
  assign n16843 = ~n16858;
  assign n16852 = n16827 & n16859;
  assign n16846 = ~n16863;
  assign n16853 = ~n16827;
  assign n16864 = n16872 & n16873;
  assign n16866 = n16769 & n16874;
  assign n16865 = ~n16769;
  assign n16867 = n16882 ^ n16883;
  assign n16884 = ~n16882;
  assign n16800 = n14897 & n14886;
  assign n16826 = n16843 & n16844;
  assign n16829 = n16845 ^ n16846;
  assign n16831 = ~n16852;
  assign n16847 = n16853 & n170;
  assign n16854 = ~n16864;
  assign n16860 = n16865 & n16796;
  assign n16771 = ~n16866;
  assign n13073 = n16867 ^ n14223;
  assign n16877 = n16884 & n16885;
  assign n16778 = n16800 ^ n16801;
  assign n16774 = n16800 ^ n16802;
  assign n16806 = n16826 ^ n16827;
  assign n16815 = n16828 ^ n16829;
  assign n16780 = n16829 & n16828;
  assign n16830 = ~n16826;
  assign n16810 = ~n16847;
  assign n16836 = n16854 & n16855;
  assign n16840 = n13073 & n15551;
  assign n16798 = ~n16860;
  assign n13080 = ~n13073;
  assign n16868 = ~n16877;
  assign n14734 = n391 ^ n16774;
  assign n16752 = n16778 & n16779;
  assign n16578 = n16774 & n391;
  assign n16781 = n170 ^ n16806;
  assign n16808 = n16815 & n13692;
  assign n16807 = ~n16815;
  assign n16823 = n16830 & n16831;
  assign n16783 = ~n16780;
  assign n16816 = n16836 ^ n16837;
  assign n16824 = n16840 ^ n14223;
  assign n16838 = ~n16836;
  assign n16848 = n16868 & n16869;
  assign n16676 = n16752 ^ n16753;
  assign n16756 = n16752 & n16753;
  assign n16352 = ~n14734;
  assign n16754 = ~n16752;
  assign n16765 = n16780 ^ n16781;
  assign n16782 = ~n16781;
  assign n16804 = n16807 & n13680;
  assign n16759 = ~n16808;
  assign n16803 = n16816 ^ n16817;
  assign n16809 = ~n16823;
  assign n16820 = n16824 & n16825;
  assign n16821 = ~n16824;
  assign n16832 = n16838 & n16839;
  assign n16833 = n16848 ^ n16849;
  assign n16850 = ~n16848;
  assign n16746 = n16754 & n16755;
  assign n16658 = ~n16756;
  assign n16757 = n16765 & n13619;
  assign n16727 = ~n16765;
  assign n16708 = n16782 & n16783;
  assign n16794 = n16803 & n169;
  assign n16784 = ~n16804;
  assign n16735 = n16809 & n16810;
  assign n16792 = ~n16803;
  assign n16718 = ~n16820;
  assign n16811 = n16821 & n16822;
  assign n16818 = ~n16832;
  assign n12979 = n16833 ^ n14227;
  assign n16842 = n16850 & n16851;
  assign n16683 = ~n16746;
  assign n16747 = n16727 & n13626;
  assign n16724 = ~n16757;
  assign n16711 = ~n16708;
  assign n16775 = n16784 & n16748;
  assign n16776 = n16784 & n16759;
  assign n16785 = n16792 & n16793;
  assign n16737 = ~n16794;
  assign n16767 = ~n16735;
  assign n16744 = ~n16811;
  assign n16795 = n16818 & n16819;
  assign n16799 = n12979 & n15474;
  assign n13018 = ~n12979;
  assign n16834 = ~n16842;
  assign n16699 = ~n16747;
  assign n16758 = ~n16775;
  assign n16749 = ~n16776;
  assign n16766 = ~n16785;
  assign n16768 = n16795 ^ n16796;
  assign n16787 = n16718 & n16744;
  assign n16691 = n16799 ^ n14231;
  assign n16797 = ~n16795;
  assign n16812 = n16834 & n16835;
  assign n12700 = n16748 ^ n16749;
  assign n16726 = n16758 & n16759;
  assign n16760 = n16766 & n16767;
  assign n16734 = n16766 & n16737;
  assign n16750 = n16768 ^ n16769;
  assign n16772 = n16691 & n16777;
  assign n16742 = ~n16787;
  assign n16773 = ~n16691;
  assign n16786 = n16797 & n16798;
  assign n16789 = n16812 ^ n14153;
  assign n16813 = ~n16812;
  assign n16697 = n16726 ^ n16727;
  assign n16700 = n12700 & n14864;
  assign n16709 = n16734 ^ n16735;
  assign n12711 = ~n12700;
  assign n16725 = ~n16726;
  assign n16740 = n16750 & n168;
  assign n16736 = ~n16760;
  assign n16738 = ~n16750;
  assign n16693 = ~n16772;
  assign n16761 = n16773 & n16668;
  assign n16770 = ~n16786;
  assign n12944 = n16788 ^ n16789;
  assign n16805 = n16813 & n16814;
  assign n12565 = n13626 ^ n16697;
  assign n16677 = n16700 ^ n13680;
  assign n16695 = n16708 ^ n16709;
  assign n16721 = n16724 & n16725;
  assign n16710 = ~n16709;
  assign n16687 = n16736 & n16737;
  assign n16728 = n16738 & n16739;
  assign n16689 = ~n16740;
  assign n16670 = ~n16761;
  assign n16741 = n16770 & n16771;
  assign n16745 = n12944 & n15452;
  assign n12994 = ~n12944;
  assign n16790 = ~n16805;
  assign n16656 = n16676 ^ n16677;
  assign n16655 = n12565 & n14799;
  assign n16678 = n16677 & n16683;
  assign n12613 = ~n12565;
  assign n16684 = n16695 & n13571;
  assign n16685 = ~n16695;
  assign n16661 = n16710 & n16711;
  assign n16698 = ~n16721;
  assign n16712 = ~n16687;
  assign n16713 = ~n16728;
  assign n16722 = n16741 ^ n16742;
  assign n16600 = n16745 ^ n14153;
  assign n16743 = ~n16741;
  assign n16762 = n16790 & n16791;
  assign n16621 = n16655 ^ n13626;
  assign n16647 = n16656 & n390;
  assign n16645 = ~n16656;
  assign n16657 = ~n16678;
  assign n16627 = ~n16684;
  assign n16679 = n16685 & n13540;
  assign n16625 = n16698 & n16699;
  assign n16675 = ~n16661;
  assign n16701 = n16712 & n16713;
  assign n16686 = n16713 & n16689;
  assign n16716 = n16722 & n183;
  assign n16719 = n16600 & n16723;
  assign n16714 = ~n16722;
  assign n16720 = ~n16600;
  assign n16729 = n16743 & n16744;
  assign n16731 = n16762 ^ n14172;
  assign n16763 = ~n16762;
  assign n16604 = ~n16621;
  assign n16642 = n16645 & n16646;
  assign n16580 = ~n16647;
  assign n16620 = n16657 & n16658;
  assign n16660 = ~n16679;
  assign n16662 = n16686 ^ n16687;
  assign n16659 = ~n16625;
  assign n16688 = ~n16701;
  assign n16702 = n16714 & n16715;
  assign n16631 = ~n16716;
  assign n16602 = ~n16719;
  assign n16703 = n16720 & n16636;
  assign n16717 = ~n16729;
  assign n12906 = n16730 ^ n16731;
  assign n16751 = n16763 & n16764;
  assign n16589 = n16620 ^ n16621;
  assign n16611 = ~n16642;
  assign n16623 = n16620 & n16643;
  assign n16622 = ~n16620;
  assign n16648 = n16659 & n16660;
  assign n16624 = n16660 & n16627;
  assign n16572 = n16661 ^ n16662;
  assign n16628 = n16662 & n16675;
  assign n16664 = n16688 & n16689;
  assign n16666 = ~n16702;
  assign n16638 = ~n16703;
  assign n16690 = n16717 & n16718;
  assign n16694 = n12906 & n15392;
  assign n12937 = ~n12906;
  assign n16732 = ~n16751;
  assign n16567 = n16589 ^ n16590;
  assign n16606 = n16611 & n16578;
  assign n16577 = n16611 & n16580;
  assign n16612 = n16622 & n16590;
  assign n16605 = ~n16623;
  assign n12551 = n16624 ^ n16625;
  assign n16626 = ~n16648;
  assign n16665 = ~n16664;
  assign n16663 = n16666 & n16631;
  assign n16667 = n16690 ^ n16691;
  assign n16527 = n16694 ^ n14172;
  assign n16692 = ~n16690;
  assign n16705 = n16732 & n16733;
  assign n16552 = n16567 & n389;
  assign n16550 = ~n16567;
  assign n16537 = n16577 ^ n16578;
  assign n16591 = n16604 & n16605;
  assign n16579 = ~n16606;
  assign n16570 = n12551 & n14766;
  assign n16569 = ~n16612;
  assign n12568 = ~n12551;
  assign n16607 = n16626 & n16627;
  assign n16629 = n16663 ^ n16664;
  assign n16649 = n16665 & n16666;
  assign n16596 = n16667 ^ n16668;
  assign n16671 = n16527 & n16561;
  assign n16672 = ~n16527;
  assign n16680 = n16692 & n16693;
  assign n12893 = n16704 ^ n16705;
  assign n16706 = ~n16705;
  assign n16314 = n16537 ^ n14734;
  assign n16536 = n16550 & n16551;
  assign n16488 = ~n16552;
  assign n16538 = n16570 ^ n13540;
  assign n16540 = ~n16537;
  assign n16486 = n16579 & n16580;
  assign n16568 = ~n16591;
  assign n16593 = n16607 & n13519;
  assign n16581 = ~n16607;
  assign n16608 = n16628 ^ n16629;
  assign n16522 = n16629 & n16628;
  assign n16634 = n16596 & n182;
  assign n16630 = ~n16649;
  assign n16632 = ~n16596;
  assign n16529 = ~n16671;
  assign n16650 = n16672 & n16673;
  assign n16669 = ~n16680;
  assign n16674 = n12893 & n15374;
  assign n12904 = ~n12893;
  assign n16696 = n16706 & n16707;
  assign n16296 = ~n16314;
  assign n16519 = ~n16536;
  assign n16530 = n16538 & n16539;
  assign n16450 = n16540 & n16352;
  assign n16531 = ~n16538;
  assign n16456 = n16568 & n16569;
  assign n16520 = ~n16486;
  assign n16541 = n16581 ^ n16572;
  assign n16582 = n16581 & n13534;
  assign n16571 = ~n16593;
  assign n16594 = n16608 & n13486;
  assign n16592 = ~n16608;
  assign n16595 = n16630 & n16631;
  assign n16613 = n16632 & n16633;
  assign n16556 = ~n16634;
  assign n16563 = ~n16650;
  assign n16635 = n16669 & n16670;
  assign n16466 = n16674 ^ n14135;
  assign n16681 = ~n16696;
  assign n16512 = n16519 & n16520;
  assign n16485 = n16519 & n16488;
  assign n16470 = ~n16530;
  assign n16521 = n16531 & n16532;
  assign n16453 = ~n16450;
  assign n12381 = n13534 ^ n16541;
  assign n16504 = ~n16456;
  assign n16553 = n16571 & n16572;
  assign n16534 = ~n16582;
  assign n16583 = n16592 & n13496;
  assign n16509 = ~n16594;
  assign n16554 = n16595 ^ n16596;
  assign n16598 = ~n16595;
  assign n16597 = ~n16613;
  assign n16599 = n16635 ^ n16636;
  assign n16639 = n16466 & n16500;
  assign n16637 = ~n16635;
  assign n16640 = ~n16466;
  assign n16652 = n16681 & n16682;
  assign n16451 = n16485 ^ n16486;
  assign n16487 = ~n16512;
  assign n16503 = ~n16521;
  assign n12437 = ~n12381;
  assign n16533 = ~n16553;
  assign n16523 = n182 ^ n16554;
  assign n16472 = ~n16583;
  assign n16584 = n16597 & n16598;
  assign n16573 = n16599 ^ n16600;
  assign n16614 = n16637 & n16638;
  assign n16502 = ~n16639;
  assign n16615 = n16640 & n16641;
  assign n12784 = n16651 ^ n16652;
  assign n16653 = ~n16652;
  assign n16181 = n16450 ^ n16451;
  assign n16452 = ~n16451;
  assign n16410 = n16487 & n16488;
  assign n16489 = n16503 & n16504;
  assign n16490 = n16470 & n16503;
  assign n16474 = n12437 & n14694;
  assign n16505 = n16522 ^ n16523;
  assign n16506 = n16533 & n16534;
  assign n16458 = n16523 & n16522;
  assign n16542 = n16509 & n16472;
  assign n16559 = n16573 & n181;
  assign n16555 = ~n16584;
  assign n16557 = ~n16573;
  assign n16601 = ~n16614;
  assign n16468 = ~n16615;
  assign n16616 = n12784 & n16609;
  assign n16603 = n12784 & n15329;
  assign n12845 = ~n12784;
  assign n16644 = n16653 & n16654;
  assign n16191 = ~n16181;
  assign n16327 = n16452 & n16453;
  assign n16370 = ~n16410;
  assign n16454 = n16474 ^ n13519;
  assign n16469 = ~n16489;
  assign n16457 = ~n16490;
  assign n16491 = n16505 & n13401;
  assign n16433 = ~n16505;
  assign n16508 = ~n16506;
  assign n16461 = ~n16458;
  assign n16507 = ~n16542;
  assign n16494 = n16555 & n16556;
  assign n16543 = n16557 & n16558;
  assign n16496 = ~n16559;
  assign n16560 = n16601 & n16602;
  assign n16574 = n16603 ^ n14018;
  assign n15384 = n16609 ^ n12845;
  assign n15386 = ~n16616;
  assign n16610 = n12845 & n16617;
  assign n16618 = ~n16644;
  assign n16442 = n16454 & n16455;
  assign n16411 = n16456 ^ n16457;
  assign n16349 = n16469 & n16470;
  assign n16440 = ~n16454;
  assign n16475 = n16433 & n13458;
  assign n16434 = ~n16491;
  assign n12265 = n16506 ^ n16507;
  assign n16492 = n16508 & n16509;
  assign n16524 = ~n16494;
  assign n16525 = ~n16543;
  assign n16526 = n16560 ^ n16561;
  assign n16564 = n16574 & n16575;
  assign n16562 = ~n16560;
  assign n16565 = ~n16574;
  assign n15360 = ~n16610;
  assign n16585 = n16618 & n16619;
  assign n16368 = n16410 ^ n16411;
  assign n16414 = n16411 & n388;
  assign n16430 = n16440 & n16441;
  assign n16359 = ~n16442;
  assign n16412 = ~n16411;
  assign n16399 = ~n16349;
  assign n16393 = ~n16475;
  assign n12386 = ~n12265;
  assign n16471 = ~n16492;
  assign n16513 = n16524 & n16525;
  assign n16493 = n16525 & n16496;
  assign n16419 = n16526 ^ n16527;
  assign n16544 = n16562 & n16563;
  assign n16381 = ~n16564;
  assign n16545 = n16565 & n16566;
  assign n12838 = n16585 ^ n16586;
  assign n16587 = ~n16585;
  assign n16328 = n388 ^ n16368;
  assign n16400 = n16412 & n16413;
  assign n16331 = ~n16414;
  assign n16398 = ~n16430;
  assign n16431 = n12386 & n14707;
  assign n16432 = n16471 & n16472;
  assign n16459 = n16493 ^ n16494;
  assign n16497 = n16419 & n16510;
  assign n16495 = ~n16513;
  assign n16498 = ~n16419;
  assign n16528 = ~n16544;
  assign n16427 = ~n16545;
  assign n16546 = n12838 & n15322;
  assign n12830 = ~n12838;
  assign n16576 = n16587 & n16588;
  assign n14628 = n16327 ^ n16328;
  assign n16329 = ~n16328;
  assign n16386 = n16398 & n16399;
  assign n16369 = ~n16400;
  assign n16387 = n16359 & n16398;
  assign n16401 = n16431 ^ n13486;
  assign n16391 = n16432 ^ n16433;
  assign n16435 = ~n16432;
  assign n16436 = n16458 ^ n16459;
  assign n16460 = ~n16459;
  assign n16462 = n16495 & n16496;
  assign n16464 = ~n16497;
  assign n16476 = n16498 & n180;
  assign n16499 = n16528 & n16529;
  assign n16514 = n16427 & n16381;
  assign n15324 = ~n16546;
  assign n16535 = n12830 & n16547;
  assign n16515 = n12830 & n15261;
  assign n16548 = ~n16576;
  assign n16126 = ~n14628;
  assign n16158 = n16329 & n16327;
  assign n16360 = n16369 & n16370;
  assign n16358 = ~n16386;
  assign n16350 = ~n16387;
  assign n12297 = n16391 ^ n13458;
  assign n16388 = n16401 & n16402;
  assign n16389 = ~n16401;
  assign n16415 = n16434 & n16435;
  assign n16416 = n16436 & n13397;
  assign n16417 = ~n16436;
  assign n16372 = n16460 & n16461;
  assign n16418 = n180 ^ n16462;
  assign n16463 = ~n16462;
  assign n16421 = ~n16476;
  assign n16465 = n16499 ^ n16500;
  assign n16501 = ~n16499;
  assign n16425 = ~n16514;
  assign n16344 = n16515 ^ n14000;
  assign n15342 = ~n16535;
  assign n16516 = n16548 & n16549;
  assign n16317 = n16349 ^ n16350;
  assign n16293 = n16358 & n16359;
  assign n16330 = ~n16360;
  assign n16318 = n12297 & n14673;
  assign n16351 = n12297 & n14734;
  assign n12308 = ~n12297;
  assign n16284 = ~n16388;
  assign n16371 = n16389 & n16390;
  assign n16392 = ~n16415;
  assign n16316 = ~n16416;
  assign n16403 = n16417 & n13391;
  assign n16373 = n16418 ^ n16419;
  assign n16443 = n16463 & n16464;
  assign n16340 = n16465 ^ n16466;
  assign n16477 = n16501 & n16502;
  assign n16478 = n16344 & n16306;
  assign n16479 = ~n16344;
  assign n16482 = n16516 ^ n13958;
  assign n16517 = ~n16516;
  assign n16312 = n16317 & n387;
  assign n16221 = n16318 ^ n13401;
  assign n16200 = n16330 & n16331;
  assign n16310 = ~n16317;
  assign n16319 = ~n16293;
  assign n14736 = ~n16351;
  assign n16333 = n12308 & n16352;
  assign n16320 = ~n16371;
  assign n16274 = n16372 ^ n16373;
  assign n16337 = n16392 & n16393;
  assign n16297 = n16373 & n16372;
  assign n16354 = ~n16403;
  assign n16422 = n16340 & n16437;
  assign n16420 = ~n16443;
  assign n16423 = ~n16340;
  assign n16467 = ~n16477;
  assign n16308 = ~n16478;
  assign n16473 = n16479 & n16480;
  assign n12706 = n16481 ^ n16482;
  assign n16511 = n16517 & n16518;
  assign n16282 = n16221 & n16178;
  assign n16292 = n16310 & n16311;
  assign n16219 = ~n16312;
  assign n16280 = ~n16221;
  assign n16313 = n16319 & n16320;
  assign n16267 = ~n16200;
  assign n14721 = ~n16333;
  assign n16332 = n16320 & n16284;
  assign n16335 = n16274 & n13360;
  assign n16334 = ~n16274;
  assign n16353 = ~n16337;
  assign n16336 = n16354 & n16316;
  assign n16300 = ~n16297;
  assign n16374 = n16420 & n16421;
  assign n16376 = ~n16422;
  assign n16404 = n16423 & n179;
  assign n16424 = n16467 & n16468;
  assign n16428 = n12706 & n15228;
  assign n16445 = n12706 & n15278;
  assign n16346 = ~n16473;
  assign n12777 = ~n12706;
  assign n16483 = ~n16511;
  assign n16268 = n16280 & n16281;
  assign n16189 = ~n16282;
  assign n16266 = ~n16292;
  assign n16283 = ~n16313;
  assign n16294 = ~n16332;
  assign n16321 = n16334 & n13349;
  assign n16228 = ~n16335;
  assign n12235 = n16336 ^ n16337;
  assign n16338 = n16353 & n16354;
  assign n16339 = n179 ^ n16374;
  assign n16375 = ~n16374;
  assign n16342 = ~n16404;
  assign n16394 = n16424 ^ n16425;
  assign n16395 = n16428 ^ n13958;
  assign n16426 = ~n16424;
  assign n16438 = n12777 & n16444;
  assign n15302 = ~n16445;
  assign n16447 = n16483 & n16484;
  assign n16244 = n16266 & n16267;
  assign n16247 = n16266 & n16219;
  assign n16233 = ~n16268;
  assign n16270 = n16283 & n16284;
  assign n16269 = n16293 ^ n16294;
  assign n16271 = n12235 & n14654;
  assign n16295 = n12235 & n16314;
  assign n16276 = ~n16321;
  assign n12248 = ~n12235;
  assign n16315 = ~n16338;
  assign n16298 = n16339 ^ n16340;
  assign n16361 = n16375 & n16376;
  assign n16379 = n16394 & n178;
  assign n16382 = n16395 & n16396;
  assign n16377 = ~n16394;
  assign n16383 = ~n16395;
  assign n16405 = n16426 & n16427;
  assign n15281 = ~n16438;
  assign n12725 = n16446 ^ n16447;
  assign n16448 = ~n16447;
  assign n16218 = ~n16244;
  assign n16201 = ~n16247;
  assign n16248 = n16269 & n386;
  assign n16220 = ~n16270;
  assign n16235 = n16271 ^ n13391;
  assign n16245 = ~n16269;
  assign n14701 = ~n16295;
  assign n16285 = n12248 & n16296;
  assign n16272 = n16297 ^ n16298;
  assign n16273 = n16315 & n16316;
  assign n16299 = ~n16298;
  assign n16341 = ~n16361;
  assign n16362 = n16377 & n16378;
  assign n16257 = ~n16379;
  assign n16212 = ~n16382;
  assign n16363 = n16383 & n16384;
  assign n16380 = ~n16405;
  assign n16385 = n12725 & n15211;
  assign n16407 = n12725 & n16429;
  assign n12739 = ~n12725;
  assign n16439 = n16448 & n16449;
  assign n16159 = n16200 ^ n16201;
  assign n16149 = n16218 & n16219;
  assign n16177 = n16220 ^ n16221;
  assign n16217 = n16233 & n16220;
  assign n16222 = n16235 & n16236;
  assign n16234 = n16245 & n16246;
  assign n16142 = ~n16248;
  assign n16223 = ~n16235;
  assign n16250 = n16272 & n13296;
  assign n16225 = n16273 ^ n16274;
  assign n14684 = ~n16285;
  assign n16249 = ~n16272;
  assign n16275 = ~n16273;
  assign n16251 = n16299 & n16300;
  assign n16302 = n16341 & n16342;
  assign n16304 = ~n16362;
  assign n16263 = ~n16363;
  assign n16343 = n16380 & n16381;
  assign n16134 = n16385 ^ n13946;
  assign n16397 = n12739 & n16406;
  assign n15266 = ~n16407;
  assign n16408 = ~n16439;
  assign n16059 = n16158 ^ n16159;
  assign n16104 = n16159 & n16158;
  assign n16075 = n16177 ^ n16178;
  assign n16179 = ~n16149;
  assign n16188 = ~n16217;
  assign n16107 = ~n16222;
  assign n16202 = n16223 & n16224;
  assign n12110 = n13360 ^ n16225;
  assign n16180 = ~n16234;
  assign n14698 = n14701 & n14684;
  assign n16237 = n16249 & n13327;
  assign n16183 = ~n16250;
  assign n16253 = n16275 & n16276;
  assign n16255 = ~n16251;
  assign n16303 = ~n16302;
  assign n16301 = n16304 & n16257;
  assign n16305 = n16343 ^ n16344;
  assign n16260 = n16263 & n16212;
  assign n16347 = n16134 & n16355;
  assign n16345 = ~n16343;
  assign n16348 = ~n16134;
  assign n15238 = ~n16397;
  assign n16364 = n16408 & n16409;
  assign n16139 = n16075 & n385;
  assign n16048 = ~n16059;
  assign n16137 = ~n16075;
  assign n16160 = n16179 & n16180;
  assign n16122 = n16188 & n16189;
  assign n16148 = n12110 & n14613;
  assign n16182 = n12110 & n16191;
  assign n16190 = n16180 & n16142;
  assign n16147 = ~n16202;
  assign n12171 = ~n12110;
  assign n16144 = ~n16237;
  assign n16227 = ~n16253;
  assign n16252 = n16301 ^ n16302;
  assign n16286 = n16303 & n16304;
  assign n16206 = n16305 ^ n16306;
  assign n16322 = n16345 & n16346;
  assign n16136 = ~n16347;
  assign n16323 = n16348 & n16170;
  assign n16356 = n15266 & n15238;
  assign n16324 = n16364 ^ n16365;
  assign n16366 = ~n16364;
  assign n16119 = n16137 & n16138;
  assign n16041 = ~n16139;
  assign n16120 = n16148 ^ n13349;
  assign n16141 = ~n16160;
  assign n16146 = ~n16122;
  assign n16161 = n16107 & n16147;
  assign n16162 = n12171 & n16181;
  assign n14664 = ~n16182;
  assign n16150 = ~n16190;
  assign n16163 = n16144 & n16183;
  assign n16164 = n16227 & n16228;
  assign n16226 = n16251 ^ n16252;
  assign n16258 = n16206 & n16277;
  assign n16254 = ~n16252;
  assign n16256 = ~n16286;
  assign n16259 = ~n16206;
  assign n16307 = ~n16322;
  assign n16172 = ~n16323;
  assign n12677 = n13858 ^ n16324;
  assign n15264 = ~n16356;
  assign n16357 = n16366 & n16367;
  assign n16093 = ~n16119;
  assign n16108 = n16120 & n16121;
  assign n16124 = n16141 & n16142;
  assign n16109 = ~n16120;
  assign n16140 = n16146 & n16147;
  assign n16105 = n16149 ^ n16150;
  assign n16123 = ~n16161;
  assign n14645 = ~n16162;
  assign n12094 = n16163 ^ n16164;
  assign n16184 = ~n16164;
  assign n16204 = n16226 & n13303;
  assign n16203 = ~n16226;
  assign n16128 = n16254 & n16255;
  assign n16205 = n16256 & n16257;
  assign n16208 = ~n16258;
  assign n16238 = n16259 & n177;
  assign n16261 = n16307 & n16308;
  assign n16264 = n12677 & n15148;
  assign n16287 = n12677 & n16309;
  assign n12543 = ~n12677;
  assign n16325 = ~n16357;
  assign n15941 = n16104 ^ n16105;
  assign n16019 = ~n16108;
  assign n16095 = n16109 & n16110;
  assign n15980 = n16105 & n16104;
  assign n16094 = n16122 ^ n16123;
  assign n16074 = ~n16124;
  assign n16106 = ~n16140;
  assign n16125 = n12094 & n14628;
  assign n16127 = n14664 & n14645;
  assign n16096 = n12094 & n14559;
  assign n12060 = ~n12094;
  assign n16165 = n16183 & n16184;
  assign n16192 = n16203 & n13235;
  assign n16050 = ~n16204;
  assign n16166 = n16205 ^ n16206;
  assign n16207 = ~n16205;
  assign n16168 = ~n16238;
  assign n16080 = n16260 ^ n16261;
  assign n16230 = n16264 ^ n13910;
  assign n16262 = ~n16261;
  assign n16278 = n12543 & n15200;
  assign n15221 = ~n16287;
  assign n16289 = n16325 & n16326;
  assign n16026 = n16074 ^ n16075;
  assign n16070 = n16093 & n16074;
  assign n16073 = n16094 & n384;
  assign n15964 = ~n15941;
  assign n16054 = ~n16095;
  assign n16057 = n16096 ^ n13296;
  assign n16008 = n16106 & n16107;
  assign n15983 = ~n15980;
  assign n16071 = ~n16094;
  assign n14630 = ~n16125;
  assign n16111 = n12060 & n16126;
  assign n14662 = ~n16127;
  assign n16143 = ~n16165;
  assign n16129 = n177 ^ n16166;
  assign n16101 = ~n16192;
  assign n16193 = n16207 & n16208;
  assign n16209 = n16080 & n16229;
  assign n16213 = n16230 & n16231;
  assign n16210 = ~n16080;
  assign n16214 = ~n16230;
  assign n16239 = n16262 & n16263;
  assign n15203 = ~n16278;
  assign n12574 = n16288 ^ n16289;
  assign n16290 = ~n16289;
  assign n15981 = n385 ^ n16026;
  assign n16043 = n16019 & n16054;
  assign n16046 = n16057 & n16058;
  assign n16040 = ~n16070;
  assign n16056 = n16071 & n16072;
  assign n15956 = ~n16073;
  assign n16044 = ~n16057;
  assign n16055 = ~n16008;
  assign n14610 = ~n16111;
  assign n16097 = n16128 ^ n16129;
  assign n16098 = n16143 & n16144;
  assign n16029 = n16129 & n16128;
  assign n16151 = n16101 & n16050;
  assign n16167 = ~n16193;
  assign n16132 = ~n16209;
  assign n16194 = n16210 & n176;
  assign n16038 = ~n16213;
  assign n16195 = n16214 & n16215;
  assign n16211 = ~n16239;
  assign n16216 = n12574 & n15132;
  assign n16240 = n12574 & n16265;
  assign n12582 = ~n12574;
  assign n16279 = n16290 & n16291;
  assign n15871 = n15980 ^ n15981;
  assign n15982 = ~n15981;
  assign n15985 = n16040 & n16041;
  assign n16009 = ~n16043;
  assign n16027 = n16044 & n16045;
  assign n15925 = ~n16046;
  assign n16042 = n16054 & n16055;
  assign n16007 = ~n16056;
  assign n16076 = n16097 & n13277;
  assign n16077 = ~n16097;
  assign n16100 = ~n16098;
  assign n16032 = ~n16029;
  assign n16099 = ~n16151;
  assign n16130 = n16167 & n16168;
  assign n16082 = ~n16194;
  assign n16089 = ~n16195;
  assign n16169 = n16211 & n16212;
  assign n16185 = n16216 ^ n13835;
  assign n15180 = ~n16240;
  assign n16232 = n12582 & n16241;
  assign n16242 = ~n16279;
  assign n15850 = ~n15871;
  assign n15935 = n15982 & n15983;
  assign n15969 = n16008 ^ n16009;
  assign n16006 = ~n15985;
  assign n15984 = n16007 & n15956;
  assign n15971 = ~n16027;
  assign n16018 = ~n16042;
  assign n15966 = ~n16076;
  assign n16060 = n16077 & n13268;
  assign n12051 = n16098 ^ n16099;
  assign n16078 = n16100 & n16101;
  assign n16079 = n176 ^ n16130;
  assign n16131 = ~n16130;
  assign n16133 = n16169 ^ n16170;
  assign n16086 = n16089 & n16038;
  assign n16175 = n16185 & n16186;
  assign n16171 = ~n16169;
  assign n16173 = ~n16185;
  assign n15165 = ~n16232;
  assign n16196 = n16242 & n16243;
  assign n15959 = n15969 & n399;
  assign n15936 = n15984 ^ n15985;
  assign n15957 = ~n15969;
  assign n15986 = n16006 & n16007;
  assign n15987 = n15925 & n15971;
  assign n15938 = n16018 & n16019;
  assign n16047 = n12051 & n16059;
  assign n16013 = ~n16060;
  assign n12016 = ~n12051;
  assign n16049 = ~n16078;
  assign n16030 = n16079 ^ n16080;
  assign n16112 = n16131 & n16132;
  assign n16102 = n16133 ^ n16134;
  assign n16152 = n16171 & n16172;
  assign n16153 = n16173 & n16174;
  assign n15954 = ~n16175;
  assign n15177 = n15180 & n15165;
  assign n12392 = n16196 ^ n16197;
  assign n16198 = ~n16196;
  assign n14465 = n15935 ^ n15936;
  assign n15827 = n15936 & n15935;
  assign n15937 = n15957 & n15958;
  assign n15870 = ~n15959;
  assign n15955 = ~n15986;
  assign n15939 = ~n15987;
  assign n15970 = ~n15938;
  assign n15989 = n16013 & n15966;
  assign n16011 = n16029 ^ n16030;
  assign n14572 = ~n16047;
  assign n16028 = n12016 & n16048;
  assign n16010 = n12016 & n14523;
  assign n15990 = n16049 & n16050;
  assign n16031 = ~n16030;
  assign n16085 = n16102 & n191;
  assign n16081 = ~n16112;
  assign n16083 = ~n16102;
  assign n16135 = ~n16152;
  assign n16001 = ~n16153;
  assign n16154 = n12392 & n16176;
  assign n12506 = ~n12392;
  assign n16187 = n16198 & n16199;
  assign n15759 = ~n14465;
  assign n15917 = ~n15937;
  assign n15919 = n15938 ^ n15939;
  assign n15868 = n15955 & n15956;
  assign n15960 = n15970 & n15971;
  assign n12000 = n15989 ^ n15990;
  assign n15972 = n16010 ^ n13235;
  assign n15991 = n16011 & n13233;
  assign n15992 = ~n16011;
  assign n14591 = ~n16028;
  assign n16012 = ~n15990;
  assign n15943 = n16031 & n16032;
  assign n15995 = n16081 & n16082;
  assign n16061 = n16083 & n16084;
  assign n15997 = ~n16085;
  assign n16087 = n16135 & n16136;
  assign n16113 = n16001 & n15954;
  assign n16114 = n12506 & n15088;
  assign n15117 = ~n16154;
  assign n16145 = n12506 & n16155;
  assign n16156 = ~n16187;
  assign n15867 = n15917 & n15870;
  assign n15898 = n15919 & n398;
  assign n15896 = ~n15919;
  assign n15918 = ~n15868;
  assign n15924 = ~n15960;
  assign n15920 = n12000 & n14498;
  assign n15942 = n12000 & n15964;
  assign n15961 = n15972 & n15973;
  assign n12011 = ~n12000;
  assign n15962 = ~n15972;
  assign n15922 = ~n15991;
  assign n15974 = n15992 & n13239;
  assign n15988 = n14591 & n14572;
  assign n15993 = n16012 & n16013;
  assign n15946 = ~n15943;
  assign n16033 = ~n15995;
  assign n16034 = ~n16061;
  assign n15906 = n16086 ^ n16087;
  assign n16088 = ~n16087;
  assign n15999 = ~n16113;
  assign n16090 = n16114 ^ n13839;
  assign n15144 = ~n16145;
  assign n16116 = n16156 & n16157;
  assign n15828 = n15867 ^ n15868;
  assign n15884 = n15896 & n15897;
  assign n15783 = ~n15898;
  assign n15895 = n15917 & n15918;
  assign n15794 = n15920 ^ n13277;
  assign n15852 = n15924 & n15925;
  assign n15926 = n12011 & n15941;
  assign n14548 = ~n15942;
  assign n15841 = ~n15961;
  assign n15940 = n15962 & n15963;
  assign n15877 = ~n15974;
  assign n14589 = ~n15988;
  assign n15965 = ~n15993;
  assign n16020 = n16033 & n16034;
  assign n15994 = n16034 & n15997;
  assign n16035 = n15906 & n16051;
  assign n16036 = ~n15906;
  assign n16062 = n16088 & n16089;
  assign n16065 = n16090 & n16091;
  assign n16063 = ~n16090;
  assign n15141 = n15144 & n15117;
  assign n12448 = n16115 ^ n16116;
  assign n16117 = ~n16116;
  assign n15716 = n15827 ^ n15828;
  assign n15766 = n15828 & n15827;
  assign n15830 = ~n15884;
  assign n15875 = n15794 & n15756;
  assign n15869 = ~n15895;
  assign n15873 = ~n15794;
  assign n15882 = ~n15852;
  assign n14528 = ~n15926;
  assign n15883 = ~n15940;
  assign n15900 = n15877 & n15922;
  assign n15901 = n15965 & n15966;
  assign n15944 = n15994 ^ n15995;
  assign n15996 = ~n16020;
  assign n15949 = ~n16035;
  assign n16021 = n16036 & n190;
  assign n16037 = ~n16062;
  assign n16052 = n16063 & n16064;
  assign n15863 = ~n16065;
  assign n16039 = n12448 & n15044;
  assign n16066 = n12448 & n16092;
  assign n12459 = ~n12448;
  assign n16103 = n16117 & n16118;
  assign n15700 = ~n15716;
  assign n15769 = ~n15766;
  assign n15809 = n15830 & n15783;
  assign n15810 = n15869 & n15870;
  assign n15854 = n15873 & n15874;
  assign n15796 = ~n15875;
  assign n15872 = n15882 & n15883;
  assign n14545 = n14548 & n14528;
  assign n11939 = n15900 ^ n15901;
  assign n15899 = n15841 & n15883;
  assign n15921 = ~n15901;
  assign n15788 = n15943 ^ n15944;
  assign n15945 = ~n15944;
  assign n15947 = n15996 & n15997;
  assign n15908 = ~n16021;
  assign n15998 = n16037 & n16038;
  assign n16014 = n16039 ^ n13792;
  assign n15912 = ~n16052;
  assign n15097 = ~n16066;
  assign n16053 = n12459 & n16067;
  assign n16068 = ~n16103;
  assign n15767 = n15809 ^ n15810;
  assign n15829 = ~n15810;
  assign n15758 = ~n15854;
  assign n15851 = n11939 & n15871;
  assign n15840 = ~n15872;
  assign n15832 = n11939 & n14454;
  assign n11978 = ~n11939;
  assign n15853 = ~n15899;
  assign n15902 = n15921 & n15922;
  assign n15903 = n15788 & n13178;
  assign n15904 = ~n15788;
  assign n15855 = n15945 & n15946;
  assign n15905 = n190 ^ n15947;
  assign n15948 = ~n15947;
  assign n15967 = n15998 ^ n15999;
  assign n16002 = n16014 & n16015;
  assign n16000 = ~n15998;
  assign n16016 = n15912 & n15863;
  assign n16003 = ~n16014;
  assign n15075 = ~n16053;
  assign n16022 = n16068 & n16069;
  assign n15657 = n15766 ^ n15767;
  assign n15768 = ~n15767;
  assign n15811 = n15829 & n15830;
  assign n15798 = n15832 ^ n13233;
  assign n15793 = n15840 & n15841;
  assign n15842 = n11978 & n15850;
  assign n14505 = ~n15851;
  assign n15831 = n15852 ^ n15853;
  assign n15876 = ~n15902;
  assign n15791 = ~n15903;
  assign n15885 = n15904 & n13139;
  assign n15856 = n15905 ^ n15906;
  assign n15927 = n15948 & n15949;
  assign n15952 = n15967 & n189;
  assign n15950 = ~n15967;
  assign n15975 = n16000 & n16001;
  assign n15780 = ~n16002;
  assign n15976 = n16003 & n16004;
  assign n15910 = ~n16016;
  assign n15094 = n15097 & n15075;
  assign n12240 = n16022 ^ n16023;
  assign n16024 = ~n16022;
  assign n15651 = ~n15657;
  assign n15696 = n15768 & n15769;
  assign n15755 = n15793 ^ n15794;
  assign n15785 = n15798 & n15799;
  assign n15782 = ~n15811;
  assign n15786 = ~n15798;
  assign n15814 = n15831 & n397;
  assign n15795 = ~n15793;
  assign n14484 = ~n15842;
  assign n15812 = ~n15831;
  assign n15833 = n15855 ^ n15856;
  assign n15834 = n15876 & n15877;
  assign n15801 = n15856 & n15855;
  assign n15836 = ~n15885;
  assign n15907 = ~n15927;
  assign n15928 = n15950 & n15951;
  assign n15819 = ~n15952;
  assign n15953 = ~n15975;
  assign n15823 = ~n15976;
  assign n15977 = n12240 & n16005;
  assign n12355 = ~n12240;
  assign n16017 = n16024 & n16025;
  assign n15643 = n15755 ^ n15756;
  assign n15734 = n15782 & n15783;
  assign n15690 = ~n15785;
  assign n15770 = n15786 & n15787;
  assign n15784 = n15795 & n15796;
  assign n15797 = n15812 & n15813;
  assign n14502 = n14505 & n14484;
  assign n15715 = ~n15814;
  assign n15816 = n15833 & n13160;
  assign n15789 = n15834 ^ n13139;
  assign n15815 = ~n15833;
  assign n15835 = ~n15834;
  assign n15804 = ~n15801;
  assign n15843 = n15907 & n15908;
  assign n15858 = ~n15928;
  assign n15909 = n15953 & n15954;
  assign n15929 = n15823 & n15780;
  assign n15930 = n12355 & n14928;
  assign n15968 = n12355 & n15051;
  assign n15033 = ~n15977;
  assign n15978 = ~n16017;
  assign n15723 = n15643 & n15732;
  assign n15724 = ~n15643;
  assign n15749 = ~n15734;
  assign n15726 = ~n15770;
  assign n15757 = ~n15784;
  assign n11936 = n15788 ^ n15789;
  assign n15750 = ~n15797;
  assign n15800 = n15815 & n13152;
  assign n15720 = ~n15816;
  assign n15817 = n15835 & n15836;
  assign n15857 = ~n15843;
  assign n15886 = n15858 & n15819;
  assign n15878 = n15909 ^ n15910;
  assign n15911 = ~n15909;
  assign n15821 = ~n15929;
  assign n15710 = n15930 ^ n13664;
  assign n15053 = ~n15968;
  assign n15932 = n15978 & n15979;
  assign n15677 = ~n15723;
  assign n15713 = n15724 & n396;
  assign n15735 = n15749 & n15750;
  assign n15736 = n15690 & n15726;
  assign n15701 = n15757 & n15758;
  assign n15751 = n11936 & n15759;
  assign n15733 = n15750 & n15715;
  assign n11931 = ~n11936;
  assign n15753 = ~n15800;
  assign n15790 = ~n15817;
  assign n15845 = n15857 & n15858;
  assign n15861 = n15878 & n188;
  assign n15844 = ~n15886;
  assign n15859 = ~n15878;
  assign n15887 = n15911 & n15912;
  assign n15889 = n15710 & n15913;
  assign n15888 = ~n15710;
  assign n12260 = n15931 ^ n15932;
  assign n15934 = n15932 & n15893;
  assign n15933 = ~n15932;
  assign n15645 = ~n15713;
  assign n15697 = n15733 ^ n15734;
  assign n15714 = ~n15735;
  assign n15702 = ~n15736;
  assign n15725 = ~n15701;
  assign n15718 = n11931 & n14340;
  assign n14443 = ~n15751;
  assign n15737 = n11931 & n14465;
  assign n15738 = n15753 & n15720;
  assign n15739 = n15790 & n15791;
  assign n15802 = n15843 ^ n15844;
  assign n15818 = ~n15845;
  assign n15846 = n15859 & n15860;
  assign n15743 = ~n15861;
  assign n15862 = ~n15887;
  assign n15879 = n15888 & n15745;
  assign n15712 = ~n15889;
  assign n15864 = n12260 & n14913;
  assign n15891 = n12260 & n15914;
  assign n12272 = ~n12260;
  assign n15923 = n15933 & n15916;
  assign n15915 = ~n15934;
  assign n14323 = n15696 ^ n15697;
  assign n15587 = n15701 ^ n15702;
  assign n15679 = n15714 & n15715;
  assign n15691 = n15718 ^ n13139;
  assign n15698 = ~n15697;
  assign n15717 = n15725 & n15726;
  assign n14467 = ~n15737;
  assign n11862 = n15738 ^ n15739;
  assign n15752 = ~n15739;
  assign n15771 = n15801 ^ n15802;
  assign n15773 = n15818 & n15819;
  assign n15803 = ~n15802;
  assign n15775 = ~n15846;
  assign n15820 = n15862 & n15863;
  assign n15837 = n15864 ^ n13677;
  assign n15747 = ~n15879;
  assign n15880 = n12272 & n15890;
  assign n15005 = ~n15891;
  assign n15894 = n15915 & n15916;
  assign n15892 = ~n15923;
  assign n15642 = n396 ^ n15679;
  assign n15663 = n15587 & n395;
  assign n15594 = ~n14323;
  assign n15682 = n15691 & n15692;
  assign n15661 = ~n15587;
  assign n15612 = n15698 & n15696;
  assign n15678 = ~n15679;
  assign n15680 = ~n15691;
  assign n15699 = n11862 & n15716;
  assign n15689 = ~n15717;
  assign n15683 = n11862 & n14373;
  assign n11891 = ~n11862;
  assign n15740 = n15752 & n15753;
  assign n15761 = n15771 & n13087;
  assign n15760 = ~n15771;
  assign n15727 = n15803 & n15804;
  assign n15774 = ~n15773;
  assign n15772 = n15775 & n15743;
  assign n15792 = n15820 ^ n15821;
  assign n15824 = n15837 & n15838;
  assign n15822 = ~n15820;
  assign n15825 = ~n15837;
  assign n14996 = ~n15880;
  assign n15881 = n15892 & n15893;
  assign n15865 = ~n15894;
  assign n15613 = n15642 ^ n15643;
  assign n15655 = n15661 & n15662;
  assign n15589 = ~n15663;
  assign n15660 = n15677 & n15678;
  assign n15664 = n15680 & n15681;
  assign n15620 = ~n15682;
  assign n15564 = n15683 ^ n13152;
  assign n15615 = ~n15612;
  assign n15603 = n15689 & n15690;
  assign n14427 = ~n15699;
  assign n15693 = n11891 & n15700;
  assign n15719 = ~n15740;
  assign n15754 = n15760 & n13094;
  assign n15687 = ~n15761;
  assign n15741 = n15772 ^ n15773;
  assign n15762 = n15774 & n15775;
  assign n15778 = n15792 & n187;
  assign n15776 = ~n15792;
  assign n15805 = n15822 & n15823;
  assign n15641 = ~n15824;
  assign n15806 = n15825 & n15826;
  assign n15015 = n15005 & n14996;
  assign n15849 = n15865 & n15866;
  assign n15847 = ~n15881;
  assign n15512 = n15612 ^ n15613;
  assign n15614 = ~n15613;
  assign n15618 = ~n15655;
  assign n15648 = n15564 & n15656;
  assign n15644 = ~n15660;
  assign n15646 = ~n15664;
  assign n15649 = ~n15564;
  assign n15647 = ~n15603;
  assign n14406 = ~n15693;
  assign n15684 = n15719 & n15720;
  assign n15722 = n15727 ^ n15741;
  assign n15653 = ~n15754;
  assign n15666 = n15741 & n15727;
  assign n15728 = ~n15741;
  assign n15742 = ~n15762;
  assign n15763 = n15776 & n15777;
  assign n15669 = ~n15778;
  assign n15779 = ~n15805;
  assign n15676 = ~n15806;
  assign n15839 = n15847 & n15848;
  assign n15808 = ~n15849;
  assign n14285 = ~n15512;
  assign n15558 = n15614 & n15615;
  assign n15616 = n15644 & n15645;
  assign n15629 = n15646 & n15647;
  assign n15630 = n15620 & n15646;
  assign n15566 = ~n15648;
  assign n15631 = n15649 & n15591;
  assign n14424 = n14427 & n14406;
  assign n15686 = ~n15684;
  assign n15704 = n15722 & n13073;
  assign n15721 = n15653 & n15687;
  assign n15703 = n15727 ^ n15728;
  assign n15706 = n15742 & n15743;
  assign n15708 = ~n15763;
  assign n15744 = n15779 & n15780;
  assign n15764 = n15676 & n15641;
  assign n15807 = ~n15839;
  assign n15586 = n395 ^ n15616;
  assign n15617 = ~n15616;
  assign n15619 = ~n15629;
  assign n15604 = ~n15630;
  assign n15593 = ~n15631;
  assign n15665 = n15686 & n15687;
  assign n15694 = n15703 & n13080;
  assign n15625 = ~n15704;
  assign n15685 = ~n15721;
  assign n15707 = ~n15706;
  assign n15705 = n15708 & n15669;
  assign n15709 = n15744 ^ n15745;
  assign n15746 = ~n15744;
  assign n15674 = ~n15764;
  assign n12158 = n15807 & n15808;
  assign n15559 = n15586 ^ n15587;
  assign n15540 = n15603 ^ n15604;
  assign n15602 = n15617 & n15618;
  assign n15590 = n15619 & n15620;
  assign n15652 = ~n15665;
  assign n11785 = n15684 ^ n15685;
  assign n15599 = ~n15694;
  assign n15667 = n15705 ^ n15706;
  assign n15695 = n15707 & n15708;
  assign n15688 = n15709 ^ n15710;
  assign n15729 = n15746 & n15747;
  assign n15730 = n15765 ^ n12158;
  assign n15748 = n12158 & n15781;
  assign n13651 = ~n12158;
  assign n14266 = n15558 ^ n15559;
  assign n15505 = n15559 & n15558;
  assign n15563 = n15590 ^ n15591;
  assign n15588 = ~n15602;
  assign n15592 = ~n15590;
  assign n15623 = n15652 & n15653;
  assign n15650 = n11785 & n15657;
  assign n11854 = ~n11785;
  assign n15622 = n15625 & n15599;
  assign n15568 = n15666 ^ n15667;
  assign n15580 = n15667 & n15666;
  assign n15672 = n15688 & n186;
  assign n15668 = ~n15695;
  assign n15670 = ~n15688;
  assign n15711 = ~n15729;
  assign n14970 = n15730 ^ n15731;
  assign n15585 = n15748 ^ n13557;
  assign n15476 = ~n14266;
  assign n15508 = ~n15505;
  assign n15541 = n15563 ^ n15564;
  assign n15560 = n15588 & n15589;
  assign n15577 = n15592 & n15593;
  assign n11832 = n15622 ^ n15623;
  assign n15624 = ~n15623;
  assign n14360 = ~n15650;
  assign n15632 = n11854 & n15651;
  assign n15621 = n11854 & n14337;
  assign n15634 = n15568 & n12979;
  assign n15633 = ~n15568;
  assign n15607 = n15668 & n15669;
  assign n15658 = n15670 & n15671;
  assign n15609 = ~n15672;
  assign n15673 = n15711 & n15712;
  assign n14978 = ~n14970;
  assign n15530 = n15541 & n393;
  assign n15528 = ~n15541;
  assign n15526 = n15560 ^ n15540;
  assign n15562 = n15560 & n15572;
  assign n15561 = ~n15560;
  assign n15565 = ~n15577;
  assign n15595 = n11832 & n14323;
  assign n15573 = n11832 & n14276;
  assign n11843 = ~n11832;
  assign n15532 = n15621 ^ n13094;
  assign n15605 = n15624 & n15625;
  assign n14385 = ~n15632;
  assign n15626 = n15633 & n13018;
  assign n15570 = ~n15634;
  assign n15635 = ~n15607;
  assign n15636 = ~n15658;
  assign n15654 = n15673 ^ n15674;
  assign n15675 = ~n15673;
  assign n15506 = n394 ^ n15526;
  assign n15522 = n15528 & n15529;
  assign n15471 = ~n15530;
  assign n15549 = n15561 & n394;
  assign n15539 = ~n15562;
  assign n15531 = n15565 & n15566;
  assign n15550 = n15573 ^ n13073;
  assign n15578 = n11843 & n15594;
  assign n14345 = ~n15595;
  assign n15597 = n15532 & n15600;
  assign n15596 = ~n15532;
  assign n15598 = ~n15605;
  assign n14382 = n14385 & n14360;
  assign n15538 = ~n15626;
  assign n15627 = n15635 & n15636;
  assign n15606 = n15636 & n15609;
  assign n15639 = n15654 & n185;
  assign n15637 = ~n15654;
  assign n15659 = n15675 & n15676;
  assign n15435 = n15505 ^ n15506;
  assign n15507 = ~n15506;
  assign n15497 = ~n15522;
  assign n15509 = n15531 ^ n15532;
  assign n15527 = n15539 & n15540;
  assign n15519 = ~n15549;
  assign n15533 = ~n15531;
  assign n15544 = n15550 & n15551;
  assign n15542 = ~n15550;
  assign n14326 = ~n15578;
  assign n15579 = n15596 & n15510;
  assign n15534 = ~n15597;
  assign n15567 = n15598 & n15599;
  assign n15581 = n15606 ^ n15607;
  assign n15608 = ~n15627;
  assign n15628 = n15637 & n15638;
  assign n15557 = ~n15639;
  assign n15640 = ~n15659;
  assign n15421 = ~n15435;
  assign n15453 = n15507 & n15508;
  assign n15498 = n15497 & n15471;
  assign n15432 = n15509 ^ n15510;
  assign n15518 = ~n15527;
  assign n15523 = n15533 & n15534;
  assign n15535 = n15542 & n15543;
  assign n15463 = ~n15544;
  assign n15536 = n15567 ^ n15568;
  assign n15514 = ~n15579;
  assign n15569 = ~n15567;
  assign n15571 = n15580 ^ n15581;
  assign n15546 = n15581 & n15580;
  assign n15574 = n15608 & n15609;
  assign n15583 = ~n15628;
  assign n15610 = n15640 & n15641;
  assign n15487 = n15432 & n392;
  assign n15456 = ~n15453;
  assign n15479 = ~n15498;
  assign n15485 = ~n15432;
  assign n15478 = n15518 & n15519;
  assign n15513 = ~n15523;
  assign n15491 = ~n15535;
  assign n11739 = n15536 ^ n13018;
  assign n15552 = n15569 & n15570;
  assign n15554 = n15571 & n12944;
  assign n15553 = ~n15571;
  assign n15582 = ~n15574;
  assign n15601 = n15583 & n15557;
  assign n15584 = n15610 ^ n15611;
  assign n15454 = n15478 ^ n15479;
  assign n15480 = n15485 & n15486;
  assign n15434 = ~n15487;
  assign n15496 = ~n15478;
  assign n15489 = n15513 & n15514;
  assign n15511 = n11739 & n14285;
  assign n15488 = n15463 & n15491;
  assign n11726 = ~n11739;
  assign n15537 = ~n15552;
  assign n15545 = n15553 & n12994;
  assign n15516 = ~n15554;
  assign n15576 = n15582 & n15583;
  assign n15555 = n15584 ^ n15585;
  assign n15575 = ~n15601;
  assign n15418 = n15453 ^ n15454;
  assign n15455 = ~n15454;
  assign n15451 = ~n15480;
  assign n15388 = n15488 ^ n15489;
  assign n15484 = n15496 & n15497;
  assign n15490 = ~n15489;
  assign n14288 = ~n15511;
  assign n15499 = n11726 & n15512;
  assign n15492 = n11726 & n14231;
  assign n15503 = n15537 & n15538;
  assign n15495 = ~n15545;
  assign n15525 = n184 ^ n15555;
  assign n15547 = n15574 ^ n15575;
  assign n15556 = ~n15576;
  assign n15401 = ~n15418;
  assign n15410 = n15455 & n15456;
  assign n15460 = n15388 & n15473;
  assign n15461 = ~n15388;
  assign n15470 = ~n15484;
  assign n15481 = n15490 & n15491;
  assign n15424 = n15492 ^ n12979;
  assign n14308 = ~n15499;
  assign n15515 = ~n15503;
  assign n15502 = n15516 & n15495;
  assign n15445 = n15546 ^ n15547;
  assign n15524 = n15556 & n15557;
  assign n15548 = ~n15547;
  assign n15413 = ~n15410;
  assign n15416 = ~n15460;
  assign n15457 = n15461 & n407;
  assign n15449 = n15470 & n15471;
  assign n15465 = n15424 & n15474;
  assign n15462 = ~n15481;
  assign n15464 = ~n15424;
  assign n11635 = n15502 ^ n15503;
  assign n15504 = n15515 & n15516;
  assign n15521 = n15445 & n12937;
  assign n15501 = n15524 ^ n15525;
  assign n15520 = ~n15445;
  assign n15500 = n15548 & n15546;
  assign n15431 = n392 ^ n15449;
  assign n15390 = ~n15457;
  assign n15450 = ~n15449;
  assign n15439 = n15462 & n15463;
  assign n15458 = n15464 & n15440;
  assign n15426 = ~n15465;
  assign n15477 = n11635 & n14266;
  assign n15466 = n11635 & n14186;
  assign n11709 = ~n11635;
  assign n15493 = n15500 ^ n15501;
  assign n15494 = ~n15504;
  assign n15517 = n15520 & n12906;
  assign n15448 = ~n15521;
  assign n15411 = n15431 ^ n15432;
  assign n15423 = n15439 ^ n15440;
  assign n15438 = n15450 & n15451;
  assign n15441 = ~n15439;
  assign n15442 = ~n15458;
  assign n15377 = n15466 ^ n12944;
  assign n15472 = n11709 & n15476;
  assign n14268 = ~n15477;
  assign n15483 = n15493 & n12893;
  assign n15467 = n15494 & n15495;
  assign n15482 = ~n15493;
  assign n15469 = ~n15517;
  assign n15365 = n15410 ^ n15411;
  assign n15412 = ~n15411;
  assign n15417 = n15423 ^ n15424;
  assign n15433 = ~n15438;
  assign n15436 = n15441 & n15442;
  assign n15444 = n15377 & n15452;
  assign n15443 = ~n15377;
  assign n15446 = n15467 ^ n12906;
  assign n14243 = ~n15472;
  assign n15475 = n15482 & n12904;
  assign n15430 = ~n15483;
  assign n15468 = ~n15467;
  assign n15348 = ~n15365;
  assign n15361 = n15412 & n15413;
  assign n15400 = n15417 & n406;
  assign n15398 = ~n15417;
  assign n15414 = n15433 & n15434;
  assign n15425 = ~n15436;
  assign n15437 = n15443 & n15404;
  assign n15379 = ~n15444;
  assign n11659 = n15445 ^ n15446;
  assign n15459 = n15468 & n15469;
  assign n15409 = ~n15475;
  assign n15364 = ~n15361;
  assign n15394 = n15398 & n15399;
  assign n15344 = ~n15400;
  assign n15387 = n407 ^ n15414;
  assign n15415 = ~n15414;
  assign n15403 = n15425 & n15426;
  assign n15422 = n11659 & n15435;
  assign n15406 = ~n15437;
  assign n11576 = ~n11659;
  assign n15427 = n15430 & n15409;
  assign n15447 = ~n15459;
  assign n15362 = n15387 ^ n15388;
  assign n15367 = ~n15394;
  assign n15376 = n15403 ^ n15404;
  assign n15397 = n15415 & n15416;
  assign n15405 = ~n15403;
  assign n15419 = n11576 & n15421;
  assign n14196 = ~n15422;
  assign n15407 = n11576 & n14095;
  assign n15428 = n15447 & n15448;
  assign n15294 = n15361 ^ n15362;
  assign n15363 = ~n15362;
  assign n15350 = n15367 & n15344;
  assign n15368 = n15376 ^ n15377;
  assign n15389 = ~n15397;
  assign n15396 = n15405 & n15406;
  assign n15391 = n15407 ^ n12906;
  assign n14220 = ~n15419;
  assign n11503 = n15427 ^ n15428;
  assign n15429 = ~n15428;
  assign n15303 = ~n15294;
  assign n15332 = n15363 & n15364;
  assign n15355 = n15368 & n405;
  assign n15353 = ~n15368;
  assign n15351 = n15389 & n15390;
  assign n15380 = n15391 & n15392;
  assign n15378 = ~n15396;
  assign n15381 = ~n15391;
  assign n14217 = n14220 & n14196;
  assign n15402 = n11503 & n15418;
  assign n15393 = n11503 & n14135;
  assign n11574 = ~n11503;
  assign n15420 = n15429 & n15430;
  assign n15333 = n15350 ^ n15351;
  assign n15346 = n15353 & n15354;
  assign n15305 = ~n15355;
  assign n15366 = ~n15351;
  assign n15335 = n15378 & n15379;
  assign n15337 = ~n15380;
  assign n15372 = n15381 & n15382;
  assign n15373 = n15393 ^ n12893;
  assign n15395 = n11574 & n15401;
  assign n14177 = ~n15402;
  assign n15408 = ~n15420;
  assign n14058 = n15332 ^ n15333;
  assign n15289 = n15333 & n15332;
  assign n15326 = ~n15346;
  assign n15352 = n15366 & n15367;
  assign n15356 = ~n15335;
  assign n15357 = ~n15372;
  assign n15371 = n15373 & n15374;
  assign n15369 = ~n15373;
  assign n14160 = ~n15395;
  assign n15383 = n15408 & n15409;
  assign n15256 = ~n14058;
  assign n15292 = ~n15289;
  assign n15309 = n15326 & n15305;
  assign n15343 = ~n15352;
  assign n15347 = n15356 & n15357;
  assign n15334 = n15357 & n15337;
  assign n15358 = n15369 & n15370;
  assign n15299 = ~n15371;
  assign n14174 = n14177 & n14160;
  assign n11516 = n15383 ^ n15384;
  assign n15385 = ~n15383;
  assign n15268 = n15334 ^ n15335;
  assign n15310 = n15343 & n15344;
  assign n15336 = ~n15347;
  assign n15317 = ~n15358;
  assign n15349 = n11516 & n15365;
  assign n11432 = ~n11516;
  assign n15375 = n15385 & n15386;
  assign n15290 = n15309 ^ n15310;
  assign n15312 = n15268 & n15327;
  assign n15313 = ~n15268;
  assign n15325 = ~n15310;
  assign n15314 = n15336 & n15337;
  assign n15338 = n15317 & n15299;
  assign n15345 = n11432 & n15348;
  assign n14120 = ~n15349;
  assign n15339 = n11432 & n14080;
  assign n15359 = ~n15375;
  assign n14024 = n15289 ^ n15290;
  assign n15291 = ~n15290;
  assign n15284 = ~n15312;
  assign n15306 = n15313 & n404;
  assign n15311 = n15325 & n15326;
  assign n15316 = ~n15314;
  assign n15315 = ~n15338;
  assign n15328 = n15339 ^ n12784;
  assign n14144 = ~n15345;
  assign n15340 = n15359 & n15360;
  assign n15231 = ~n14024;
  assign n15239 = n15291 & n15292;
  assign n15270 = ~n15306;
  assign n15304 = ~n15311;
  assign n15244 = n15314 ^ n15315;
  assign n15307 = n15316 & n15317;
  assign n15318 = n15328 & n15329;
  assign n15319 = ~n15328;
  assign n15330 = n14144 & n14120;
  assign n15321 = n15340 ^ n12830;
  assign n15341 = ~n15340;
  assign n15242 = ~n15239;
  assign n15282 = n15304 & n15305;
  assign n15297 = n15244 & n403;
  assign n15295 = ~n15244;
  assign n15298 = ~n15307;
  assign n15259 = ~n15318;
  assign n15308 = n15319 & n15320;
  assign n11342 = n15321 ^ n15322;
  assign n14142 = ~n15330;
  assign n15331 = n15341 & n15342;
  assign n15267 = n404 ^ n15282;
  assign n15283 = ~n15282;
  assign n15286 = n15295 & n15296;
  assign n15224 = ~n15297;
  assign n15271 = n15298 & n15299;
  assign n15293 = n11342 & n15303;
  assign n15276 = ~n15308;
  assign n11417 = ~n11342;
  assign n15323 = ~n15331;
  assign n15240 = n15267 ^ n15268;
  assign n15274 = n15283 & n15284;
  assign n15246 = ~n15286;
  assign n15275 = ~n15271;
  assign n14084 = ~n15293;
  assign n15285 = n11417 & n15294;
  assign n15287 = n15276 & n15259;
  assign n15277 = n11417 & n14043;
  assign n15300 = n15323 & n15324;
  assign n13984 = n15239 ^ n15240;
  assign n15241 = ~n15240;
  assign n15269 = ~n15274;
  assign n15273 = n15275 & n15276;
  assign n15214 = n15277 ^ n12838;
  assign n14102 = ~n15285;
  assign n15272 = ~n15287;
  assign n15279 = n15300 ^ n12706;
  assign n15301 = ~n15300;
  assign n15185 = ~n13984;
  assign n15204 = n15241 & n15242;
  assign n15243 = n15269 & n15270;
  assign n15262 = n15214 & n15234;
  assign n15257 = n15271 ^ n15272;
  assign n15258 = ~n15273;
  assign n15260 = ~n15214;
  assign n14099 = n14102 & n14084;
  assign n11257 = n15278 ^ n15279;
  assign n15288 = n15301 & n15302;
  assign n15222 = n15243 ^ n15244;
  assign n15245 = ~n15243;
  assign n15252 = n15257 & n402;
  assign n15233 = n15258 & n15259;
  assign n15253 = n15260 & n15261;
  assign n15236 = ~n15262;
  assign n15255 = n11257 & n14058;
  assign n15250 = ~n15257;
  assign n15248 = n11257 & n13994;
  assign n11329 = ~n11257;
  assign n15280 = ~n15288;
  assign n15205 = n403 ^ n15222;
  assign n15213 = n15233 ^ n15234;
  assign n15230 = n15245 & n15246;
  assign n15174 = n15248 ^ n12706;
  assign n15247 = n15250 & n15251;
  assign n15187 = ~n15252;
  assign n15235 = ~n15233;
  assign n15216 = ~n15253;
  assign n14060 = ~n15255;
  assign n15249 = n11329 & n15256;
  assign n15263 = n15280 & n15281;
  assign n13941 = n15204 ^ n15205;
  assign n15181 = n15205 & n15204;
  assign n15167 = n15213 ^ n15214;
  assign n15226 = n15174 & n15228;
  assign n15223 = ~n15230;
  assign n15229 = n15235 & n15236;
  assign n15225 = ~n15174;
  assign n15209 = ~n15247;
  assign n14040 = ~n15249;
  assign n11303 = n15263 ^ n15264;
  assign n15265 = ~n15263;
  assign n15153 = ~n13941;
  assign n15184 = ~n15181;
  assign n15192 = n15167 & n15210;
  assign n15193 = ~n15167;
  assign n15207 = n15223 & n15224;
  assign n15217 = n15225 & n15195;
  assign n15176 = ~n15226;
  assign n15206 = n15209 & n15187;
  assign n15215 = ~n15229;
  assign n15232 = n11303 & n14024;
  assign n11285 = ~n11303;
  assign n15254 = n15265 & n15266;
  assign n15169 = ~n15192;
  assign n15188 = n15193 & n401;
  assign n15182 = n15206 ^ n15207;
  assign n15208 = ~n15207;
  assign n15194 = n15215 & n15216;
  assign n15196 = ~n15217;
  assign n15227 = n11285 & n15231;
  assign n14005 = ~n15232;
  assign n15218 = n11285 & n13953;
  assign n15237 = ~n15254;
  assign n15105 = n15181 ^ n15182;
  assign n15147 = ~n15188;
  assign n15183 = ~n15182;
  assign n15173 = n15194 ^ n15195;
  assign n15191 = n15208 & n15209;
  assign n15197 = ~n15194;
  assign n15136 = n15218 ^ n12725;
  assign n14026 = ~n15227;
  assign n15219 = n15237 & n15238;
  assign n15122 = ~n15105;
  assign n15124 = n15173 ^ n15174;
  assign n15118 = n15183 & n15184;
  assign n15186 = ~n15191;
  assign n15189 = n15196 & n15197;
  assign n15198 = n15136 & n15211;
  assign n15199 = ~n15136;
  assign n15201 = n15219 ^ n12677;
  assign n15220 = ~n15219;
  assign n15158 = n15124 & n400;
  assign n15156 = ~n15124;
  assign n15121 = ~n15118;
  assign n15166 = n15186 & n15187;
  assign n15175 = ~n15189;
  assign n15138 = ~n15198;
  assign n15190 = n15199 & n15160;
  assign n11209 = n15200 ^ n15201;
  assign n15212 = n15220 & n15221;
  assign n15151 = n15156 & n15157;
  assign n15100 = ~n15158;
  assign n15145 = n15166 ^ n15167;
  assign n15168 = ~n15166;
  assign n15159 = n15175 & n15176;
  assign n15172 = n11209 & n15185;
  assign n15162 = ~n15190;
  assign n11089 = ~n11209;
  assign n15202 = ~n15212;
  assign n15119 = n401 ^ n15145;
  assign n15126 = ~n15151;
  assign n15135 = n15159 ^ n15160;
  assign n15155 = n15168 & n15169;
  assign n15161 = ~n15159;
  assign n15170 = n11089 & n13984;
  assign n13963 = ~n15172;
  assign n15163 = n11089 & n13858;
  assign n15178 = n15202 & n15203;
  assign n15080 = n15118 ^ n15119;
  assign n15120 = ~n15119;
  assign n15127 = n15135 ^ n15136;
  assign n15146 = ~n15155;
  assign n15152 = n15161 & n15162;
  assign n15091 = n15163 ^ n12677;
  assign n13986 = ~n15170;
  assign n11002 = n15177 ^ n15178;
  assign n15179 = ~n15178;
  assign n15063 = ~n15080;
  assign n15076 = n15120 & n15121;
  assign n15110 = n15127 & n415;
  assign n15108 = ~n15127;
  assign n15123 = n15146 & n15147;
  assign n15140 = n15091 & n15148;
  assign n15137 = ~n15152;
  assign n15139 = ~n15091;
  assign n15154 = n11002 & n13941;
  assign n15149 = n11002 & n13868;
  assign n11126 = ~n11002;
  assign n15171 = n15179 & n15180;
  assign n15079 = ~n15076;
  assign n15103 = n15108 & n15109;
  assign n15055 = ~n15110;
  assign n15098 = n15123 ^ n15124;
  assign n15125 = ~n15123;
  assign n15111 = n15137 & n15138;
  assign n15133 = n15139 & n15112;
  assign n15093 = ~n15140;
  assign n15131 = n15149 ^ n12574;
  assign n15150 = n11126 & n15153;
  assign n13943 = ~n15154;
  assign n15164 = ~n15171;
  assign n15077 = n400 ^ n15098;
  assign n15082 = ~n15103;
  assign n15090 = n15111 ^ n15112;
  assign n15107 = n15125 & n15126;
  assign n15113 = ~n15111;
  assign n15128 = n15131 & n15132;
  assign n15114 = ~n15133;
  assign n15129 = ~n15131;
  assign n13925 = ~n15150;
  assign n15142 = n15164 & n15165;
  assign n15019 = n15076 ^ n15077;
  assign n15078 = ~n15077;
  assign n15087 = n15082 & n15055;
  assign n15083 = n15090 ^ n15091;
  assign n15099 = ~n15107;
  assign n15104 = n15113 & n15114;
  assign n15049 = ~n15128;
  assign n15115 = n15129 & n15130;
  assign n11041 = n15141 ^ n15142;
  assign n15143 = ~n15142;
  assign n15009 = ~n15019;
  assign n15038 = n15078 & n15079;
  assign n15068 = n15083 & n414;
  assign n15060 = ~n15087;
  assign n15066 = ~n15083;
  assign n15059 = n15099 & n15100;
  assign n15092 = ~n15104;
  assign n15072 = ~n15115;
  assign n15106 = n11041 & n15122;
  assign n15101 = n11041 & n13847;
  assign n11052 = ~n11041;
  assign n15134 = n15143 & n15144;
  assign n15039 = n15059 ^ n15060;
  assign n15041 = ~n15038;
  assign n15061 = n15066 & n15067;
  assign n15021 = ~n15068;
  assign n15081 = ~n15059;
  assign n15070 = n15092 & n15093;
  assign n15069 = n15072 & n15049;
  assign n15011 = n15101 ^ n12506;
  assign n15102 = n11052 & n15105;
  assign n13907 = ~n15106;
  assign n15116 = ~n15134;
  assign n14998 = n15038 ^ n15039;
  assign n15040 = ~n15039;
  assign n15035 = ~n15061;
  assign n15000 = n15069 ^ n15070;
  assign n15065 = n15081 & n15082;
  assign n15071 = ~n15070;
  assign n15084 = n15011 & n15088;
  assign n15085 = ~n15011;
  assign n13885 = ~n15102;
  assign n15095 = n15116 & n15117;
  assign n14984 = ~n14998;
  assign n14903 = n15040 & n15041;
  assign n15042 = n15035 & n15021;
  assign n15046 = n15000 & n15056;
  assign n15047 = ~n15000;
  assign n15054 = ~n15065;
  assign n15062 = n15071 & n15072;
  assign n15014 = ~n15084;
  assign n15073 = n15085 & n15027;
  assign n15086 = n13907 & n13885;
  assign n10934 = n15094 ^ n15095;
  assign n15096 = ~n15095;
  assign n15008 = ~n14903;
  assign n15023 = ~n15042;
  assign n15002 = ~n15046;
  assign n15043 = n15047 & n413;
  assign n15022 = n15054 & n15055;
  assign n15048 = ~n15062;
  assign n15029 = ~n15073;
  assign n15064 = n10934 & n15080;
  assign n15057 = n10934 & n13803;
  assign n13905 = ~n15086;
  assign n10957 = ~n10934;
  assign n15089 = n15096 & n15097;
  assign n14922 = n15022 ^ n15023;
  assign n14974 = ~n15043;
  assign n15034 = ~n15022;
  assign n15026 = n15048 & n15049;
  assign n14964 = n15057 ^ n12448;
  assign n15058 = n10957 & n15063;
  assign n13867 = ~n15064;
  assign n15074 = ~n15089;
  assign n14951 = n14922 & n15008;
  assign n15012 = n15026 ^ n15027;
  assign n15025 = n15034 & n15035;
  assign n15028 = ~n15026;
  assign n15036 = n14964 & n15044;
  assign n15037 = ~n14964;
  assign n13844 = ~n15058;
  assign n15050 = n15074 & n15075;
  assign n14954 = ~n14951;
  assign n15003 = n15011 ^ n15012;
  assign n15020 = ~n15025;
  assign n15024 = n15028 & n15029;
  assign n14966 = ~n15036;
  assign n15030 = n15037 & n14991;
  assign n13864 = n13867 & n13844;
  assign n15031 = n15050 ^ n15051;
  assign n15052 = ~n15050;
  assign n14989 = n15003 & n412;
  assign n14987 = ~n15003;
  assign n14999 = n15020 & n15021;
  assign n15013 = ~n15024;
  assign n14993 = ~n15030;
  assign n10863 = n15031 ^ n12240;
  assign n15045 = n15052 & n15053;
  assign n14981 = n14987 & n14988;
  assign n14934 = ~n14989;
  assign n14972 = n14999 ^ n15000;
  assign n15001 = ~n14999;
  assign n14990 = n15013 & n15014;
  assign n15010 = n10863 & n15019;
  assign n10843 = ~n10863;
  assign n15032 = ~n15045;
  assign n14952 = n413 ^ n14972;
  assign n14956 = ~n14981;
  assign n14963 = n14990 ^ n14991;
  assign n14986 = n15001 & n15002;
  assign n14992 = ~n14990;
  assign n15006 = n10843 & n15009;
  assign n13783 = ~n15010;
  assign n14994 = n10843 & n13729;
  assign n15016 = n15032 & n15033;
  assign n13869 = n14951 ^ n14952;
  assign n14953 = ~n14952;
  assign n14938 = n14956 & n14934;
  assign n14957 = n14963 ^ n14964;
  assign n14973 = ~n14986;
  assign n14982 = n14992 & n14993;
  assign n14945 = n14994 ^ n12240;
  assign n13817 = ~n15006;
  assign n10742 = n15015 ^ n15016;
  assign n15018 = n15016 & n14996;
  assign n15017 = ~n15016;
  assign n13808 = n14931 ^ n13869;
  assign n13809 = n13869 ^ n12791;
  assign n14932 = ~n13869;
  assign n14923 = n14953 & n14954;
  assign n14943 = n14957 & n411;
  assign n14941 = ~n14957;
  assign n14939 = n14973 & n14974;
  assign n14967 = n14945 & n14975;
  assign n14965 = ~n14982;
  assign n14968 = ~n14945;
  assign n14979 = n13817 & n13783;
  assign n14985 = n10742 & n14998;
  assign n14976 = n10742 & n13689;
  assign n10749 = ~n10742;
  assign n15007 = n15017 & n15005;
  assign n15004 = ~n15018;
  assign n14896 = n13809 & n13785;
  assign n11790 = ~n13809;
  assign n14869 = n14932 & n12791;
  assign n14926 = ~n14923;
  assign n14924 = n14938 ^ n14939;
  assign n14936 = n14941 & n14942;
  assign n14893 = ~n14943;
  assign n14955 = ~n14939;
  assign n14944 = n14965 & n14966;
  assign n14947 = ~n14967;
  assign n14961 = n14968 & n14928;
  assign n14889 = n14976 ^ n12260;
  assign n13815 = ~n14979;
  assign n14980 = n10749 & n14984;
  assign n13738 = ~n14985;
  assign n14997 = n15004 & n15005;
  assign n14995 = ~n15007;
  assign n14885 = n14896 ^ n14897;
  assign n14880 = n14896 ^ n14898;
  assign n14916 = n14923 ^ n14924;
  assign n14925 = ~n14924;
  assign n14918 = ~n14936;
  assign n14927 = n14944 ^ n14945;
  assign n14940 = n14955 & n14956;
  assign n14946 = ~n14944;
  assign n14960 = n14889 & n14913;
  assign n14930 = ~n14961;
  assign n14958 = ~n14889;
  assign n13731 = ~n14980;
  assign n14983 = n14995 & n14996;
  assign n14977 = ~n14997;
  assign n14575 = n103 ^ n14880;
  assign n14780 = n14880 & n103;
  assign n14863 = n14885 & n14886;
  assign n14907 = n14916 & n12711;
  assign n14906 = ~n14916;
  assign n14882 = n14925 & n14926;
  assign n14921 = n14918 & n14893;
  assign n14919 = n14927 ^ n14928;
  assign n14933 = ~n14940;
  assign n14937 = n14946 & n14947;
  assign n14948 = n14958 & n14959;
  assign n14891 = ~n14960;
  assign n13753 = n13738 & n13731;
  assign n14971 = n14977 & n14978;
  assign n14969 = ~n14983;
  assign n14825 = n14863 ^ n14864;
  assign n14867 = n14863 & n14864;
  assign n14570 = ~n14575;
  assign n14865 = ~n14863;
  assign n14899 = n14906 & n12700;
  assign n14871 = ~n14907;
  assign n14911 = n14919 & n410;
  assign n14901 = ~n14921;
  assign n14909 = ~n14919;
  assign n14900 = n14933 & n14934;
  assign n14929 = ~n14937;
  assign n14915 = ~n14948;
  assign n14962 = n14969 & n14970;
  assign n14950 = ~n14971;
  assign n14857 = n14865 & n14866;
  assign n14815 = ~n14867;
  assign n14887 = ~n14899;
  assign n14883 = n14900 ^ n14901;
  assign n14902 = n14909 & n14910;
  assign n14856 = ~n14911;
  assign n14917 = ~n14900;
  assign n14912 = n14929 & n14930;
  assign n14949 = ~n14962;
  assign n14828 = ~n14857;
  assign n14838 = n14882 ^ n14883;
  assign n14881 = n14887 & n14869;
  assign n14868 = n14887 & n14871;
  assign n14849 = n14883 & n14882;
  assign n14878 = ~n14902;
  assign n14888 = n14912 ^ n14913;
  assign n14908 = n14917 & n14918;
  assign n14914 = ~n14912;
  assign n10610 = n14949 & n14950;
  assign n11759 = n14868 ^ n14869;
  assign n14858 = n14838 & n12613;
  assign n14859 = ~n14838;
  assign n14870 = ~n14881;
  assign n14852 = ~n14849;
  assign n14884 = n14878 & n14856;
  assign n14830 = n14888 ^ n14889;
  assign n14892 = ~n14908;
  assign n14905 = n14914 & n14915;
  assign n14920 = n10610 & n14935;
  assign n12228 = ~n10610;
  assign n11761 = ~n11759;
  assign n14835 = ~n14858;
  assign n14854 = n14859 & n12565;
  assign n14853 = n14870 & n14871;
  assign n14873 = n14830 & n14879;
  assign n14861 = ~n14884;
  assign n14874 = ~n14830;
  assign n14860 = n14892 & n14893;
  assign n14890 = ~n14905;
  assign n14894 = n14920 ^ n12158;
  assign n14904 = n14922 ^ n12228;
  assign n14840 = n11761 & n13692;
  assign n14839 = n14853 ^ n12565;
  assign n14847 = ~n14854;
  assign n14848 = ~n14853;
  assign n14850 = n14860 ^ n14861;
  assign n14846 = ~n14873;
  assign n14862 = n14874 & n409;
  assign n14877 = ~n14860;
  assign n14875 = n14890 & n14891;
  assign n14876 = n14894 ^ n14895;
  assign n13701 = n14903 ^ n14904;
  assign n11617 = n14838 ^ n14839;
  assign n14826 = n14840 ^ n12700;
  assign n14843 = n14847 & n14848;
  assign n14841 = n14849 ^ n14850;
  assign n14851 = ~n14850;
  assign n14833 = ~n14862;
  assign n14822 = n14875 ^ n14876;
  assign n14872 = n14877 & n14878;
  assign n13709 = ~n13701;
  assign n14813 = n14825 ^ n14826;
  assign n14827 = n14828 & n14826;
  assign n11611 = ~n11617;
  assign n14836 = n14841 & n12551;
  assign n14834 = ~n14843;
  assign n14837 = ~n14841;
  assign n14816 = n14851 & n14852;
  assign n14855 = ~n14872;
  assign n14811 = n14813 & n102;
  assign n14809 = ~n14813;
  assign n14814 = ~n14827;
  assign n14812 = n11611 & n13626;
  assign n14804 = n14834 & n14835;
  assign n14823 = ~n14836;
  assign n14831 = n14837 & n12568;
  assign n14844 = n14855 & n14856;
  assign n14806 = n14809 & n14810;
  assign n14784 = ~n14811;
  assign n14798 = n14812 ^ n12565;
  assign n14763 = n14814 & n14815;
  assign n14824 = ~n14804;
  assign n14808 = ~n14831;
  assign n14829 = n409 ^ n14844;
  assign n14845 = ~n14844;
  assign n14794 = n14798 & n14799;
  assign n14793 = ~n14806;
  assign n14795 = ~n14798;
  assign n14782 = ~n14763;
  assign n14818 = n14823 & n14824;
  assign n14820 = n14823 & n14808;
  assign n14817 = n14829 ^ n14830;
  assign n14842 = n14845 & n14846;
  assign n14791 = n14793 & n14780;
  assign n14779 = n14793 & n14784;
  assign n14768 = ~n14794;
  assign n14792 = n14795 & n14796;
  assign n14790 = n14816 ^ n14817;
  assign n14807 = ~n14818;
  assign n14805 = ~n14820;
  assign n14819 = ~n14817;
  assign n14832 = ~n14842;
  assign n14524 = n14779 ^ n14780;
  assign n14783 = ~n14791;
  assign n14781 = ~n14792;
  assign n11471 = n14804 ^ n14805;
  assign n14800 = n14790 & n12381;
  assign n14802 = n14807 & n14808;
  assign n14801 = ~n14790;
  assign n14788 = n14819 & n14816;
  assign n14821 = n14832 & n14833;
  assign n14526 = ~n14524;
  assign n14776 = n14781 & n14782;
  assign n14712 = n14783 & n14784;
  assign n14777 = n14781 & n14768;
  assign n11545 = ~n11471;
  assign n14772 = ~n14800;
  assign n14797 = n14801 & n12437;
  assign n14787 = ~n14802;
  assign n14803 = n14821 ^ n14822;
  assign n14767 = ~n14776;
  assign n14738 = ~n14712;
  assign n14764 = ~n14777;
  assign n14770 = n14787 ^ n14790;
  assign n14775 = n11545 & n13571;
  assign n14786 = ~n14797;
  assign n14789 = n408 ^ n14803;
  assign n14755 = n14763 ^ n14764;
  assign n14725 = n14767 & n14768;
  assign n11441 = n14770 ^ n12437;
  assign n14765 = n14775 ^ n12551;
  assign n14785 = n14786 & n14787;
  assign n14778 = n14788 ^ n14789;
  assign n14753 = n14755 & n101;
  assign n14751 = ~n14755;
  assign n14746 = ~n14725;
  assign n14754 = n11441 & n13534;
  assign n14760 = n14765 & n14766;
  assign n11463 = ~n11441;
  assign n14761 = ~n14765;
  assign n14773 = n14778 & n12265;
  assign n14771 = ~n14785;
  assign n14774 = ~n14778;
  assign n14744 = n14751 & n14752;
  assign n14723 = ~n14753;
  assign n14715 = n14754 ^ n12381;
  assign n14731 = ~n14760;
  assign n14757 = n14761 & n14762;
  assign n14748 = n14771 & n14772;
  assign n14750 = ~n14773;
  assign n14769 = n14774 & n12386;
  assign n14740 = n14715 & n14741;
  assign n14737 = ~n14744;
  assign n14739 = ~n14715;
  assign n14745 = ~n14757;
  assign n14758 = ~n14748;
  assign n14759 = ~n14769;
  assign n14728 = n14737 & n14738;
  assign n14729 = n14737 & n14723;
  assign n14732 = n14739 & n14694;
  assign n14716 = ~n14740;
  assign n14742 = n14745 & n14746;
  assign n14743 = n14745 & n14731;
  assign n14756 = n14758 & n14759;
  assign n14747 = n14759 & n14750;
  assign n14722 = ~n14728;
  assign n14713 = ~n14729;
  assign n14696 = ~n14732;
  assign n14730 = ~n14742;
  assign n14726 = ~n14743;
  assign n11392 = n14747 ^ n14748;
  assign n14749 = ~n14756;
  assign n14692 = n14712 ^ n14713;
  assign n14669 = n14722 & n14723;
  assign n14718 = n14725 ^ n14726;
  assign n14714 = n14730 & n14731;
  assign n14724 = n11392 & n13496;
  assign n11403 = ~n11392;
  assign n14733 = n14749 & n14750;
  assign n14481 = n14692 ^ n14524;
  assign n14647 = n14692 & n14524;
  assign n14690 = ~n14669;
  assign n14693 = n14714 ^ n14715;
  assign n14711 = n14718 & n100;
  assign n14706 = n14724 ^ n12386;
  assign n14709 = ~n14718;
  assign n14717 = ~n14714;
  assign n14719 = n14733 ^ n14734;
  assign n14735 = ~n14733;
  assign n14494 = ~n14481;
  assign n14685 = n14693 ^ n14694;
  assign n14702 = n14706 & n14707;
  assign n14705 = n14709 & n14710;
  assign n14675 = ~n14711;
  assign n14708 = n14716 & n14717;
  assign n11296 = n14719 ^ n12297;
  assign n14703 = ~n14706;
  assign n14727 = n14735 & n14736;
  assign n14679 = n14685 & n99;
  assign n14677 = ~n14685;
  assign n14686 = n11296 & n13458;
  assign n14660 = ~n14702;
  assign n14697 = n14703 & n14704;
  assign n14689 = ~n14705;
  assign n14695 = ~n14708;
  assign n11310 = ~n11296;
  assign n14720 = ~n14727;
  assign n14671 = n14677 & n14678;
  assign n14634 = ~n14679;
  assign n14672 = n14686 ^ n12297;
  assign n14687 = n14689 & n14690;
  assign n14688 = n14689 & n14675;
  assign n14657 = n14695 & n14696;
  assign n14681 = ~n14697;
  assign n14699 = n14720 & n14721;
  assign n14651 = ~n14671;
  assign n14667 = n14672 & n14673;
  assign n14665 = ~n14672;
  assign n14674 = ~n14687;
  assign n14682 = n14681 & n14660;
  assign n14670 = ~n14688;
  assign n14680 = ~n14657;
  assign n11108 = n14698 ^ n14699;
  assign n14700 = ~n14699;
  assign n14653 = n14651 & n14634;
  assign n14656 = n14665 & n14666;
  assign n14625 = ~n14667;
  assign n14648 = n14669 ^ n14670;
  assign n14631 = n14674 & n14675;
  assign n14676 = n14680 & n14681;
  assign n14658 = ~n14682;
  assign n14668 = n11108 & n13397;
  assign n11218 = ~n11108;
  assign n14691 = n14700 & n14701;
  assign n13226 = n14647 ^ n14648;
  assign n14632 = ~n14653;
  assign n14614 = n14648 & n14647;
  assign n14637 = ~n14656;
  assign n14593 = n14657 ^ n14658;
  assign n14652 = ~n14631;
  assign n14585 = n14668 ^ n12235;
  assign n14659 = ~n14676;
  assign n14683 = ~n14691;
  assign n14615 = n14631 ^ n14632;
  assign n14428 = ~n13226;
  assign n14641 = n14637 & n14625;
  assign n14642 = n14593 & n98;
  assign n14617 = ~n14614;
  assign n14646 = n14651 & n14652;
  assign n14649 = n14585 & n14654;
  assign n14639 = ~n14593;
  assign n14622 = n14659 & n14660;
  assign n14650 = ~n14585;
  assign n14661 = n14683 & n14684;
  assign n14409 = n14614 ^ n14615;
  assign n14616 = ~n14615;
  assign n14636 = n14639 & n14640;
  assign n14623 = ~n14641;
  assign n14595 = ~n14642;
  assign n14633 = ~n14646;
  assign n14587 = ~n14649;
  assign n14643 = n14650 & n14603;
  assign n14638 = ~n14622;
  assign n11132 = n14661 ^ n14662;
  assign n14663 = ~n14661;
  assign n14404 = ~n14409;
  assign n14576 = n14616 & n14617;
  assign n14611 = n14622 ^ n14623;
  assign n14618 = n14633 & n14634;
  assign n14620 = ~n14636;
  assign n14635 = n14637 & n14638;
  assign n14605 = ~n14643;
  assign n11115 = ~n11132;
  assign n14655 = n14663 & n14664;
  assign n14579 = ~n14576;
  assign n14601 = n14611 & n97;
  assign n14592 = n98 ^ n14618;
  assign n14599 = ~n14611;
  assign n14619 = ~n14618;
  assign n14624 = ~n14635;
  assign n14626 = n11115 & n13360;
  assign n14644 = ~n14655;
  assign n14577 = n14592 ^ n14593;
  assign n14596 = n14599 & n14600;
  assign n14557 = ~n14601;
  assign n14612 = n14619 & n14620;
  assign n14602 = n14624 & n14625;
  assign n14540 = n14626 ^ n12110;
  assign n14627 = n14644 & n14645;
  assign n13154 = n14576 ^ n14577;
  assign n14578 = ~n14577;
  assign n14580 = ~n14596;
  assign n14584 = n14602 ^ n14603;
  assign n14594 = ~n14612;
  assign n14606 = n14540 & n14613;
  assign n14604 = ~n14602;
  assign n14607 = ~n14540;
  assign n14608 = n14627 ^ n14628;
  assign n14629 = ~n14627;
  assign n14364 = ~n13154;
  assign n14530 = n14578 & n14579;
  assign n14534 = n14584 ^ n14585;
  assign n14582 = n14580 & n14557;
  assign n14554 = n14594 & n14595;
  assign n14597 = n14604 & n14605;
  assign n14542 = ~n14606;
  assign n14598 = n14607 & n14566;
  assign n11045 = n12094 ^ n14608;
  assign n14621 = n14629 & n14630;
  assign n14564 = n14534 & n96;
  assign n14562 = ~n14534;
  assign n14555 = ~n14582;
  assign n14581 = ~n14554;
  assign n14574 = n11045 & n13327;
  assign n14586 = ~n14597;
  assign n14568 = ~n14598;
  assign n11063 = ~n11045;
  assign n14609 = ~n14621;
  assign n14535 = n14554 ^ n14555;
  assign n14553 = n14562 & n14563;
  assign n14511 = ~n14564;
  assign n14558 = n14574 ^ n12094;
  assign n14573 = n14580 & n14581;
  assign n14565 = n14586 & n14587;
  assign n14588 = n14609 & n14610;
  assign n14305 = n14530 ^ n14535;
  assign n14485 = n14535 & n14530;
  assign n14531 = ~n14535;
  assign n14536 = ~n14553;
  assign n14550 = n14558 & n14559;
  assign n14539 = n14565 ^ n14566;
  assign n14551 = ~n14558;
  assign n14556 = ~n14573;
  assign n14567 = ~n14565;
  assign n10973 = n14588 ^ n14589;
  assign n14590 = ~n14588;
  assign n14309 = n14530 ^ n14531;
  assign n14488 = ~n14485;
  assign n14529 = n14539 ^ n14540;
  assign n14501 = ~n14550;
  assign n14543 = n14551 & n14552;
  assign n14549 = n14556 & n14557;
  assign n14560 = n14567 & n14568;
  assign n14569 = n10973 & n14575;
  assign n10961 = ~n10973;
  assign n14583 = n14590 & n14591;
  assign n14518 = n14529 & n111;
  assign n14516 = ~n14529;
  assign n14519 = ~n14543;
  assign n14533 = ~n14549;
  assign n14541 = ~n14560;
  assign n14544 = n10961 & n13303;
  assign n13338 = ~n14569;
  assign n14561 = n10961 & n14570;
  assign n14571 = ~n14583;
  assign n14512 = n14516 & n14517;
  assign n14470 = ~n14518;
  assign n14506 = n14533 ^ n14534;
  assign n14507 = n14519 & n14501;
  assign n14532 = n14536 & n14533;
  assign n14508 = n14541 & n14542;
  assign n14461 = n14544 ^ n12051;
  assign n13353 = ~n14561;
  assign n14546 = n14571 & n14572;
  assign n14486 = n96 ^ n14506;
  assign n14450 = n14507 ^ n14508;
  assign n14496 = ~n14512;
  assign n14510 = ~n14532;
  assign n14521 = n14461 & n14477;
  assign n14520 = ~n14508;
  assign n14522 = ~n14461;
  assign n14537 = n13353 & n13338;
  assign n10867 = n14545 ^ n14546;
  assign n14547 = ~n14546;
  assign n13066 = n14485 ^ n14486;
  assign n14490 = n14450 & n14497;
  assign n14473 = n14496 & n14470;
  assign n14487 = ~n14486;
  assign n14491 = ~n14450;
  assign n14474 = n14510 & n14511;
  assign n14513 = n14519 & n14520;
  assign n14479 = ~n14521;
  assign n14514 = n14522 & n14523;
  assign n13324 = n14524 ^ n10867;
  assign n14509 = n10867 & n13277;
  assign n14525 = n10867 & n14524;
  assign n13351 = ~n14537;
  assign n10882 = ~n10867;
  assign n14538 = n14547 & n14548;
  assign n14264 = ~n13066;
  assign n14457 = n14473 ^ n14474;
  assign n14456 = n14487 & n14488;
  assign n14452 = ~n14490;
  assign n14475 = n14491 & n110;
  assign n14495 = ~n14474;
  assign n14419 = n14509 ^ n12000;
  assign n14500 = ~n14513;
  assign n14463 = ~n14514;
  assign n13326 = ~n14525;
  assign n14515 = n10882 & n14526;
  assign n14527 = ~n14538;
  assign n14229 = n14456 ^ n14457;
  assign n14458 = ~n14457;
  assign n14459 = ~n14456;
  assign n14431 = ~n14475;
  assign n14489 = n14495 & n14496;
  assign n14493 = n14419 & n14498;
  assign n14476 = n14500 & n14501;
  assign n14492 = ~n14419;
  assign n13306 = ~n14515;
  assign n14503 = n14527 & n14528;
  assign n14215 = ~n14229;
  assign n14410 = n14458 & n14459;
  assign n14460 = n14476 ^ n14477;
  assign n14469 = ~n14489;
  assign n14480 = n14492 & n14437;
  assign n14421 = ~n14493;
  assign n14478 = ~n14476;
  assign n10726 = n14502 ^ n14503;
  assign n14504 = ~n14503;
  assign n14413 = n14460 ^ n14461;
  assign n14449 = n14469 & n14470;
  assign n14471 = n14478 & n14479;
  assign n14439 = ~n14480;
  assign n14468 = n10726 & n13239;
  assign n14482 = n10726 & n14494;
  assign n10728 = ~n10726;
  assign n14499 = n14504 & n14505;
  assign n14434 = n14413 & n14444;
  assign n14429 = n14449 ^ n14450;
  assign n14435 = ~n14413;
  assign n14451 = ~n14449;
  assign n14453 = n14468 ^ n11939;
  assign n14462 = ~n14471;
  assign n14472 = n10728 & n14481;
  assign n13285 = ~n14482;
  assign n14483 = ~n14499;
  assign n14411 = n110 ^ n14429;
  assign n14414 = ~n14434;
  assign n14432 = n14435 & n109;
  assign n14445 = n14451 & n14452;
  assign n14448 = n14453 & n14454;
  assign n14436 = n14462 & n14463;
  assign n14446 = ~n14453;
  assign n13266 = ~n14472;
  assign n14464 = n14483 & n14484;
  assign n12989 = n14410 ^ n14411;
  assign n14365 = n14411 & n14410;
  assign n14391 = ~n14432;
  assign n14418 = n14436 ^ n14437;
  assign n14430 = ~n14445;
  assign n14440 = n14446 & n14447;
  assign n14380 = ~n14448;
  assign n14438 = ~n14436;
  assign n13282 = n13285 & n13266;
  assign n14441 = n14464 ^ n14465;
  assign n14466 = ~n14464;
  assign n14205 = ~n12989;
  assign n14368 = ~n14365;
  assign n14348 = n14418 ^ n14419;
  assign n14412 = n14430 & n14431;
  assign n14433 = n14438 & n14439;
  assign n14402 = ~n14440;
  assign n10697 = n14441 ^ n11931;
  assign n14455 = n14466 & n14467;
  assign n14398 = n14348 & n108;
  assign n14389 = n14412 ^ n14413;
  assign n14396 = ~n14348;
  assign n14415 = ~n14412;
  assign n14422 = n14402 & n14380;
  assign n14408 = n10697 & n13178;
  assign n14423 = n10697 & n14428;
  assign n14420 = ~n14433;
  assign n10712 = ~n10697;
  assign n14442 = ~n14455;
  assign n14366 = n109 ^ n14389;
  assign n14392 = n14396 & n14397;
  assign n14350 = ~n14398;
  assign n14354 = n14408 ^ n11936;
  assign n14407 = n14414 & n14415;
  assign n14399 = n14420 & n14421;
  assign n14400 = ~n14422;
  assign n13248 = ~n14423;
  assign n14416 = n10712 & n13226;
  assign n14425 = n14442 & n14443;
  assign n12970 = n14365 ^ n14366;
  assign n14367 = ~n14366;
  assign n14371 = ~n14392;
  assign n14387 = n14354 & n14393;
  assign n14334 = n14399 ^ n14400;
  assign n14386 = ~n14354;
  assign n14390 = ~n14407;
  assign n14401 = ~n14399;
  assign n13229 = ~n14416;
  assign n10619 = n14424 ^ n14425;
  assign n14426 = ~n14425;
  assign n14158 = ~n12970;
  assign n14331 = n14367 & n14368;
  assign n14378 = n14334 & n107;
  assign n14381 = n14386 & n14340;
  assign n14355 = ~n14387;
  assign n14369 = n14390 & n14391;
  assign n14376 = ~n14334;
  assign n14394 = n14401 & n14402;
  assign n14388 = n10619 & n13160;
  assign n14403 = n10619 & n14409;
  assign n10626 = ~n10619;
  assign n14417 = n14426 & n14427;
  assign n14347 = n108 ^ n14369;
  assign n14372 = n14376 & n14377;
  assign n14312 = ~n14378;
  assign n14342 = ~n14381;
  assign n14370 = ~n14369;
  assign n14301 = n14388 ^ n11862;
  assign n14379 = ~n14394;
  assign n13207 = ~n14403;
  assign n14395 = n10626 & n14404;
  assign n14405 = ~n14417;
  assign n14332 = n14347 ^ n14348;
  assign n14361 = n14370 & n14371;
  assign n14336 = ~n14372;
  assign n14363 = n14301 & n14373;
  assign n14353 = n14379 & n14380;
  assign n14362 = ~n14301;
  assign n13192 = ~n14395;
  assign n14383 = n14405 & n14406;
  assign n12933 = n14331 ^ n14332;
  assign n14298 = n14332 & n14331;
  assign n14339 = n14353 ^ n14354;
  assign n14349 = ~n14361;
  assign n14357 = n14362 & n14319;
  assign n14303 = ~n14363;
  assign n14356 = ~n14353;
  assign n14374 = n13207 & n13192;
  assign n10546 = n14382 ^ n14383;
  assign n14384 = ~n14383;
  assign n14126 = ~n12933;
  assign n14292 = ~n14298;
  assign n14327 = n14339 ^ n14340;
  assign n14333 = n14349 & n14350;
  assign n14351 = n14355 & n14356;
  assign n14321 = ~n14357;
  assign n14346 = n10546 & n13094;
  assign n14358 = n10546 & n14364;
  assign n13205 = ~n14374;
  assign n10559 = ~n10546;
  assign n14375 = n14384 & n14385;
  assign n14317 = n14327 & n106;
  assign n14310 = n14333 ^ n14334;
  assign n14315 = ~n14327;
  assign n14335 = ~n14333;
  assign n14258 = n14346 ^ n11854;
  assign n14341 = ~n14351;
  assign n13177 = ~n14358;
  assign n14352 = n10559 & n13154;
  assign n14359 = ~n14375;
  assign n14299 = n107 ^ n14310;
  assign n14313 = n14315 & n14316;
  assign n14274 = ~n14317;
  assign n14328 = n14335 & n14336;
  assign n14329 = n14258 & n14337;
  assign n14318 = n14341 & n14342;
  assign n14330 = ~n14258;
  assign n13157 = ~n14352;
  assign n14343 = n14359 & n14360;
  assign n14081 = n14298 ^ n14299;
  assign n14291 = ~n14299;
  assign n14294 = ~n14313;
  assign n14300 = n14318 ^ n14319;
  assign n14311 = ~n14328;
  assign n14261 = ~n14329;
  assign n14322 = n14330 & n14282;
  assign n14320 = ~n14318;
  assign n14324 = n14343 ^ n11832;
  assign n14344 = ~n14343;
  assign n14087 = ~n14081;
  assign n14252 = n14291 & n14292;
  assign n14295 = n14294 & n14274;
  assign n14255 = n14300 ^ n14301;
  assign n14271 = n14311 & n14312;
  assign n14314 = n14320 & n14321;
  assign n14284 = ~n14322;
  assign n10531 = n14323 ^ n14324;
  assign n14338 = n14344 & n14345;
  assign n14280 = n14255 & n105;
  assign n14272 = ~n14295;
  assign n14278 = ~n14255;
  assign n14293 = ~n14271;
  assign n14290 = n10531 & n13080;
  assign n14304 = n10531 & n14309;
  assign n14302 = ~n14314;
  assign n10539 = ~n10531;
  assign n14325 = ~n14338;
  assign n14253 = n14271 ^ n14272;
  assign n14275 = n14278 & n14279;
  assign n14235 = ~n14280;
  assign n14238 = n14290 ^ n11832;
  assign n14289 = n14293 & n14294;
  assign n14281 = n14302 & n14303;
  assign n13134 = ~n14304;
  assign n14296 = n10539 & n14305;
  assign n14306 = n14325 & n14326;
  assign n14022 = n14252 ^ n14253;
  assign n14206 = n14253 & n14252;
  assign n14256 = ~n14275;
  assign n14270 = n14238 & n14276;
  assign n14259 = n14281 ^ n14282;
  assign n14269 = ~n14238;
  assign n14273 = ~n14289;
  assign n14283 = ~n14281;
  assign n13115 = ~n14296;
  assign n14286 = n14306 ^ n11739;
  assign n14307 = ~n14306;
  assign n14027 = ~n14022;
  assign n14221 = ~n14206;
  assign n14248 = n14258 ^ n14259;
  assign n14262 = n14269 & n14223;
  assign n14225 = ~n14270;
  assign n14254 = n14273 & n14274;
  assign n14277 = n14283 & n14284;
  assign n13131 = n13134 & n13115;
  assign n10461 = n14285 ^ n14286;
  assign n14297 = n14307 & n14308;
  assign n14246 = n14248 & n104;
  assign n14244 = ~n14248;
  assign n14233 = n14254 ^ n14255;
  assign n14240 = ~n14262;
  assign n14257 = ~n14254;
  assign n14247 = n10461 & n13018;
  assign n14263 = n10461 & n13066;
  assign n14260 = ~n14277;
  assign n10420 = ~n10461;
  assign n14287 = ~n14297;
  assign n14211 = n105 ^ n14233;
  assign n14236 = n14244 & n14245;
  assign n14191 = ~n14246;
  assign n14230 = n14247 ^ n11726;
  assign n14249 = n14256 & n14257;
  assign n14237 = n14260 & n14261;
  assign n13091 = ~n14263;
  assign n14250 = n10420 & n14264;
  assign n14265 = n14287 & n14288;
  assign n13982 = n14206 ^ n14211;
  assign n14178 = n14211 & n14221;
  assign n14207 = ~n14211;
  assign n14228 = n14230 & n14231;
  assign n14213 = ~n14236;
  assign n14222 = n14237 ^ n14238;
  assign n14226 = ~n14230;
  assign n14234 = ~n14249;
  assign n14239 = ~n14237;
  assign n13069 = ~n14250;
  assign n14241 = n14265 ^ n14266;
  assign n14267 = ~n14265;
  assign n13989 = n14206 ^ n14207;
  assign n14197 = n14213 & n14191;
  assign n14168 = n14222 ^ n14223;
  assign n14214 = n14226 & n14227;
  assign n14181 = ~n14228;
  assign n14198 = n14234 & n14235;
  assign n14232 = n14239 & n14240;
  assign n10401 = n14241 ^ n11709;
  assign n14251 = n14267 & n14268;
  assign n14179 = n14197 ^ n14198;
  assign n14201 = n14168 & n119;
  assign n14199 = ~n14168;
  assign n14202 = ~n14214;
  assign n14216 = n10401 & n14229;
  assign n14212 = ~n14198;
  assign n14224 = ~n14232;
  assign n10444 = ~n10401;
  assign n14242 = ~n14251;
  assign n13938 = n14178 ^ n14179;
  assign n14127 = n14179 & n14178;
  assign n14192 = n14199 & n14200;
  assign n14148 = ~n14201;
  assign n14184 = n14202 & n14181;
  assign n14208 = n14212 & n14213;
  assign n14204 = n10444 & n12994;
  assign n14209 = n10444 & n14215;
  assign n13032 = ~n14216;
  assign n14185 = n14224 & n14225;
  assign n14218 = n14242 & n14243;
  assign n13947 = ~n13938;
  assign n14130 = ~n14127;
  assign n14104 = n14184 ^ n14185;
  assign n14170 = ~n14192;
  assign n14138 = n14204 ^ n11635;
  assign n14190 = ~n14208;
  assign n13051 = ~n14209;
  assign n14203 = ~n14185;
  assign n10364 = n14217 ^ n14218;
  assign n14219 = ~n14218;
  assign n14162 = n14104 & n14171;
  assign n14163 = ~n14104;
  assign n14182 = n14138 & n14186;
  assign n14167 = n14190 & n14191;
  assign n14183 = ~n14138;
  assign n14188 = n13051 & n13032;
  assign n14193 = n14202 & n14203;
  assign n14187 = n10364 & n12937;
  assign n14194 = n10364 & n14205;
  assign n10366 = ~n10364;
  assign n14210 = n14219 & n14220;
  assign n14133 = ~n14162;
  assign n14151 = n14163 & n118;
  assign n14146 = n14167 ^ n14168;
  assign n14140 = ~n14182;
  assign n14173 = n14183 & n14153;
  assign n14169 = ~n14167;
  assign n14114 = n14187 ^ n11659;
  assign n13049 = ~n14188;
  assign n14180 = ~n14193;
  assign n13010 = ~n14194;
  assign n14189 = n10366 & n12989;
  assign n14195 = ~n14210;
  assign n14128 = n119 ^ n14146;
  assign n14106 = ~n14151;
  assign n14161 = n14169 & n14170;
  assign n14164 = n14114 & n14172;
  assign n14155 = ~n14173;
  assign n14152 = n14180 & n14181;
  assign n14165 = ~n14114;
  assign n12992 = ~n14189;
  assign n14175 = n14195 & n14196;
  assign n12690 = n14127 ^ n14128;
  assign n14129 = ~n14128;
  assign n14137 = n14152 ^ n14153;
  assign n14147 = ~n14161;
  assign n14116 = ~n14164;
  assign n14156 = n14165 & n14095;
  assign n14154 = ~n14152;
  assign n10321 = n14174 ^ n14175;
  assign n14176 = ~n14175;
  assign n13903 = ~n12690;
  assign n14088 = n14129 & n14130;
  assign n14121 = n14137 ^ n14138;
  assign n14131 = n14147 & n14148;
  assign n14149 = n14154 & n14155;
  assign n14097 = ~n14156;
  assign n14145 = n10321 & n12904;
  assign n14157 = n10321 & n12970;
  assign n10289 = ~n10321;
  assign n14166 = n14176 & n14177;
  assign n14112 = n14121 & n117;
  assign n14103 = n118 ^ n14131;
  assign n14110 = ~n14121;
  assign n14132 = ~n14131;
  assign n14134 = n14145 ^ n11503;
  assign n14139 = ~n14149;
  assign n12972 = ~n14157;
  assign n14150 = n10289 & n14158;
  assign n14159 = ~n14166;
  assign n14089 = n14103 ^ n14104;
  assign n14107 = n14110 & n14111;
  assign n14066 = ~n14112;
  assign n14122 = n14132 & n14133;
  assign n14125 = n14134 & n14135;
  assign n14113 = n14139 & n14140;
  assign n14123 = ~n14134;
  assign n12956 = ~n14150;
  assign n14141 = n14159 & n14160;
  assign n12634 = n14088 ^ n14089;
  assign n14045 = n14089 & n14088;
  assign n14090 = ~n14107;
  assign n14094 = n14113 ^ n14114;
  assign n14105 = ~n14122;
  assign n14117 = n14123 & n14124;
  assign n14056 = ~n14125;
  assign n14115 = ~n14113;
  assign n10315 = n14141 ^ n14142;
  assign n14143 = ~n14141;
  assign n13882 = ~n12634;
  assign n14048 = ~n14045;
  assign n14092 = n14090 & n14066;
  assign n14085 = n14094 ^ n14095;
  assign n14063 = n14105 & n14106;
  assign n14108 = n14115 & n14116;
  assign n14077 = ~n14117;
  assign n14118 = n10315 & n14126;
  assign n10258 = ~n10315;
  assign n14136 = n14143 & n14144;
  assign n14073 = n14085 & n116;
  assign n14064 = ~n14092;
  assign n14071 = ~n14085;
  assign n14091 = ~n14063;
  assign n14074 = n14077 & n14056;
  assign n14096 = ~n14108;
  assign n14098 = n10258 & n12845;
  assign n12914 = ~n14118;
  assign n14109 = n10258 & n12933;
  assign n14119 = ~n14136;
  assign n14046 = n14063 ^ n14064;
  assign n14067 = n14071 & n14072;
  assign n14029 = ~n14073;
  assign n14086 = n14090 & n14091;
  assign n14075 = n14096 & n14097;
  assign n14034 = n14098 ^ n11516;
  assign n12935 = ~n14109;
  assign n14100 = n14119 & n14120;
  assign n13848 = n14045 ^ n14046;
  assign n14047 = ~n14046;
  assign n14050 = ~n14067;
  assign n14010 = n14074 ^ n14075;
  assign n14065 = ~n14086;
  assign n14078 = n14034 & n14018;
  assign n14076 = ~n14075;
  assign n14079 = ~n14034;
  assign n10291 = n14099 ^ n14100;
  assign n14101 = ~n14100;
  assign n13842 = ~n13848;
  assign n14015 = n14047 & n14048;
  assign n14031 = n14050 & n14029;
  assign n14053 = n14010 & n14061;
  assign n14032 = n14065 & n14066;
  assign n14054 = ~n14010;
  assign n14068 = n14076 & n14077;
  assign n14036 = ~n14078;
  assign n14069 = n14079 & n14080;
  assign n14062 = n10291 & n12838;
  assign n14082 = n10291 & n14087;
  assign n10298 = ~n10291;
  assign n14093 = n14101 & n14102;
  assign n14016 = n14031 ^ n14032;
  assign n14012 = ~n14053;
  assign n14051 = n14054 & n115;
  assign n14049 = ~n14032;
  assign n13977 = n14062 ^ n11342;
  assign n14055 = ~n14068;
  assign n14020 = ~n14069;
  assign n14070 = n10298 & n14081;
  assign n12890 = ~n14082;
  assign n14083 = ~n14093;
  assign n12450 = n14015 ^ n14016;
  assign n13967 = n14016 & n14015;
  assign n14041 = n14049 & n14050;
  assign n13992 = ~n14051;
  assign n14044 = n13977 & n14000;
  assign n14033 = n14055 & n14056;
  assign n14042 = ~n13977;
  assign n12872 = ~n14070;
  assign n14057 = n14083 & n14084;
  assign n13793 = ~n12450;
  assign n13975 = ~n13967;
  assign n14017 = n14033 ^ n14034;
  assign n14028 = ~n14041;
  assign n14037 = n14042 & n14043;
  assign n14002 = ~n14044;
  assign n14035 = ~n14033;
  assign n12887 = n12890 & n12872;
  assign n14038 = n14057 ^ n14058;
  assign n14059 = ~n14057;
  assign n13970 = n14017 ^ n14018;
  assign n14009 = n14028 & n14029;
  assign n14030 = n14035 & n14036;
  assign n13979 = ~n14037;
  assign n10182 = n11257 ^ n14038;
  assign n14052 = n14059 & n14060;
  assign n13997 = n13970 & n14006;
  assign n13990 = n14009 ^ n14010;
  assign n13998 = ~n13970;
  assign n14011 = ~n14009;
  assign n14008 = n10182 & n12777;
  assign n14021 = n10182 & n14027;
  assign n14019 = ~n14030;
  assign n10261 = ~n10182;
  assign n14039 = ~n14052;
  assign n13968 = n115 ^ n13990;
  assign n13972 = ~n13997;
  assign n13993 = n13998 & n114;
  assign n13934 = n14008 ^ n11257;
  assign n14007 = n14011 & n14012;
  assign n13999 = n14019 & n14020;
  assign n12850 = ~n14021;
  assign n14013 = n10261 & n14022;
  assign n14023 = n14039 & n14040;
  assign n12371 = n13967 ^ n13968;
  assign n13646 = n13968 & n13975;
  assign n13950 = ~n13993;
  assign n13987 = n13934 & n13994;
  assign n13976 = n13999 ^ n14000;
  assign n13988 = ~n13934;
  assign n13991 = ~n14007;
  assign n14001 = ~n13999;
  assign n12823 = ~n14013;
  assign n14003 = n14023 ^ n14024;
  assign n14025 = ~n14023;
  assign n12406 = ~n12371;
  assign n13912 = n13976 ^ n13977;
  assign n13936 = ~n13987;
  assign n13980 = n13988 & n13958;
  assign n13969 = n13991 & n13992;
  assign n13995 = n14001 & n14002;
  assign n13996 = n12850 & n12823;
  assign n10123 = n11303 ^ n14003;
  assign n14014 = n14025 & n14026;
  assign n13955 = n13912 & n13964;
  assign n13948 = n13969 ^ n13970;
  assign n13956 = ~n13912;
  assign n13960 = ~n13980;
  assign n13971 = ~n13969;
  assign n13981 = n10123 & n13989;
  assign n13966 = n10123 & n12739;
  assign n13978 = ~n13995;
  assign n12848 = ~n13996;
  assign n10224 = ~n10123;
  assign n14004 = ~n14014;
  assign n13616 = n114 ^ n13948;
  assign n13930 = ~n13955;
  assign n13951 = n13956 & n113;
  assign n13952 = n13966 ^ n11285;
  assign n13965 = n13971 & n13972;
  assign n13957 = n13978 & n13979;
  assign n12799 = ~n13981;
  assign n13973 = n10224 & n13982;
  assign n13983 = n14004 & n14005;
  assign n13889 = n13616 & n13646;
  assign n13914 = ~n13951;
  assign n13944 = n13952 & n13953;
  assign n13933 = n13957 ^ n13958;
  assign n13945 = ~n13952;
  assign n13949 = ~n13965;
  assign n13959 = ~n13957;
  assign n12775 = ~n13973;
  assign n13961 = n13983 ^ n13984;
  assign n13985 = ~n13983;
  assign n13926 = n13933 ^ n13934;
  assign n13899 = ~n13944;
  assign n13937 = n13945 & n13946;
  assign n13928 = n13949 & n13950;
  assign n13954 = n13959 & n13960;
  assign n12796 = n12799 & n12775;
  assign n10177 = n13961 ^ n11209;
  assign n13974 = n13985 & n13986;
  assign n13919 = n13926 & n112;
  assign n13911 = n113 ^ n13928;
  assign n13917 = ~n13926;
  assign n13921 = ~n13937;
  assign n13929 = ~n13928;
  assign n13939 = n10177 & n13947;
  assign n13935 = ~n13954;
  assign n10080 = ~n10177;
  assign n13962 = ~n13974;
  assign n13890 = n13911 ^ n13912;
  assign n13915 = n13917 & n13918;
  assign n13873 = ~n13919;
  assign n13908 = n13921 & n13899;
  assign n13927 = n13929 & n13930;
  assign n13909 = n13935 & n13936;
  assign n13931 = n10080 & n13938;
  assign n13922 = n10080 & n12543;
  assign n12721 = ~n13939;
  assign n13940 = n13962 & n13963;
  assign n11746 = n13889 ^ n13890;
  assign n13849 = n13890 & n13889;
  assign n13852 = n13908 ^ n13909;
  assign n13892 = ~n13915;
  assign n13878 = n13922 ^ n11209;
  assign n13913 = ~n13927;
  assign n13920 = ~n13909;
  assign n12748 = ~n13931;
  assign n13923 = n13940 ^ n13941;
  assign n13942 = ~n13940;
  assign n12814 = n11746 ^ n13869;
  assign n13758 = n11746 & n11790;
  assign n11744 = ~n11746;
  assign n13887 = n13852 & n13893;
  assign n13894 = n13892 & n13873;
  assign n13888 = ~n13852;
  assign n13901 = n13878 & n13910;
  assign n13870 = n13913 & n13914;
  assign n13900 = ~n13878;
  assign n13916 = n13920 & n13921;
  assign n12745 = n12748 & n12721;
  assign n10127 = n13923 ^ n11126;
  assign n13932 = n13942 & n13943;
  assign n13829 = n12814 ^ n12791;
  assign n13854 = ~n13887;
  assign n13876 = n13888 & n127;
  assign n13871 = ~n13894;
  assign n13895 = n13900 & n13858;
  assign n13880 = ~n13901;
  assign n13891 = ~n13870;
  assign n13902 = n10127 & n12690;
  assign n13898 = ~n13916;
  assign n10114 = ~n10127;
  assign n13924 = ~n13932;
  assign n13807 = n13829 & n12791;
  assign n9893 = ~n13829;
  assign n13850 = n13870 ^ n13871;
  assign n13824 = ~n13876;
  assign n13886 = n13891 & n13892;
  assign n13860 = ~n13895;
  assign n13877 = n13898 & n13899;
  assign n12667 = ~n13902;
  assign n13881 = n10114 & n12582;
  assign n13896 = n10114 & n13903;
  assign n13904 = n13924 & n13925;
  assign n13773 = n13807 ^ n13808;
  assign n13784 = n13807 ^ n13809;
  assign n13830 = n13849 ^ n13850;
  assign n13794 = n13850 & n13849;
  assign n13857 = n13877 ^ n13878;
  assign n13811 = n13881 ^ n11002;
  assign n13872 = ~n13886;
  assign n13879 = ~n13877;
  assign n12692 = ~n13896;
  assign n10093 = n13904 ^ n13905;
  assign n13906 = ~n13904;
  assign n11921 = n327 ^ n13773;
  assign n13628 = n13784 & n13785;
  assign n13545 = n13773 & n327;
  assign n13820 = n13830 & n11759;
  assign n13821 = ~n13830;
  assign n13797 = ~n13794;
  assign n13765 = n13857 ^ n13858;
  assign n13862 = n13811 & n13868;
  assign n13851 = n13872 & n13873;
  assign n13861 = ~n13811;
  assign n13874 = n13879 & n13880;
  assign n13883 = n10093 & n12634;
  assign n10017 = ~n10093;
  assign n13897 = n13906 & n13907;
  assign n13136 = ~n11921;
  assign n13763 = ~n13820;
  assign n13818 = n13821 & n11761;
  assign n13833 = n13765 & n126;
  assign n13822 = n13851 ^ n13852;
  assign n13831 = ~n13765;
  assign n13855 = n13861 & n13835;
  assign n13813 = ~n13862;
  assign n13853 = ~n13851;
  assign n13859 = ~n13874;
  assign n13863 = n10017 & n12392;
  assign n13875 = n10017 & n13882;
  assign n12601 = ~n13883;
  assign n13884 = ~n13897;
  assign n13798 = ~n13818;
  assign n13795 = n127 ^ n13822;
  assign n13825 = n13831 & n13832;
  assign n13767 = ~n13833;
  assign n13845 = n13853 & n13854;
  assign n13837 = ~n13855;
  assign n13834 = n13859 & n13860;
  assign n13846 = n13863 ^ n11041;
  assign n12636 = ~n13875;
  assign n13865 = n13884 & n13885;
  assign n13774 = n13794 ^ n13795;
  assign n13786 = n13798 & n13758;
  assign n13787 = n13798 & n13763;
  assign n13796 = ~n13795;
  assign n13801 = ~n13825;
  assign n13810 = n13834 ^ n13835;
  assign n13823 = ~n13845;
  assign n13840 = n13846 & n13847;
  assign n13836 = ~n13834;
  assign n13838 = ~n13846;
  assign n9979 = n13864 ^ n13865;
  assign n13866 = ~n13865;
  assign n13761 = n13774 & n11611;
  assign n13703 = ~n13774;
  assign n13762 = ~n13786;
  assign n13759 = ~n13787;
  assign n13740 = n13796 & n13797;
  assign n13788 = n13810 ^ n13811;
  assign n13799 = n13823 & n13824;
  assign n13826 = n13836 & n13837;
  assign n13827 = n13838 & n13839;
  assign n13750 = ~n13840;
  assign n13841 = n9979 & n13848;
  assign n13819 = n9979 & n12459;
  assign n10033 = ~n9979;
  assign n13856 = n13866 & n13867;
  assign n9828 = n13758 ^ n13759;
  assign n13757 = n13703 & n11617;
  assign n13739 = ~n13761;
  assign n13760 = n13762 & n13763;
  assign n13777 = n13788 & n125;
  assign n13764 = n126 ^ n13799;
  assign n13775 = ~n13788;
  assign n13800 = ~n13799;
  assign n13802 = n13819 ^ n10934;
  assign n13812 = ~n13826;
  assign n13779 = ~n13827;
  assign n12563 = ~n13841;
  assign n13828 = n10033 & n13842;
  assign n13843 = ~n13856;
  assign n13710 = n9828 & n12711;
  assign n9836 = ~n9828;
  assign n13712 = ~n13757;
  assign n13734 = ~n13760;
  assign n13741 = n13764 ^ n13765;
  assign n13768 = n13775 & n13776;
  assign n13716 = ~n13777;
  assign n13789 = n13800 & n13801;
  assign n13790 = n13802 & n13803;
  assign n13769 = n13812 & n13813;
  assign n13804 = n13779 & n13750;
  assign n13791 = ~n13802;
  assign n12525 = ~n13828;
  assign n13814 = n13843 & n13844;
  assign n13691 = n13710 ^ n11761;
  assign n13704 = n13734 ^ n11617;
  assign n13733 = n13739 & n13734;
  assign n13720 = n13740 ^ n13741;
  assign n13693 = n13741 & n13740;
  assign n13743 = ~n13768;
  assign n13766 = ~n13789;
  assign n13699 = ~n13790;
  assign n13780 = n13791 & n13792;
  assign n13778 = ~n13769;
  assign n13770 = ~n13804;
  assign n13805 = n12563 & n12525;
  assign n9923 = n13814 ^ n13815;
  assign n13816 = ~n13814;
  assign n13678 = n13691 & n13692;
  assign n9786 = n13703 ^ n13704;
  assign n13679 = ~n13691;
  assign n13713 = n13720 & n11545;
  assign n13711 = ~n13733;
  assign n13714 = ~n13720;
  assign n13721 = n13743 & n13716;
  assign n13722 = n13766 & n13767;
  assign n13748 = n13769 ^ n13770;
  assign n13771 = n13778 & n13779;
  assign n13726 = ~n13780;
  assign n13781 = n9923 & n13793;
  assign n12561 = ~n13805;
  assign n10006 = ~n9923;
  assign n13806 = n13816 & n13817;
  assign n13630 = ~n13678;
  assign n13670 = n13679 & n13680;
  assign n9811 = ~n9786;
  assign n13649 = n13711 & n13712;
  assign n13682 = ~n13713;
  assign n13705 = n13714 & n11471;
  assign n13694 = n13721 ^ n13722;
  assign n13746 = n13748 & n124;
  assign n13742 = ~n13722;
  assign n13744 = ~n13748;
  assign n13751 = n13726 & n13699;
  assign n13749 = ~n13771;
  assign n12452 = ~n13781;
  assign n13772 = n10006 & n12450;
  assign n13752 = n10006 & n12240;
  assign n13782 = ~n13806;
  assign n13647 = n9811 & n12613;
  assign n13652 = ~n13670;
  assign n13673 = n13693 ^ n13694;
  assign n13681 = ~n13649;
  assign n13654 = ~n13705;
  assign n13656 = n13694 & n13693;
  assign n13735 = n13742 & n13743;
  assign n13736 = n13744 & n13745;
  assign n13659 = ~n13746;
  assign n13723 = n13749 & n13750;
  assign n13724 = ~n13751;
  assign n13642 = n13752 ^ n10863;
  assign n12485 = ~n13772;
  assign n13754 = n13782 & n13783;
  assign n13625 = n13647 ^ n11611;
  assign n13648 = n13652 & n13628;
  assign n13627 = n13652 & n13630;
  assign n13661 = n13673 & n11441;
  assign n13671 = n13681 & n13682;
  assign n13672 = n13682 & n13654;
  assign n13662 = ~n13673;
  assign n13706 = n13723 ^ n13724;
  assign n13715 = ~n13735;
  assign n13686 = ~n13736;
  assign n13727 = n13642 & n13664;
  assign n13725 = ~n13723;
  assign n13728 = ~n13642;
  assign n9946 = n13753 ^ n13754;
  assign n13756 = n13754 & n13731;
  assign n13755 = ~n13754;
  assign n13617 = n13625 & n13626;
  assign n13607 = n13627 ^ n13628;
  assign n13618 = ~n13625;
  assign n13629 = ~n13648;
  assign n13632 = ~n13661;
  assign n13655 = n13662 & n11463;
  assign n13653 = ~n13671;
  assign n13650 = ~n13672;
  assign n13697 = n13706 & n123;
  assign n13684 = n13715 & n13716;
  assign n13683 = n13686 & n13659;
  assign n13695 = ~n13706;
  assign n13717 = n13725 & n13726;
  assign n13666 = ~n13727;
  assign n13718 = n13728 & n13729;
  assign n13707 = n9946 & n12272;
  assign n9951 = ~n9946;
  assign n13747 = n13755 & n13738;
  assign n13737 = ~n13756;
  assign n13594 = n13607 & n326;
  assign n13561 = ~n13617;
  assign n13608 = n13618 & n13619;
  assign n13592 = ~n13607;
  assign n13559 = n13629 & n13630;
  assign n9742 = n13649 ^ n13650;
  assign n13597 = n13653 & n13654;
  assign n13596 = ~n13655;
  assign n13657 = n13683 ^ n13684;
  assign n13687 = n13695 & n13696;
  assign n13604 = ~n13697;
  assign n13685 = ~n13684;
  assign n13688 = n13707 ^ n10742;
  assign n13698 = ~n13717;
  assign n13644 = ~n13718;
  assign n13732 = n13737 & n13738;
  assign n13730 = ~n13747;
  assign n13589 = n13592 & n13593;
  assign n13547 = ~n13594;
  assign n13587 = ~n13608;
  assign n13588 = ~n13559;
  assign n9775 = ~n9742;
  assign n13633 = n13632 & n13596;
  assign n13631 = ~n13597;
  assign n13640 = n13656 ^ n13657;
  assign n13599 = n13657 & n13656;
  assign n13674 = n13685 & n13686;
  assign n13639 = ~n13687;
  assign n13675 = n13688 & n13689;
  assign n13663 = n13698 & n13699;
  assign n13676 = ~n13688;
  assign n13719 = n13730 & n13731;
  assign n13708 = ~n13732;
  assign n13580 = n13587 & n13588;
  assign n13570 = ~n13589;
  assign n13558 = n13587 & n13561;
  assign n13590 = n9775 & n12568;
  assign n13620 = n13631 & n13632;
  assign n13598 = ~n13633;
  assign n13635 = n13640 & n11392;
  assign n13634 = ~n13640;
  assign n13602 = ~n13599;
  assign n13636 = n13639 & n13604;
  assign n13641 = n13663 ^ n13664;
  assign n13658 = ~n13674;
  assign n13586 = ~n13675;
  assign n13667 = n13676 & n13677;
  assign n13665 = ~n13663;
  assign n13702 = n13708 & n13709;
  assign n13700 = ~n13719;
  assign n13492 = n13558 ^ n13559;
  assign n13562 = n13570 & n13545;
  assign n13544 = n13570 & n13547;
  assign n13560 = ~n13580;
  assign n13505 = n13590 ^ n11545;
  assign n9732 = n13597 ^ n13598;
  assign n13595 = ~n13620;
  assign n13621 = n13634 & n11403;
  assign n13573 = ~n13635;
  assign n13552 = n13641 ^ n13642;
  assign n13637 = n13658 & n13659;
  assign n13660 = n13665 & n13666;
  assign n13614 = ~n13667;
  assign n13690 = n13700 & n13701;
  assign n13669 = ~n13702;
  assign n13537 = n13492 & n13543;
  assign n13514 = n13544 ^ n13545;
  assign n13538 = ~n13492;
  assign n13539 = n13560 & n13561;
  assign n13546 = ~n13562;
  assign n13563 = n13505 & n13571;
  assign n13564 = ~n13505;
  assign n9707 = ~n9732;
  assign n13565 = n13595 & n13596;
  assign n13550 = ~n13621;
  assign n13609 = n13552 & n13622;
  assign n13600 = n13636 ^ n13637;
  assign n13610 = ~n13552;
  assign n13638 = ~n13637;
  assign n13645 = n13614 & n13586;
  assign n13643 = ~n13660;
  assign n13668 = ~n13690;
  assign n13112 = n13514 ^ n11921;
  assign n13116 = n13514 ^ n13136;
  assign n13464 = n13514 & n11921;
  assign n13515 = ~n13537;
  assign n13531 = n13538 & n325;
  assign n13506 = n13539 ^ n13540;
  assign n13517 = n13546 & n13547;
  assign n13542 = ~n13539;
  assign n13509 = ~n13563;
  assign n13555 = n13564 & n13540;
  assign n13548 = n9707 & n12381;
  assign n13572 = ~n13565;
  assign n13591 = n13550 & n13573;
  assign n13581 = n13599 ^ n13600;
  assign n13578 = ~n13609;
  assign n13605 = n13610 & n122;
  assign n13601 = ~n13600;
  assign n13623 = n13638 & n13639;
  assign n13611 = n13643 & n13644;
  assign n13612 = ~n13645;
  assign n9873 = n13668 & n13669;
  assign n13490 = n13505 ^ n13506;
  assign n13467 = ~n13464;
  assign n13491 = n325 ^ n13517;
  assign n13494 = ~n13531;
  assign n13516 = ~n13517;
  assign n13533 = n13548 ^ n11441;
  assign n13541 = ~n13555;
  assign n13567 = n13572 & n13573;
  assign n13574 = n13581 & n11310;
  assign n13566 = ~n13591;
  assign n13575 = ~n13581;
  assign n13525 = n13601 & n13602;
  assign n13554 = ~n13605;
  assign n13528 = n13611 ^ n13612;
  assign n13603 = ~n13623;
  assign n13613 = ~n13611;
  assign n13615 = n13646 ^ n9873;
  assign n13624 = n9873 & n13651;
  assign n10694 = ~n9873;
  assign n13482 = n13490 & n324;
  assign n13465 = n13491 ^ n13492;
  assign n13480 = ~n13490;
  assign n13507 = n13515 & n13516;
  assign n13520 = n13533 & n13534;
  assign n13532 = n13541 & n13542;
  assign n13518 = ~n13533;
  assign n9729 = n13565 ^ n13566;
  assign n13549 = ~n13567;
  assign n13498 = ~n13574;
  assign n13568 = n13575 & n11296;
  assign n13584 = n13528 & n121;
  assign n13576 = n13603 & n13604;
  assign n13582 = ~n13528;
  assign n13606 = n13613 & n13614;
  assign n12305 = n13615 ^ n13616;
  assign n13535 = n13624 ^ n10610;
  assign n11849 = n13464 ^ n13465;
  assign n13476 = n13480 & n13481;
  assign n13435 = ~n13482;
  assign n13466 = ~n13465;
  assign n13493 = ~n13507;
  assign n13511 = n13518 & n13519;
  assign n13460 = ~n13520;
  assign n13508 = ~n13532;
  assign n13522 = n13549 & n13550;
  assign n9719 = ~n9729;
  assign n13524 = ~n13568;
  assign n13551 = n122 ^ n13576;
  assign n13579 = n13582 & n13583;
  assign n13503 = ~n13584;
  assign n13577 = ~n13576;
  assign n13585 = ~n13606;
  assign n12290 = ~n12305;
  assign n13046 = ~n11849;
  assign n13413 = n13466 & n13467;
  assign n13456 = ~n13476;
  assign n13433 = n13493 & n13494;
  assign n13461 = n13508 & n13509;
  assign n13484 = ~n13511;
  assign n13510 = n9719 & n12265;
  assign n13523 = ~n13522;
  assign n13521 = n13524 & n13498;
  assign n13526 = n13551 ^ n13552;
  assign n13569 = n13577 & n13578;
  assign n13530 = ~n13579;
  assign n13556 = n13585 & n13586;
  assign n13432 = n13456 & n13435;
  assign n13457 = ~n13433;
  assign n13488 = n13484 & n13460;
  assign n13483 = ~n13461;
  assign n13495 = n13510 ^ n11392;
  assign n9689 = n13521 ^ n13522;
  assign n13512 = n13523 & n13524;
  assign n13445 = n13525 ^ n13526;
  assign n13471 = n13526 & n13525;
  assign n13536 = n13556 ^ n13557;
  assign n13553 = ~n13569;
  assign n13414 = n13432 ^ n13433;
  assign n13452 = n13456 & n13457;
  assign n13478 = n13483 & n13484;
  assign n13462 = ~n13488;
  assign n13487 = n13495 & n13496;
  assign n13477 = n9689 & n12308;
  assign n13485 = ~n13495;
  assign n13499 = n13445 & n11218;
  assign n9639 = ~n9689;
  assign n13497 = ~n13512;
  assign n13500 = ~n13445;
  assign n13504 = n13535 ^ n13536;
  assign n13527 = n13553 & n13554;
  assign n13030 = n13413 ^ n13414;
  assign n13376 = n13414 & n13413;
  assign n13434 = ~n13452;
  assign n13443 = n13461 ^ n13462;
  assign n13381 = n13477 ^ n11296;
  assign n13459 = ~n13478;
  assign n13479 = n13485 & n13486;
  assign n13419 = ~n13487;
  assign n13468 = n13497 & n13498;
  assign n13447 = ~n13499;
  assign n13489 = n13500 & n11108;
  assign n13475 = n120 ^ n13504;
  assign n13501 = n13527 ^ n13528;
  assign n13529 = ~n13527;
  assign n13034 = ~n13030;
  assign n13399 = n13434 & n13435;
  assign n13440 = n13443 & n323;
  assign n13438 = ~n13443;
  assign n13454 = n13381 & n13458;
  assign n13428 = n13459 & n13460;
  assign n13453 = ~n13381;
  assign n13444 = n13468 ^ n11218;
  assign n13437 = ~n13479;
  assign n13469 = ~n13468;
  assign n13470 = ~n13489;
  assign n13472 = n121 ^ n13501;
  assign n13513 = n13529 & n13530;
  assign n13416 = ~n13399;
  assign n13431 = n13438 & n13439;
  assign n13395 = ~n13440;
  assign n9633 = n13444 ^ n13445;
  assign n13442 = n13453 & n13401;
  assign n13383 = ~n13454;
  assign n13436 = ~n13428;
  assign n13455 = n13437 & n13419;
  assign n13463 = n13469 & n13470;
  assign n13423 = n13471 ^ n13472;
  assign n13473 = ~n13472;
  assign n13502 = ~n13513;
  assign n13409 = n9633 & n12248;
  assign n13415 = ~n13431;
  assign n13430 = n13436 & n13437;
  assign n9644 = ~n9633;
  assign n13403 = ~n13442;
  assign n13429 = ~n13455;
  assign n13449 = n13423 & n11115;
  assign n13446 = ~n13463;
  assign n13448 = ~n13423;
  assign n13450 = n13473 & n13471;
  assign n13474 = n13502 & n13503;
  assign n13396 = n13409 ^ n11108;
  assign n13408 = n13415 & n13416;
  assign n13398 = n13415 & n13395;
  assign n13417 = n13428 ^ n13429;
  assign n13418 = ~n13430;
  assign n13422 = n13446 & n13447;
  assign n13441 = n13448 & n11132;
  assign n13425 = ~n13449;
  assign n13451 = n13474 ^ n13475;
  assign n13392 = n13396 & n13397;
  assign n13377 = n13398 ^ n13399;
  assign n13390 = ~n13396;
  assign n13394 = ~n13408;
  assign n13412 = n13417 & n322;
  assign n13400 = n13418 & n13419;
  assign n13410 = ~n13417;
  assign n13405 = n13422 ^ n13423;
  assign n13424 = ~n13422;
  assign n13407 = ~n13441;
  assign n13387 = n13450 ^ n13451;
  assign n12968 = n13376 ^ n13377;
  assign n13354 = n13377 & n13376;
  assign n13385 = n13390 & n13391;
  assign n13344 = ~n13392;
  assign n13374 = n13394 & n13395;
  assign n13380 = n13400 ^ n13401;
  assign n9565 = n11132 ^ n13405;
  assign n13404 = n13410 & n13411;
  assign n13363 = ~n13412;
  assign n13402 = ~n13400;
  assign n13420 = n13424 & n13425;
  assign n13427 = n13387 & n11063;
  assign n13426 = ~n13387;
  assign n12974 = ~n12968;
  assign n13330 = n13380 ^ n13381;
  assign n13367 = ~n13385;
  assign n13379 = ~n13374;
  assign n13393 = n13402 & n13403;
  assign n9626 = ~n9565;
  assign n13378 = ~n13404;
  assign n13406 = ~n13420;
  assign n13421 = n13426 & n11045;
  assign n13372 = ~n13427;
  assign n13366 = n13330 & n321;
  assign n13356 = n13367 & n13344;
  assign n13364 = ~n13330;
  assign n13375 = n13378 & n13379;
  assign n13369 = n9626 & n12171;
  assign n13373 = n13378 & n13363;
  assign n13382 = ~n13393;
  assign n13386 = n13406 & n13407;
  assign n13389 = ~n13421;
  assign n13358 = n13364 & n13365;
  assign n13332 = ~n13366;
  assign n13359 = n13369 ^ n11115;
  assign n13355 = n13373 ^ n13374;
  assign n13362 = ~n13375;
  assign n13357 = n13382 & n13383;
  assign n13370 = n13386 ^ n13387;
  assign n13388 = ~n13386;
  assign n11677 = n13354 ^ n13355;
  assign n13290 = n13356 ^ n13357;
  assign n13341 = ~n13358;
  assign n13347 = n13359 & n13360;
  assign n13308 = n13355 & n13354;
  assign n13340 = n13362 & n13363;
  assign n13348 = ~n13359;
  assign n9523 = n11045 ^ n13370;
  assign n13368 = ~n13357;
  assign n13384 = n13388 & n13389;
  assign n13329 = n321 ^ n13340;
  assign n12930 = ~n11677;
  assign n13301 = ~n13290;
  assign n13316 = ~n13347;
  assign n13345 = n13348 & n13349;
  assign n13342 = ~n13340;
  assign n13361 = n13367 & n13368;
  assign n9590 = ~n9523;
  assign n13371 = ~n13384;
  assign n13309 = n13329 ^ n13330;
  assign n13339 = n13341 & n13342;
  assign n13333 = ~n13345;
  assign n13336 = n9590 & n12060;
  assign n13343 = ~n13361;
  assign n13350 = n13371 & n13372;
  assign n12885 = n13308 ^ n13309;
  assign n13270 = n13309 & n13308;
  assign n13335 = n13333 & n13316;
  assign n13273 = n13336 ^ n11045;
  assign n13331 = ~n13339;
  assign n13313 = n13343 & n13344;
  assign n9534 = n13350 ^ n13351;
  assign n13352 = ~n13350;
  assign n12896 = ~n12885;
  assign n13279 = ~n13270;
  assign n13320 = n13273 & n13327;
  assign n13310 = n13331 & n13332;
  assign n13314 = ~n13335;
  assign n13321 = ~n13273;
  assign n13334 = ~n13313;
  assign n9528 = ~n9534;
  assign n13346 = n13352 & n13353;
  assign n13289 = n320 ^ n13310;
  assign n13242 = n13313 ^ n13314;
  assign n13312 = n13310 & n13319;
  assign n13275 = ~n13320;
  assign n13317 = n13321 & n13296;
  assign n13311 = ~n13310;
  assign n13328 = n13333 & n13334;
  assign n13322 = n9528 & n12051;
  assign n13337 = ~n13346;
  assign n13271 = n13289 ^ n13290;
  assign n13294 = n13242 & n335;
  assign n13292 = ~n13242;
  assign n13307 = n13311 & n320;
  assign n13300 = ~n13312;
  assign n13297 = ~n13317;
  assign n13257 = n13322 ^ n10973;
  assign n13315 = ~n13328;
  assign n13323 = n13337 & n13338;
  assign n11517 = n13270 ^ n13271;
  assign n13219 = n13271 & n13279;
  assign n13286 = n13292 & n13293;
  assign n13244 = ~n13294;
  assign n13291 = n13300 & n13301;
  assign n13281 = ~n13307;
  assign n13304 = n13257 & n13235;
  assign n13295 = n13315 & n13316;
  assign n13302 = ~n13257;
  assign n9463 = n13323 ^ n13324;
  assign n13325 = ~n13323;
  assign n12870 = ~n11517;
  assign n13263 = ~n13286;
  assign n13280 = ~n13291;
  assign n13272 = n13295 ^ n13296;
  assign n13299 = n13302 & n13303;
  assign n13259 = ~n13304;
  assign n13298 = ~n13295;
  assign n13288 = n9463 & n12011;
  assign n9520 = ~n9463;
  assign n13318 = n13325 & n13326;
  assign n13260 = n13272 ^ n13273;
  assign n13261 = n13280 & n13281;
  assign n13276 = n13288 ^ n10867;
  assign n13287 = n13297 & n13298;
  assign n13237 = ~n13299;
  assign n13305 = ~n13318;
  assign n13254 = n13260 & n334;
  assign n13241 = n335 ^ n13261;
  assign n13252 = ~n13260;
  assign n13262 = ~n13261;
  assign n13269 = n13276 & n13277;
  assign n13267 = ~n13276;
  assign n13274 = ~n13287;
  assign n13283 = n13305 & n13306;
  assign n13220 = n13241 ^ n13242;
  assign n13249 = n13252 & n13253;
  assign n13202 = ~n13254;
  assign n13255 = n13262 & n13263;
  assign n13264 = n13267 & n13268;
  assign n13199 = ~n13269;
  assign n13256 = n13274 & n13275;
  assign n9472 = n13282 ^ n13283;
  assign n13284 = ~n13283;
  assign n11478 = n13219 ^ n13220;
  assign n13221 = ~n13220;
  assign n13224 = ~n13249;
  assign n13243 = ~n13255;
  assign n13234 = n13256 ^ n13257;
  assign n13218 = ~n13264;
  assign n13258 = ~n13256;
  assign n13251 = n9472 & n11978;
  assign n9481 = ~n9472;
  assign n13278 = n13284 & n13285;
  assign n12832 = ~n11478;
  assign n13185 = n13221 & n13219;
  assign n13230 = n13224 & n13202;
  assign n13168 = n13234 ^ n13235;
  assign n13208 = n13243 & n13244;
  assign n13245 = n13218 & n13199;
  assign n13238 = n13251 ^ n10726;
  assign n13250 = n13258 & n13259;
  assign n13265 = ~n13278;
  assign n13212 = n13168 & n13222;
  assign n13209 = ~n13230;
  assign n13213 = ~n13168;
  assign n13223 = ~n13208;
  assign n13231 = n13238 & n13239;
  assign n13216 = ~n13245;
  assign n13232 = ~n13238;
  assign n13236 = ~n13250;
  assign n13246 = n13265 & n13266;
  assign n13193 = n13208 ^ n13209;
  assign n13189 = ~n13212;
  assign n13210 = n13213 & n333;
  assign n13214 = n13223 & n13224;
  assign n13164 = ~n13231;
  assign n13225 = n13232 & n13233;
  assign n13215 = n13236 & n13237;
  assign n13227 = n13246 ^ n10697;
  assign n13247 = ~n13246;
  assign n12772 = n13185 ^ n13193;
  assign n13143 = n13193 & n13185;
  assign n13186 = ~n13193;
  assign n13170 = ~n13210;
  assign n13201 = ~n13214;
  assign n13203 = n13215 ^ n13216;
  assign n13184 = ~n13225;
  assign n9417 = n13226 ^ n13227;
  assign n13217 = ~n13215;
  assign n13240 = n13247 & n13248;
  assign n12778 = n13185 ^ n13186;
  assign n13146 = ~n13143;
  assign n13187 = n13201 & n13202;
  assign n13197 = n13203 & n332;
  assign n13195 = ~n13203;
  assign n13181 = n13184 & n13164;
  assign n13211 = n13217 & n13218;
  assign n9409 = ~n9417;
  assign n13228 = ~n13240;
  assign n13167 = n333 ^ n13187;
  assign n13188 = ~n13187;
  assign n13194 = n13195 & n13196;
  assign n13129 = ~n13197;
  assign n13190 = n9409 & n11936;
  assign n13198 = ~n13211;
  assign n13204 = n13228 & n13229;
  assign n13144 = n13167 ^ n13168;
  assign n13180 = n13188 & n13189;
  assign n13118 = n13190 ^ n10697;
  assign n13150 = ~n13194;
  assign n13182 = n13198 & n13199;
  assign n9323 = n13204 ^ n13205;
  assign n13206 = ~n13204;
  assign n12727 = n13143 ^ n13144;
  assign n13145 = ~n13144;
  assign n13173 = n13118 & n13178;
  assign n13169 = ~n13180;
  assign n13147 = n13150 & n13129;
  assign n13108 = n13181 ^ n13182;
  assign n13172 = ~n13118;
  assign n13183 = ~n13182;
  assign n9396 = ~n9323;
  assign n13200 = n13206 & n13207;
  assign n12719 = ~n12727;
  assign n13124 = n13145 & n13146;
  assign n13148 = n13169 & n13170;
  assign n13161 = n13108 & n13171;
  assign n13165 = n13172 & n13139;
  assign n13120 = ~n13173;
  assign n13162 = ~n13108;
  assign n13179 = n13183 & n13184;
  assign n13174 = n9396 & n11891;
  assign n13191 = ~n13200;
  assign n13127 = ~n13124;
  assign n13125 = n13147 ^ n13148;
  assign n13149 = ~n13148;
  assign n13110 = ~n13161;
  assign n13158 = n13162 & n331;
  assign n13141 = ~n13165;
  assign n13159 = n13174 ^ n10619;
  assign n13163 = ~n13179;
  assign n13175 = n13191 & n13192;
  assign n12631 = n13124 ^ n13125;
  assign n13126 = ~n13125;
  assign n13137 = n13149 & n13150;
  assign n13085 = ~n13158;
  assign n13153 = n13159 & n13160;
  assign n13138 = n13163 & n13164;
  assign n13151 = ~n13159;
  assign n13155 = n13175 ^ n10546;
  assign n13176 = ~n13175;
  assign n12641 = ~n12631;
  assign n13059 = n13126 & n13127;
  assign n13128 = ~n13137;
  assign n13117 = n13138 ^ n13139;
  assign n13142 = n13151 & n13152;
  assign n13078 = ~n13153;
  assign n9283 = n13154 ^ n13155;
  assign n13140 = ~n13138;
  assign n13166 = n13176 & n13177;
  assign n13062 = ~n13059;
  assign n13106 = n13117 ^ n13118;
  assign n13107 = n13128 & n13129;
  assign n13130 = n9283 & n13136;
  assign n13135 = n13140 & n13141;
  assign n13104 = ~n13142;
  assign n9361 = ~n9283;
  assign n13156 = ~n13166;
  assign n13099 = n13106 & n330;
  assign n13083 = n13107 ^ n13108;
  assign n13097 = ~n13106;
  assign n13109 = ~n13107;
  assign n13121 = n13104 & n13078;
  assign n13111 = n9361 & n11785;
  assign n11906 = ~n13130;
  assign n13122 = n9361 & n11921;
  assign n13119 = ~n13135;
  assign n13132 = n13156 & n13157;
  assign n13060 = n331 ^ n13083;
  assign n13092 = n13097 & n13098;
  assign n13044 = ~n13099;
  assign n13100 = n13109 & n13110;
  assign n13093 = n13111 ^ n10546;
  assign n13101 = n13119 & n13120;
  assign n13102 = ~n13121;
  assign n11923 = ~n13122;
  assign n9288 = n13131 ^ n13132;
  assign n13133 = ~n13132;
  assign n12576 = n13059 ^ n13060;
  assign n13061 = ~n13060;
  assign n13064 = ~n13092;
  assign n13088 = n13093 & n13094;
  assign n13084 = ~n13100;
  assign n13002 = n13101 ^ n13102;
  assign n13086 = ~n13093;
  assign n13103 = ~n13101;
  assign n13096 = n9288 & n11843;
  assign n13113 = n9288 & n13116;
  assign n9295 = ~n9288;
  assign n13123 = n13133 & n13134;
  assign n12559 = ~n12576;
  assign n13035 = n13061 & n13062;
  assign n13053 = n13064 & n13044;
  assign n13054 = n13084 & n13085;
  assign n13076 = n13002 & n329;
  assign n13081 = n13086 & n13087;
  assign n13040 = ~n13088;
  assign n13074 = ~n13002;
  assign n13079 = n13096 ^ n10531;
  assign n13095 = n13103 & n13104;
  assign n13105 = n9295 & n13112;
  assign n11886 = ~n13113;
  assign n13114 = ~n13123;
  assign n13036 = n13053 ^ n13054;
  assign n13063 = ~n13054;
  assign n13070 = n13074 & n13075;
  assign n13004 = ~n13076;
  assign n13071 = n13079 & n13080;
  assign n13057 = ~n13081;
  assign n13072 = ~n13079;
  assign n13077 = ~n13095;
  assign n11871 = ~n13105;
  assign n13089 = n13114 & n13115;
  assign n12523 = n13035 ^ n13036;
  assign n12983 = n13036 & n13035;
  assign n13055 = n13063 & n13064;
  assign n13058 = n13057 & n13040;
  assign n13027 = ~n13070;
  assign n12999 = ~n13071;
  assign n13065 = n13072 & n13073;
  assign n13037 = n13077 & n13078;
  assign n11883 = n11886 & n11871;
  assign n13067 = n13089 ^ n10461;
  assign n13090 = ~n13089;
  assign n12532 = ~n12523;
  assign n13043 = ~n13055;
  assign n13038 = ~n13058;
  assign n13023 = ~n13065;
  assign n9224 = n13066 ^ n13067;
  assign n13056 = ~n13037;
  assign n13082 = n13090 & n13091;
  assign n13028 = n13037 ^ n13038;
  assign n13025 = n13043 & n13044;
  assign n13045 = n13023 & n12999;
  assign n13033 = n9224 & n11739;
  assign n13047 = n9224 & n11849;
  assign n13052 = n13056 & n13057;
  assign n9246 = ~n9224;
  assign n13068 = ~n13082;
  assign n13001 = n329 ^ n13025;
  assign n13019 = n13028 & n328;
  assign n12960 = n13033 ^ n10461;
  assign n13016 = ~n13028;
  assign n13026 = ~n13025;
  assign n13021 = ~n13045;
  assign n13041 = n9246 & n13046;
  assign n11851 = ~n13047;
  assign n13039 = ~n13052;
  assign n13048 = n13068 & n13069;
  assign n12984 = n13001 ^ n13002;
  assign n13011 = n13016 & n13017;
  assign n13012 = n12960 & n13018;
  assign n12966 = ~n13019;
  assign n13015 = n13026 & n13027;
  assign n13013 = ~n12960;
  assign n13020 = n13039 & n13040;
  assign n11827 = ~n13041;
  assign n9212 = n13048 ^ n13049;
  assign n13050 = ~n13048;
  assign n12415 = n12983 ^ n12984;
  assign n12957 = n12984 & n12983;
  assign n12986 = ~n13011;
  assign n12962 = ~n13012;
  assign n13006 = n13013 & n12979;
  assign n13003 = ~n13015;
  assign n13005 = n13020 ^ n13021;
  assign n13022 = ~n13020;
  assign n13029 = n9212 & n13034;
  assign n9183 = ~n9212;
  assign n13042 = n13050 & n13051;
  assign n12402 = ~n12415;
  assign n12975 = n12986 & n12966;
  assign n12976 = n13003 & n13004;
  assign n12997 = n13005 & n343;
  assign n12981 = ~n13006;
  assign n12995 = ~n13005;
  assign n13014 = n13022 & n13023;
  assign n13007 = n9183 & n11709;
  assign n11769 = ~n13029;
  assign n13024 = n9183 & n13030;
  assign n13031 = ~n13042;
  assign n12958 = n12975 ^ n12976;
  assign n12985 = ~n12976;
  assign n12993 = n12995 & n12996;
  assign n12927 = ~n12997;
  assign n12918 = n13007 ^ n10444;
  assign n12998 = ~n13014;
  assign n11796 = ~n13024;
  assign n13008 = n13031 & n13032;
  assign n10889 = n12957 ^ n12958;
  assign n12916 = n12958 & n12957;
  assign n12977 = n12985 & n12986;
  assign n12952 = ~n12993;
  assign n12987 = n12918 & n12994;
  assign n12978 = n12998 & n12999;
  assign n12988 = ~n12918;
  assign n11793 = n11796 & n11769;
  assign n12990 = n13008 ^ n10364;
  assign n13009 = ~n13008;
  assign n10891 = ~n10889;
  assign n12965 = ~n12977;
  assign n12949 = n12952 & n12927;
  assign n12959 = n12978 ^ n12979;
  assign n12921 = ~n12987;
  assign n12982 = n12988 & n12944;
  assign n9118 = n12989 ^ n12990;
  assign n12980 = ~n12978;
  assign n13000 = n13009 & n13010;
  assign n12948 = n12959 ^ n12960;
  assign n12950 = n12965 & n12966;
  assign n12967 = n9118 & n12974;
  assign n12973 = n12980 & n12981;
  assign n12946 = ~n12982;
  assign n9173 = ~n9118;
  assign n12991 = ~n13000;
  assign n12941 = n12948 & n342;
  assign n12925 = n12949 ^ n12950;
  assign n12939 = ~n12948;
  assign n12951 = ~n12950;
  assign n12953 = n9173 & n11659;
  assign n11699 = ~n12967;
  assign n12963 = n9173 & n12968;
  assign n12961 = ~n12973;
  assign n12969 = n12991 & n12992;
  assign n12229 = n12916 ^ n12925;
  assign n12874 = n12925 & n12916;
  assign n12936 = n12939 & n12940;
  assign n12883 = ~n12941;
  assign n12917 = ~n12925;
  assign n12942 = n12951 & n12952;
  assign n12877 = n12953 ^ n10364;
  assign n12943 = n12961 & n12962;
  assign n11730 = ~n12963;
  assign n12954 = n12969 ^ n12970;
  assign n12971 = ~n12969;
  assign n12216 = n12916 ^ n12917;
  assign n12911 = ~n12936;
  assign n12928 = n12877 & n12937;
  assign n12926 = ~n12942;
  assign n12919 = n12943 ^ n12944;
  assign n12929 = ~n12877;
  assign n12947 = n11730 & n11699;
  assign n9101 = n10321 ^ n12954;
  assign n12945 = ~n12943;
  assign n12964 = n12971 & n12972;
  assign n12897 = n12911 & n12883;
  assign n12909 = n12918 ^ n12919;
  assign n12898 = n12926 & n12927;
  assign n12879 = ~n12928;
  assign n12922 = n12929 & n12906;
  assign n12915 = n9101 & n11574;
  assign n12931 = n9101 & n11677;
  assign n12938 = n12945 & n12946;
  assign n11728 = ~n12947;
  assign n9135 = ~n9101;
  assign n12955 = ~n12964;
  assign n12875 = n12897 ^ n12898;
  assign n12901 = n12909 & n341;
  assign n12899 = ~n12909;
  assign n12903 = n12915 ^ n10321;
  assign n12910 = ~n12898;
  assign n12908 = ~n12922;
  assign n12923 = n9135 & n12930;
  assign n11679 = ~n12931;
  assign n12920 = ~n12938;
  assign n12932 = n12955 & n12956;
  assign n11807 = n12874 ^ n12875;
  assign n12825 = n12875 & n12874;
  assign n12891 = n12899 & n12900;
  assign n12841 = ~n12901;
  assign n12894 = n12903 & n12904;
  assign n12902 = n12910 & n12911;
  assign n12892 = ~n12903;
  assign n12905 = n12920 & n12921;
  assign n11651 = ~n12923;
  assign n12912 = n12932 ^ n12933;
  assign n12934 = ~n12932;
  assign n11805 = n11807 ^ n9893;
  assign n11808 = ~n11807;
  assign n12866 = ~n12891;
  assign n12884 = n12892 & n12893;
  assign n12835 = ~n12894;
  assign n12882 = ~n12902;
  assign n12876 = n12905 ^ n12906;
  assign n9094 = n12912 ^ n10315;
  assign n12907 = ~n12905;
  assign n12924 = n12934 & n12935;
  assign n12813 = n11805 & n11790;
  assign n8831 = ~n11805;
  assign n11834 = n11808 & n9893;
  assign n12873 = n12866 & n12841;
  assign n12864 = n12876 ^ n12877;
  assign n12851 = n12882 & n12883;
  assign n12861 = ~n12884;
  assign n12886 = n9094 & n12896;
  assign n12895 = n12907 & n12908;
  assign n9086 = ~n9094;
  assign n12913 = ~n12924;
  assign n12789 = n12813 ^ n12814;
  assign n12833 = n11834 & n9836;
  assign n11820 = ~n11834;
  assign n12858 = n12864 & n340;
  assign n12852 = ~n12873;
  assign n12856 = ~n12864;
  assign n12867 = n12861 & n12835;
  assign n12865 = ~n12851;
  assign n12868 = n9086 & n11516;
  assign n12880 = n9086 & n12885;
  assign n11586 = ~n12886;
  assign n12878 = ~n12895;
  assign n12888 = n12913 & n12914;
  assign n10387 = n39 ^ n12789;
  assign n12535 = n12789 & n39;
  assign n12790 = ~n12789;
  assign n12824 = n11820 & n9828;
  assign n12780 = ~n12833;
  assign n12826 = n12851 ^ n12852;
  assign n12853 = n12856 & n12857;
  assign n12793 = ~n12858;
  assign n12859 = n12865 & n12866;
  assign n12843 = ~n12867;
  assign n12809 = n12868 ^ n10315;
  assign n12842 = n12878 & n12879;
  assign n11615 = ~n12880;
  assign n9067 = n12887 ^ n12888;
  assign n12889 = ~n12888;
  assign n11599 = ~n10387;
  assign n12643 = n12790 & n12791;
  assign n12803 = ~n12824;
  assign n12800 = n12825 ^ n12826;
  assign n12827 = ~n12826;
  assign n12828 = n12842 ^ n12843;
  assign n12816 = ~n12853;
  assign n12846 = n12809 & n12784;
  assign n12840 = ~n12859;
  assign n12844 = ~n12809;
  assign n12862 = n11615 & n11586;
  assign n12860 = ~n12842;
  assign n12855 = n9067 & n11342;
  assign n12869 = n9067 & n11517;
  assign n8994 = ~n9067;
  assign n12881 = n12889 & n12890;
  assign n12776 = n11834 ^ n12800;
  assign n12801 = n12803 & n12800;
  assign n12781 = n12827 & n12825;
  assign n12819 = n12828 & n339;
  assign n12804 = n12816 & n12793;
  assign n12817 = ~n12828;
  assign n12805 = n12840 & n12841;
  assign n12836 = n12844 & n12845;
  assign n12811 = ~n12846;
  assign n12837 = n12855 ^ n10291;
  assign n12854 = n12860 & n12861;
  assign n11613 = ~n12862;
  assign n11551 = ~n12869;
  assign n12863 = n8994 & n12870;
  assign n12871 = ~n12881;
  assign n8699 = n12776 ^ n9828;
  assign n12779 = ~n12801;
  assign n12782 = n12804 ^ n12805;
  assign n12807 = n12817 & n12818;
  assign n12744 = ~n12819;
  assign n12815 = ~n12805;
  assign n12787 = ~n12836;
  assign n12831 = n12837 & n12838;
  assign n12829 = ~n12837;
  assign n12834 = ~n12854;
  assign n11520 = ~n12863;
  assign n12847 = n12871 & n12872;
  assign n12728 = n8699 & n11759;
  assign n8712 = ~n8699;
  assign n12694 = n12779 & n12780;
  assign n12766 = n12781 ^ n12782;
  assign n12731 = n12782 & n12781;
  assign n12769 = ~n12807;
  assign n12806 = n12815 & n12816;
  assign n12820 = n12829 & n12830;
  assign n12737 = ~n12831;
  assign n12808 = n12834 & n12835;
  assign n9006 = n12847 ^ n12848;
  assign n12849 = ~n12847;
  assign n12710 = n12728 ^ n9828;
  assign n12753 = n12766 & n9811;
  assign n12741 = ~n12694;
  assign n12754 = ~n12766;
  assign n12742 = ~n12731;
  assign n12785 = n12769 & n12744;
  assign n12792 = ~n12806;
  assign n12783 = n12808 ^ n12809;
  assign n12763 = ~n12820;
  assign n12810 = ~n12808;
  assign n12821 = n9006 & n12832;
  assign n8999 = ~n9006;
  assign n12839 = n12849 & n12850;
  assign n12701 = n12710 & n12711;
  assign n12699 = ~n12710;
  assign n12730 = ~n12753;
  assign n12749 = n12754 & n9786;
  assign n12685 = n12783 ^ n12784;
  assign n12758 = ~n12785;
  assign n12757 = n12792 & n12793;
  assign n12794 = n12763 & n12737;
  assign n12802 = n12810 & n12811;
  assign n12795 = n8999 & n11329;
  assign n11448 = ~n12821;
  assign n12812 = n8999 & n11478;
  assign n12822 = ~n12839;
  assign n12693 = n12699 & n12700;
  assign n12645 = ~n12701;
  assign n12729 = n12730 & n12741;
  assign n12713 = ~n12749;
  assign n12732 = n12757 ^ n12758;
  assign n12755 = n12685 & n12767;
  assign n12756 = ~n12685;
  assign n12768 = ~n12757;
  assign n12761 = ~n12794;
  assign n12674 = n12795 ^ n10182;
  assign n12786 = ~n12802;
  assign n11480 = ~n12812;
  assign n12797 = n12822 & n12823;
  assign n12671 = ~n12693;
  assign n12712 = ~n12729;
  assign n12722 = n12713 & n12730;
  assign n12681 = n12731 ^ n12732;
  assign n12657 = n12732 & n12742;
  assign n12716 = ~n12755;
  assign n12750 = n12756 & n338;
  assign n12759 = n12768 & n12769;
  assign n12770 = n12674 & n12777;
  assign n12760 = n12786 & n12787;
  assign n12771 = ~n12674;
  assign n8935 = n12796 ^ n12797;
  assign n12798 = ~n12797;
  assign n12668 = n12671 & n12643;
  assign n12642 = n12671 & n12645;
  assign n12680 = n12712 & n12713;
  assign n12703 = n12681 & n9775;
  assign n12695 = ~n12722;
  assign n12702 = ~n12681;
  assign n12660 = ~n12657;
  assign n12687 = ~n12750;
  assign n12743 = ~n12759;
  assign n12627 = n12760 ^ n12761;
  assign n12676 = ~n12770;
  assign n12764 = n12771 & n12706;
  assign n12762 = ~n12760;
  assign n12752 = n8935 & n11303;
  assign n12773 = n8935 & n12778;
  assign n8983 = ~n8935;
  assign n12788 = n12798 & n12799;
  assign n12623 = n12642 ^ n12643;
  assign n12644 = ~n12668;
  assign n12654 = n12680 ^ n12681;
  assign n8670 = n12694 ^ n12695;
  assign n12682 = ~n12680;
  assign n12696 = n12702 & n9742;
  assign n12683 = ~n12703;
  assign n12714 = n12743 & n12744;
  assign n12735 = n12627 & n337;
  assign n12733 = ~n12627;
  assign n12738 = n12752 ^ n10123;
  assign n12751 = n12762 & n12763;
  assign n12708 = ~n12764;
  assign n12765 = n8983 & n12772;
  assign n11401 = ~n12773;
  assign n12774 = ~n12788;
  assign n12611 = n12623 & n38;
  assign n12609 = ~n12623;
  assign n12603 = n12644 & n12645;
  assign n8613 = n12654 ^ n9742;
  assign n12672 = n12682 & n12683;
  assign n8664 = ~n8670;
  assign n12656 = ~n12696;
  assign n12684 = n338 ^ n12714;
  assign n12715 = ~n12714;
  assign n12723 = n12733 & n12734;
  assign n12629 = ~n12735;
  assign n12726 = n12738 & n12739;
  assign n12724 = ~n12738;
  assign n12736 = ~n12751;
  assign n11358 = ~n12765;
  assign n12746 = n12774 & n12775;
  assign n12602 = n12609 & n12610;
  assign n12537 = ~n12611;
  assign n12614 = n12603 & n12565;
  assign n12612 = ~n12603;
  assign n8603 = ~n8613;
  assign n12637 = n8664 & n11617;
  assign n12655 = ~n12672;
  assign n12658 = n12684 ^ n12685;
  assign n12704 = n12715 & n12716;
  assign n12663 = ~n12723;
  assign n12717 = n12724 & n12725;
  assign n12620 = ~n12726;
  assign n12705 = n12736 & n12737;
  assign n11398 = n11401 & n11358;
  assign n8898 = n12745 ^ n12746;
  assign n12747 = ~n12746;
  assign n12577 = ~n12602;
  assign n12605 = n12612 & n12613;
  assign n12588 = ~n12614;
  assign n12590 = n8603 & n11471;
  assign n12604 = n12637 ^ n9786;
  assign n12539 = n12655 & n12656;
  assign n12638 = n12657 ^ n12658;
  assign n12659 = ~n12658;
  assign n12686 = ~n12704;
  assign n12673 = n12705 ^ n12706;
  assign n12653 = ~n12717;
  assign n12707 = ~n12705;
  assign n12698 = n8898 & n11209;
  assign n12718 = n8898 & n12727;
  assign n8945 = ~n8898;
  assign n12740 = n12747 & n12748;
  assign n12566 = n12577 & n12535;
  assign n12534 = n12577 & n12537;
  assign n12567 = n12590 ^ n9775;
  assign n12564 = n12603 ^ n12604;
  assign n12549 = ~n12605;
  assign n12589 = ~n12604;
  assign n12625 = n12638 & n9707;
  assign n12606 = ~n12539;
  assign n12624 = ~n12638;
  assign n12593 = n12659 & n12660;
  assign n12596 = n12673 ^ n12674;
  assign n12661 = n12686 & n12687;
  assign n12688 = n12653 & n12620;
  assign n12584 = n12698 ^ n10177;
  assign n12697 = n12707 & n12708;
  assign n11316 = ~n12718;
  assign n12709 = n8945 & n12719;
  assign n12720 = ~n12740;
  assign n12496 = n12534 ^ n12535;
  assign n12461 = n12564 ^ n12565;
  assign n12536 = ~n12566;
  assign n12552 = n12567 & n12568;
  assign n12550 = ~n12567;
  assign n12578 = n12588 & n12589;
  assign n12615 = n12624 & n9732;
  assign n12592 = ~n12625;
  assign n12648 = n12596 & n336;
  assign n12626 = n337 ^ n12661;
  assign n12646 = ~n12596;
  assign n12662 = ~n12661;
  assign n12670 = n12584 & n12677;
  assign n12651 = ~n12688;
  assign n12669 = ~n12584;
  assign n12675 = ~n12697;
  assign n11269 = ~n12709;
  assign n12689 = n12720 & n12721;
  assign n11476 = n12496 ^ n10387;
  assign n12416 = n12496 & n10387;
  assign n12526 = n12461 & n12533;
  assign n12499 = n12536 & n12537;
  assign n12527 = ~n12461;
  assign n12538 = n12550 & n12551;
  assign n12473 = ~n12552;
  assign n12548 = ~n12578;
  assign n12591 = n12592 & n12606;
  assign n12570 = ~n12615;
  assign n12594 = n12626 ^ n12627;
  assign n12639 = n12646 & n12647;
  assign n12556 = ~n12648;
  assign n12649 = n12662 & n12663;
  assign n12664 = n12669 & n12543;
  assign n12586 = ~n12670;
  assign n12650 = n12675 & n12676;
  assign n12678 = n11316 & n11269;
  assign n12665 = n12689 ^ n12690;
  assign n12691 = ~n12689;
  assign n11490 = ~n11476;
  assign n12460 = n37 ^ n12499;
  assign n12497 = ~n12526;
  assign n12510 = n12527 & n37;
  assign n12498 = ~n12499;
  assign n12511 = ~n12538;
  assign n12464 = n12548 & n12549;
  assign n12569 = ~n12591;
  assign n12579 = n12592 & n12570;
  assign n12571 = n12593 ^ n12594;
  assign n12514 = n12594 & n12593;
  assign n12598 = ~n12639;
  assign n12628 = ~n12649;
  assign n12630 = n12650 ^ n12651;
  assign n12545 = ~n12664;
  assign n8854 = n10127 ^ n12665;
  assign n12652 = ~n12650;
  assign n11314 = ~n12678;
  assign n12679 = n12691 & n12692;
  assign n12417 = n12460 ^ n12461;
  assign n12486 = n12497 & n12498;
  assign n12463 = ~n12510;
  assign n12501 = n12473 & n12511;
  assign n12512 = ~n12464;
  assign n12528 = n12569 & n12570;
  assign n12553 = n12571 & n9719;
  assign n12540 = ~n12579;
  assign n12487 = ~n12571;
  assign n12595 = n12628 & n12629;
  assign n12618 = n12630 & n351;
  assign n12616 = ~n12630;
  assign n12608 = n8854 & n11126;
  assign n12632 = n8854 & n12641;
  assign n12640 = n12652 & n12653;
  assign n8891 = ~n8854;
  assign n12666 = ~n12679;
  assign n11419 = n12416 ^ n12417;
  assign n12278 = n12417 & n12416;
  assign n12462 = ~n12486;
  assign n12465 = ~n12501;
  assign n12500 = n12511 & n12512;
  assign n12488 = n12528 ^ n9729;
  assign n8517 = n12539 ^ n12540;
  assign n12530 = ~n12528;
  assign n12541 = n12487 & n9729;
  assign n12529 = ~n12553;
  assign n12554 = n12595 ^ n12596;
  assign n12581 = n12608 ^ n10114;
  assign n12597 = ~n12595;
  assign n12607 = n12616 & n12617;
  assign n12478 = ~n12618;
  assign n12621 = n8891 & n12631;
  assign n11234 = ~n12632;
  assign n12619 = ~n12640;
  assign n12633 = n12666 & n12667;
  assign n11397 = ~n11419;
  assign n12329 = n12462 & n12463;
  assign n12436 = n12464 ^ n12465;
  assign n8500 = n12487 ^ n12488;
  assign n12472 = ~n12500;
  assign n12513 = n12529 & n12530;
  assign n8543 = ~n8517;
  assign n12490 = ~n12541;
  assign n12515 = n336 ^ n12554;
  assign n12572 = n12581 & n12582;
  assign n12580 = n12597 & n12598;
  assign n12573 = ~n12581;
  assign n12520 = ~n12607;
  assign n12583 = n12619 & n12620;
  assign n11192 = ~n12621;
  assign n12599 = n12633 ^ n12634;
  assign n12635 = ~n12633;
  assign n12420 = n12436 & n36;
  assign n12383 = ~n12329;
  assign n12418 = ~n12436;
  assign n12421 = n8500 & n11403;
  assign n12422 = n12472 & n12473;
  assign n8505 = ~n8500;
  assign n12466 = n8543 & n11463;
  assign n12489 = ~n12513;
  assign n12491 = n12514 ^ n12515;
  assign n12475 = n12515 & n12514;
  assign n12469 = ~n12572;
  assign n12557 = n12573 & n12574;
  assign n12555 = ~n12580;
  assign n12517 = n12520 & n12478;
  assign n12542 = n12583 ^ n12584;
  assign n12587 = n11234 & n11192;
  assign n8800 = n10093 ^ n12599;
  assign n12585 = ~n12583;
  assign n12622 = n12635 & n12636;
  assign n12408 = n12418 & n12419;
  assign n12346 = ~n12420;
  assign n12311 = n12421 ^ n9719;
  assign n12398 = ~n12422;
  assign n12423 = n12466 ^ n9732;
  assign n12453 = n12489 & n12490;
  assign n12474 = n12491 & n9689;
  assign n12409 = ~n12491;
  assign n12516 = n12542 ^ n12543;
  assign n12518 = n12555 & n12556;
  assign n12508 = ~n12557;
  assign n12531 = n8800 & n11052;
  assign n12558 = n8800 & n12576;
  assign n12575 = n12585 & n12586;
  assign n11232 = ~n12587;
  assign n8843 = ~n8800;
  assign n12600 = ~n12622;
  assign n12384 = n12311 & n12265;
  assign n12382 = ~n12408;
  assign n12385 = ~n12311;
  assign n12380 = n12422 ^ n12423;
  assign n12425 = n12423 & n12437;
  assign n12410 = n12453 ^ n9689;
  assign n12424 = ~n12423;
  assign n12455 = ~n12453;
  assign n12467 = n12409 & n9639;
  assign n12454 = ~n12474;
  assign n12504 = n12516 & n350;
  assign n12476 = n12517 ^ n12518;
  assign n12502 = ~n12516;
  assign n12521 = n12508 & n12469;
  assign n12432 = n12531 ^ n10093;
  assign n12519 = ~n12518;
  assign n11148 = ~n12558;
  assign n12546 = n8843 & n12559;
  assign n12544 = ~n12575;
  assign n12560 = n12600 & n12601;
  assign n12294 = n12380 ^ n12381;
  assign n12374 = n12382 & n12383;
  assign n12375 = n12382 & n12346;
  assign n12281 = ~n12384;
  assign n12376 = n12385 & n12386;
  assign n8410 = n12409 ^ n12410;
  assign n12411 = n12424 & n12381;
  assign n12399 = ~n12425;
  assign n12438 = n12454 & n12455;
  assign n12413 = ~n12467;
  assign n12456 = n12475 ^ n12476;
  assign n12389 = n12476 & n12475;
  assign n12492 = n12502 & n12503;
  assign n12401 = ~n12504;
  assign n12494 = n12432 & n12506;
  assign n12505 = n12519 & n12520;
  assign n12480 = ~n12521;
  assign n12493 = ~n12432;
  assign n12479 = n12544 & n12545;
  assign n11106 = ~n12546;
  assign n8714 = n12560 ^ n12561;
  assign n12562 = ~n12560;
  assign n12344 = n12294 & n35;
  assign n12342 = ~n12294;
  assign n12345 = ~n12374;
  assign n12330 = ~n12375;
  assign n12318 = ~n12376;
  assign n12387 = n12398 & n12399;
  assign n8475 = ~n8410;
  assign n12363 = ~n12411;
  assign n12412 = ~n12438;
  assign n12440 = n12456 & n9633;
  assign n12439 = ~n12456;
  assign n12457 = n12479 ^ n12480;
  assign n12442 = ~n12492;
  assign n12481 = n12493 & n12392;
  assign n12434 = ~n12494;
  assign n12477 = ~n12505;
  assign n11145 = n11148 & n11106;
  assign n12507 = ~n12479;
  assign n12522 = n8714 & n12532;
  assign n8818 = ~n8714;
  assign n12547 = n12562 & n12563;
  assign n12291 = n12329 ^ n12330;
  assign n12328 = n12342 & n12343;
  assign n12263 = ~n12344;
  assign n12331 = n12345 & n12346;
  assign n12332 = n8475 & n11310;
  assign n12362 = ~n12387;
  assign n12348 = n12412 & n12413;
  assign n12426 = n12439 & n9644;
  assign n12378 = ~n12440;
  assign n12445 = n12457 & n349;
  assign n12427 = n12442 & n12401;
  assign n12443 = ~n12457;
  assign n12428 = n12477 & n12478;
  assign n12394 = ~n12481;
  assign n12495 = n12507 & n12508;
  assign n12482 = n8818 & n10957;
  assign n11022 = ~n12522;
  assign n12509 = n8818 & n12523;
  assign n12524 = ~n12547;
  assign n11355 = n12278 ^ n12291;
  assign n12218 = n12291 & n12278;
  assign n12279 = ~n12291;
  assign n12306 = ~n12328;
  assign n12293 = ~n12331;
  assign n12307 = n12332 ^ n9689;
  assign n12347 = n12362 & n12363;
  assign n12377 = ~n12348;
  assign n12334 = ~n12426;
  assign n12390 = n12427 ^ n12428;
  assign n12430 = n12443 & n12444;
  assign n12322 = ~n12445;
  assign n12441 = ~n12428;
  assign n12458 = n12482 ^ n9979;
  assign n12468 = ~n12495;
  assign n11069 = ~n12509;
  assign n12483 = n12524 & n12525;
  assign n11369 = n12278 ^ n12279;
  assign n12221 = ~n12218;
  assign n12254 = n12293 ^ n12294;
  assign n12292 = n12306 & n12293;
  assign n12295 = n12307 & n12308;
  assign n12296 = ~n12307;
  assign n12310 = ~n12347;
  assign n12364 = n12377 & n12378;
  assign n12365 = n12389 ^ n12390;
  assign n12388 = n12378 & n12334;
  assign n12319 = n12390 & n12389;
  assign n12370 = ~n12430;
  assign n12429 = n12441 & n12442;
  assign n12446 = n12458 & n12459;
  assign n12431 = n12468 & n12469;
  assign n12447 = ~n12458;
  assign n12470 = n11069 & n11022;
  assign n12449 = n12483 ^ n10006;
  assign n12484 = ~n12483;
  assign n12219 = n35 ^ n12254;
  assign n12262 = ~n12292;
  assign n12208 = ~n12295;
  assign n12282 = n12296 & n12297;
  assign n12264 = n12310 ^ n12311;
  assign n12309 = n12318 & n12310;
  assign n12333 = ~n12364;
  assign n12350 = n12365 & n9626;
  assign n12299 = ~n12365;
  assign n12349 = ~n12388;
  assign n12367 = n12370 & n12322;
  assign n12400 = ~n12429;
  assign n12391 = n12431 ^ n12432;
  assign n12316 = ~n12446;
  assign n12435 = n12447 & n12448;
  assign n8718 = n12449 ^ n12450;
  assign n12433 = ~n12431;
  assign n11067 = ~n12470;
  assign n12471 = n12484 & n12485;
  assign n11267 = n12218 ^ n12219;
  assign n12220 = ~n12219;
  assign n12160 = n12262 & n12263;
  assign n12243 = n12264 ^ n12265;
  assign n12244 = ~n12282;
  assign n12280 = ~n12309;
  assign n12298 = n12333 & n12334;
  assign n8438 = n12348 ^ n12349;
  assign n12335 = n12299 & n9565;
  assign n12301 = ~n12350;
  assign n12366 = n12391 ^ n12392;
  assign n12368 = n12400 & n12401;
  assign n12379 = n8718 & n10863;
  assign n12403 = n8718 & n12415;
  assign n12414 = n12433 & n12434;
  assign n12359 = ~n12435;
  assign n8725 = ~n8718;
  assign n12451 = ~n12471;
  assign n11287 = ~n11267;
  assign n12126 = n12220 & n12221;
  assign n12232 = n12243 & n34;
  assign n12193 = ~n12160;
  assign n12246 = n12244 & n12208;
  assign n12230 = ~n12243;
  assign n12205 = n12280 & n12281;
  assign n12255 = n12298 ^ n12299;
  assign n12300 = ~n12298;
  assign n8429 = ~n8438;
  assign n12257 = ~n12335;
  assign n12353 = n12366 & n348;
  assign n12320 = n12367 ^ n12368;
  assign n12351 = ~n12366;
  assign n12274 = n12379 ^ n9923;
  assign n12369 = ~n12368;
  assign n12395 = n12359 & n12316;
  assign n12396 = n8725 & n12402;
  assign n10983 = ~n12403;
  assign n12393 = ~n12414;
  assign n12404 = n12451 & n12452;
  assign n12129 = ~n12126;
  assign n12222 = n12230 & n12231;
  assign n12162 = ~n12232;
  assign n12206 = ~n12246;
  assign n8376 = n12255 ^ n9565;
  assign n12245 = ~n12205;
  assign n12283 = n12300 & n12301;
  assign n12266 = n8429 & n11218;
  assign n12225 = n12319 ^ n12320;
  assign n12237 = n12320 & n12319;
  assign n12336 = n12351 & n12352;
  assign n12250 = ~n12353;
  assign n12337 = n12274 & n12355;
  assign n12354 = n12369 & n12370;
  assign n12338 = ~n12274;
  assign n12356 = n12393 & n12394;
  assign n12357 = ~n12395;
  assign n10938 = ~n12396;
  assign n12372 = n12404 ^ n9946;
  assign n12407 = n12404 & n12371;
  assign n12405 = ~n12404;
  assign n12183 = n12205 ^ n12206;
  assign n12194 = ~n12222;
  assign n12195 = n8376 & n11132;
  assign n12233 = n12244 & n12245;
  assign n8389 = ~n8376;
  assign n12247 = n12266 ^ n9633;
  assign n12256 = ~n12283;
  assign n12285 = n12225 & n9590;
  assign n12284 = ~n12225;
  assign n12287 = ~n12336;
  assign n12276 = ~n12337;
  assign n12324 = n12338 & n12240;
  assign n12321 = ~n12354;
  assign n12323 = n12356 ^ n12357;
  assign n12360 = n10983 & n10938;
  assign n8709 = n12371 ^ n12372;
  assign n12358 = ~n12356;
  assign n12397 = n12405 & n12406;
  assign n12327 = ~n12407;
  assign n12172 = n12183 & n33;
  assign n12184 = n12193 & n12194;
  assign n12159 = n12194 & n12162;
  assign n12084 = n12195 ^ n9626;
  assign n12169 = ~n12183;
  assign n12207 = ~n12233;
  assign n12236 = n12247 & n12248;
  assign n12234 = ~n12247;
  assign n12224 = n12256 & n12257;
  assign n12267 = n12284 & n9523;
  assign n12227 = ~n12285;
  assign n12268 = n12287 & n12250;
  assign n12269 = n12321 & n12322;
  assign n12314 = n12323 & n347;
  assign n12242 = ~n12324;
  assign n12312 = ~n12323;
  assign n12303 = n8709 & n10749;
  assign n12339 = n12358 & n12359;
  assign n10981 = ~n12360;
  assign n8607 = ~n8709;
  assign n12373 = n12327 & n9951;
  assign n12341 = ~n12397;
  assign n12127 = n12159 ^ n12160;
  assign n12163 = n12169 & n12170;
  assign n12164 = n12084 & n12171;
  assign n12104 = ~n12172;
  assign n12161 = ~n12184;
  assign n12165 = ~n12084;
  assign n12150 = n12207 & n12208;
  assign n12185 = n12224 ^ n12225;
  assign n12223 = n12234 & n12235;
  assign n12140 = ~n12236;
  assign n12226 = ~n12224;
  assign n12188 = ~n12267;
  assign n12238 = n12268 ^ n12269;
  assign n12271 = n12303 ^ n9946;
  assign n12286 = ~n12269;
  assign n12302 = n12312 & n12313;
  assign n12178 = ~n12314;
  assign n12315 = ~n12339;
  assign n12361 = n12341 & n9946;
  assign n12340 = ~n12373;
  assign n10169 = n12126 ^ n12127;
  assign n12128 = ~n12127;
  assign n12101 = n12161 & n12162;
  assign n12131 = ~n12163;
  assign n12087 = ~n12164;
  assign n12149 = n12165 & n12110;
  assign n8298 = n12185 ^ n9523;
  assign n12173 = ~n12150;
  assign n12174 = ~n12223;
  assign n12209 = n12226 & n12227;
  assign n12153 = n12237 ^ n12238;
  assign n12175 = n12238 & n12237;
  assign n12258 = n12271 & n12272;
  assign n12270 = n12286 & n12287;
  assign n12259 = ~n12271;
  assign n12214 = ~n12302;
  assign n12273 = n12315 & n12316;
  assign n12325 = n12340 & n12341;
  assign n12326 = ~n12361;
  assign n11190 = ~n10169;
  assign n12072 = n12128 & n12129;
  assign n12132 = n12131 & n12104;
  assign n12130 = ~n12101;
  assign n12112 = ~n12149;
  assign n12166 = n12173 & n12174;
  assign n8360 = ~n8298;
  assign n12186 = n12174 & n12140;
  assign n12187 = ~n12209;
  assign n12196 = n12153 & n9528;
  assign n12197 = ~n12153;
  assign n12168 = ~n12258;
  assign n12251 = n12259 & n12260;
  assign n12249 = ~n12270;
  assign n12211 = n12214 & n12178;
  assign n12239 = n12273 ^ n12274;
  assign n12275 = ~n12273;
  assign n12304 = ~n12325;
  assign n12317 = n12326 & n12327;
  assign n12075 = ~n12072;
  assign n12116 = n12130 & n12131;
  assign n12102 = ~n12132;
  assign n12120 = n8360 & n11063;
  assign n12139 = ~n12166;
  assign n12151 = ~n12186;
  assign n12152 = n12187 & n12188;
  assign n12155 = ~n12196;
  assign n12189 = n12197 & n9534;
  assign n12210 = n12239 ^ n12240;
  assign n12212 = n12249 & n12250;
  assign n12203 = ~n12251;
  assign n12261 = n12275 & n12276;
  assign n12288 = n12304 & n12305;
  assign n12289 = ~n12317;
  assign n12073 = n12101 ^ n12102;
  assign n12103 = ~n12116;
  assign n12035 = n12120 ^ n9590;
  assign n12109 = n12139 & n12140;
  assign n12133 = n12150 ^ n12151;
  assign n12121 = n12152 ^ n12153;
  assign n12154 = ~n12152;
  assign n12123 = ~n12189;
  assign n12200 = n12210 & n346;
  assign n12176 = n12211 ^ n12212;
  assign n12198 = ~n12210;
  assign n12215 = n12203 & n12168;
  assign n12213 = ~n12212;
  assign n12241 = ~n12261;
  assign n12253 = ~n12288;
  assign n12277 = n12289 & n12290;
  assign n11127 = n12072 ^ n12073;
  assign n12074 = ~n12073;
  assign n12066 = n12103 & n12104;
  assign n12095 = n12035 & n12060;
  assign n12085 = n12109 ^ n12110;
  assign n12093 = ~n12035;
  assign n8283 = n12121 ^ n9528;
  assign n12119 = n12133 & n32;
  assign n12111 = ~n12109;
  assign n12117 = ~n12133;
  assign n12141 = n12154 & n12155;
  assign n12097 = n12175 ^ n12176;
  assign n12106 = n12176 & n12175;
  assign n12190 = n12198 & n12199;
  assign n12115 = ~n12200;
  assign n12201 = n12213 & n12214;
  assign n12180 = ~n12215;
  assign n12179 = n12241 & n12242;
  assign n12252 = ~n12277;
  assign n11103 = ~n11127;
  assign n12041 = n12074 & n12075;
  assign n12006 = n12084 ^ n12085;
  assign n12076 = ~n12066;
  assign n12088 = n12093 & n12094;
  assign n12037 = ~n12095;
  assign n12078 = n8283 & n10973;
  assign n12105 = n12111 & n12112;
  assign n8337 = ~n8283;
  assign n12113 = n12117 & n12118;
  assign n12048 = ~n12119;
  assign n12122 = ~n12141;
  assign n12143 = n12097 & n9463;
  assign n12142 = ~n12097;
  assign n12156 = n12179 ^ n12180;
  assign n12145 = ~n12190;
  assign n12177 = ~n12201;
  assign n12202 = ~n12179;
  assign n8586 = n12252 & n12253;
  assign n12058 = n12006 & n47;
  assign n12056 = ~n12006;
  assign n11990 = n12078 ^ n9534;
  assign n12061 = ~n12088;
  assign n12086 = ~n12105;
  assign n12077 = ~n12113;
  assign n12096 = n12122 & n12123;
  assign n12134 = n12142 & n9520;
  assign n12099 = ~n12143;
  assign n12148 = n12156 & n345;
  assign n12135 = n12145 & n12115;
  assign n12146 = ~n12156;
  assign n12136 = n12177 & n12178;
  assign n12191 = n12202 & n12203;
  assign n12192 = n8586 & n12228;
  assign n12217 = n8586 & n12229;
  assign n9929 = ~n8586;
  assign n12046 = n12056 & n12057;
  assign n12008 = ~n12058;
  assign n12049 = n11990 & n12016;
  assign n12050 = ~n11990;
  assign n12067 = n12076 & n12077;
  assign n12059 = n12086 & n12087;
  assign n12065 = n12077 & n12048;
  assign n12068 = n12096 ^ n12097;
  assign n12098 = ~n12096;
  assign n12070 = ~n12134;
  assign n12107 = n12135 ^ n12136;
  assign n12138 = n12146 & n12147;
  assign n12064 = ~n12148;
  assign n12144 = ~n12136;
  assign n12167 = ~n12191;
  assign n12157 = n12192 ^ n9873;
  assign n12204 = n9929 & n12216;
  assign n12182 = ~n12217;
  assign n12028 = ~n12046;
  assign n12018 = ~n12049;
  assign n12043 = n12050 & n12051;
  assign n12034 = n12059 ^ n12060;
  assign n12042 = n12065 ^ n12066;
  assign n12047 = ~n12067;
  assign n8304 = n12068 ^ n9520;
  assign n12062 = ~n12059;
  assign n12089 = n12098 & n12099;
  assign n12090 = n12106 ^ n12107;
  assign n12053 = n12107 & n12106;
  assign n12092 = ~n12138;
  assign n12137 = n12144 & n12145;
  assign n12125 = n12157 ^ n12158;
  assign n12124 = n12167 & n12168;
  assign n12181 = ~n12204;
  assign n11985 = n12034 ^ n12035;
  assign n10107 = n12041 ^ n12042;
  assign n11992 = ~n12043;
  assign n11982 = n12042 & n12041;
  assign n12029 = n12047 & n12048;
  assign n12052 = n12061 & n12062;
  assign n8294 = ~n8304;
  assign n12069 = ~n12089;
  assign n12079 = n12090 & n9472;
  assign n12080 = ~n12090;
  assign n12108 = n12092 & n12064;
  assign n12100 = n12124 ^ n12125;
  assign n12114 = ~n12137;
  assign n10766 = n12181 & n12182;
  assign n12013 = n11985 & n12021;
  assign n12014 = ~n11985;
  assign n12005 = n47 ^ n12029;
  assign n11042 = ~n10107;
  assign n12027 = ~n12029;
  assign n12023 = n8294 & n10882;
  assign n12036 = ~n12052;
  assign n12031 = n12069 & n12070;
  assign n12045 = ~n12079;
  assign n12071 = n12080 & n9481;
  assign n12040 = n344 ^ n12100;
  assign n12082 = ~n12108;
  assign n12081 = n12114 & n12115;
  assign n10784 = ~n10766;
  assign n11983 = n12005 ^ n12006;
  assign n11987 = ~n12013;
  assign n12009 = n12014 & n46;
  assign n12010 = n12023 ^ n9463;
  assign n12022 = n12027 & n12028;
  assign n12015 = n12036 & n12037;
  assign n12044 = ~n12031;
  assign n12025 = ~n12071;
  assign n12054 = n12081 ^ n12082;
  assign n12091 = ~n12081;
  assign n10067 = n11982 ^ n11983;
  assign n11948 = n11983 & n11982;
  assign n11965 = ~n12009;
  assign n11998 = n12010 & n12011;
  assign n11989 = n12015 ^ n12016;
  assign n11999 = ~n12010;
  assign n12007 = ~n12022;
  assign n12017 = ~n12015;
  assign n12038 = n12044 & n12045;
  assign n12030 = n12045 & n12025;
  assign n12002 = n12053 ^ n12054;
  assign n12055 = ~n12054;
  assign n12083 = n12091 & n12092;
  assign n10958 = ~n10067;
  assign n11954 = ~n11948;
  assign n11925 = n11989 ^ n11990;
  assign n11958 = ~n11998;
  assign n11993 = n11999 & n12000;
  assign n11984 = n12007 & n12008;
  assign n12012 = n12017 & n12018;
  assign n8229 = n12030 ^ n12031;
  assign n12024 = ~n12038;
  assign n12033 = n12002 & n9417;
  assign n12032 = ~n12002;
  assign n12019 = n12055 & n12053;
  assign n12063 = ~n12083;
  assign n11969 = n11925 & n11976;
  assign n11963 = n11984 ^ n11985;
  assign n11970 = ~n11925;
  assign n11972 = ~n11993;
  assign n11986 = ~n11984;
  assign n11991 = ~n12012;
  assign n11994 = n8229 & n10728;
  assign n12001 = n12024 & n12025;
  assign n8211 = ~n8229;
  assign n12026 = n12032 & n9409;
  assign n11981 = ~n12033;
  assign n12039 = n12063 & n12064;
  assign n11949 = n46 ^ n11963;
  assign n11951 = ~n11969;
  assign n11966 = n11970 & n45;
  assign n11973 = n11972 & n11958;
  assign n11977 = n11986 & n11987;
  assign n11955 = n11991 & n11992;
  assign n11915 = n11994 ^ n9472;
  assign n11979 = n12001 ^ n12002;
  assign n12003 = ~n12001;
  assign n12004 = ~n12026;
  assign n12020 = n12039 ^ n12040;
  assign n10027 = n11948 ^ n11949;
  assign n11907 = n11949 & n11954;
  assign n11927 = ~n11966;
  assign n11956 = ~n11973;
  assign n11964 = ~n11977;
  assign n11975 = n11915 & n11978;
  assign n8198 = n11979 ^ n9417;
  assign n11971 = ~n11955;
  assign n11974 = ~n11915;
  assign n11995 = n12003 & n12004;
  assign n11945 = n12019 ^ n12020;
  assign n10029 = ~n10027;
  assign n11910 = ~n11907;
  assign n11943 = n11955 ^ n11956;
  assign n11950 = n11964 & n11965;
  assign n11953 = n8198 & n10712;
  assign n11967 = n11971 & n11972;
  assign n11968 = n11974 & n11939;
  assign n11917 = ~n11975;
  assign n8209 = ~n8198;
  assign n11980 = ~n11995;
  assign n11997 = n11945 & n9396;
  assign n11996 = ~n11945;
  assign n11937 = n11943 & n44;
  assign n11924 = n45 ^ n11950;
  assign n11935 = n11953 ^ n9409;
  assign n11933 = ~n11943;
  assign n11952 = ~n11950;
  assign n11957 = ~n11967;
  assign n11941 = ~n11968;
  assign n11960 = n11980 & n11981;
  assign n11988 = n11996 & n9323;
  assign n11962 = ~n11997;
  assign n11908 = n11924 ^ n11925;
  assign n11928 = n11933 & n11934;
  assign n11929 = n11935 & n11936;
  assign n11888 = ~n11937;
  assign n11930 = ~n11935;
  assign n11942 = n11951 & n11952;
  assign n11938 = n11957 & n11958;
  assign n11944 = n11960 ^ n9396;
  assign n11961 = ~n11960;
  assign n11947 = ~n11988;
  assign n10671 = n11907 ^ n11908;
  assign n11909 = ~n11908;
  assign n11912 = ~n11928;
  assign n11878 = ~n11929;
  assign n11919 = n11930 & n11931;
  assign n11914 = n11938 ^ n11939;
  assign n11926 = ~n11942;
  assign n8176 = n11944 ^ n11945;
  assign n11940 = ~n11938;
  assign n11959 = n11961 & n11962;
  assign n11875 = n11909 & n11910;
  assign n11901 = n11914 ^ n11915;
  assign n11897 = n11912 & n11888;
  assign n11900 = ~n11919;
  assign n11898 = n11926 & n11927;
  assign n11913 = n8176 & n10626;
  assign n11932 = n11940 & n11941;
  assign n8189 = ~n8176;
  assign n11946 = ~n11959;
  assign n11876 = n11897 ^ n11898;
  assign n11896 = n11901 & n43;
  assign n11894 = ~n11901;
  assign n11903 = n11900 & n11878;
  assign n11838 = n11913 ^ n9323;
  assign n11911 = ~n11898;
  assign n11916 = ~n11932;
  assign n11920 = n11946 & n11947;
  assign n9930 = n11875 ^ n11876;
  assign n11835 = n11876 & n11875;
  assign n11889 = n11894 & n11895;
  assign n11853 = ~n11896;
  assign n11892 = n11838 & n11862;
  assign n11881 = ~n11903;
  assign n11890 = ~n11838;
  assign n11902 = n11911 & n11912;
  assign n11880 = n11916 & n11917;
  assign n11904 = n11920 ^ n11921;
  assign n11922 = ~n11920;
  assign n7817 = n11805 ^ n9930;
  assign n9900 = n11808 ^ n9930;
  assign n11857 = ~n9930;
  assign n11874 = n11880 ^ n11881;
  assign n11873 = ~n11889;
  assign n11882 = n11890 & n11891;
  assign n11864 = ~n11892;
  assign n11887 = ~n11902;
  assign n8146 = n11904 ^ n9283;
  assign n11899 = ~n11880;
  assign n11918 = n11922 & n11923;
  assign n9899 = ~n7817;
  assign n11748 = n11857 & n8831;
  assign n11868 = n11874 & n42;
  assign n11858 = n11873 & n11853;
  assign n11866 = ~n11874;
  assign n11841 = ~n11882;
  assign n11859 = n11887 & n11888;
  assign n11893 = n11899 & n11900;
  assign n8137 = ~n8146;
  assign n11905 = ~n11918;
  assign n11804 = n9899 & n9893;
  assign n11828 = n9899 & n11834;
  assign n11836 = n11858 ^ n11859;
  assign n11860 = n11866 & n11867;
  assign n11801 = ~n11868;
  assign n11872 = ~n11859;
  assign n11869 = n8137 & n10559;
  assign n11877 = ~n11893;
  assign n11884 = n11905 & n11906;
  assign n11789 = n11804 ^ n11805;
  assign n11809 = n11804 & n11820;
  assign n11806 = ~n11804;
  assign n11777 = ~n11828;
  assign n11821 = n11835 ^ n11836;
  assign n11782 = n11836 & n11835;
  assign n11830 = ~n11860;
  assign n11817 = n11869 ^ n9283;
  assign n11865 = n11872 & n11873;
  assign n11861 = n11877 & n11878;
  assign n8048 = n11883 ^ n11884;
  assign n11885 = ~n11884;
  assign n11758 = n11789 & n11790;
  assign n11797 = n11806 & n11807;
  assign n11798 = n11777 & n11808;
  assign n11779 = ~n11809;
  assign n11810 = n11821 & n8699;
  assign n11811 = ~n11821;
  assign n11791 = ~n11782;
  assign n11839 = n11830 & n11801;
  assign n11846 = n11817 & n11854;
  assign n11837 = n11861 ^ n11862;
  assign n11847 = ~n11817;
  assign n11852 = ~n11865;
  assign n11863 = ~n11861;
  assign n11856 = n8048 & n10539;
  assign n8095 = ~n8048;
  assign n11879 = n11885 & n11886;
  assign n11660 = n11758 ^ n11759;
  assign n11762 = n11758 & n11759;
  assign n11760 = ~n11758;
  assign n11776 = ~n11797;
  assign n11778 = ~n11798;
  assign n11781 = ~n11810;
  assign n11799 = n11811 & n8712;
  assign n11773 = n11837 ^ n11838;
  assign n11815 = ~n11839;
  assign n11818 = ~n11846;
  assign n11844 = n11847 & n11785;
  assign n11814 = n11852 & n11853;
  assign n11842 = n11856 ^ n9288;
  assign n11855 = n11863 & n11864;
  assign n11870 = ~n11879;
  assign n11742 = n11760 & n11761;
  assign n11642 = ~n11762;
  assign n11770 = n11776 & n11777;
  assign n11771 = n11778 & n11779;
  assign n11780 = n11781 & n11748;
  assign n11764 = ~n11799;
  assign n11783 = n11814 ^ n11815;
  assign n11812 = n11773 & n11822;
  assign n11813 = ~n11773;
  assign n11833 = n11842 & n11843;
  assign n11787 = ~n11844;
  assign n11829 = ~n11814;
  assign n11831 = ~n11842;
  assign n11840 = ~n11855;
  assign n11848 = n11870 & n11871;
  assign n11671 = ~n11742;
  assign n11743 = ~n11770;
  assign n11745 = ~n11771;
  assign n11763 = ~n11780;
  assign n11747 = n11764 & n11781;
  assign n11721 = n11782 ^ n11783;
  assign n11700 = n11783 & n11791;
  assign n11775 = ~n11812;
  assign n11802 = n11813 & n41;
  assign n11823 = n11829 & n11830;
  assign n11824 = n11831 & n11832;
  assign n11717 = ~n11833;
  assign n11816 = n11840 & n11841;
  assign n11825 = n11848 ^ n11849;
  assign n11850 = ~n11848;
  assign n11731 = n11743 & n11744;
  assign n11732 = n11745 & n11746;
  assign n7642 = n11747 ^ n11748;
  assign n11720 = n11763 & n11764;
  assign n11750 = n11721 & n8664;
  assign n11749 = ~n11721;
  assign n11703 = ~n11700;
  assign n11736 = ~n11802;
  assign n11784 = n11816 ^ n11817;
  assign n11800 = ~n11823;
  assign n11757 = ~n11824;
  assign n8061 = n11825 ^ n9246;
  assign n11819 = ~n11816;
  assign n11845 = n11850 & n11851;
  assign n11693 = n11720 ^ n11721;
  assign n11710 = ~n11731;
  assign n11711 = ~n11732;
  assign n7792 = ~n7642;
  assign n11722 = ~n11720;
  assign n11734 = n11749 & n8670;
  assign n11723 = ~n11750;
  assign n11765 = n11784 ^ n11785;
  assign n11772 = n11800 & n11801;
  assign n11792 = n11757 & n11717;
  assign n11803 = n11818 & n11819;
  assign n8054 = ~n8061;
  assign n11826 = ~n11845;
  assign n7634 = n11693 ^ n8670;
  assign n11685 = n11710 & n11711;
  assign n11686 = n7792 & n9836;
  assign n11712 = n11722 & n11723;
  assign n11695 = ~n11734;
  assign n11753 = n11765 & n40;
  assign n11733 = n11772 ^ n11773;
  assign n11751 = ~n11765;
  assign n11774 = ~n11772;
  assign n11755 = ~n11792;
  assign n11767 = n8054 & n10420;
  assign n11786 = ~n11803;
  assign n11794 = n11826 & n11827;
  assign n7623 = ~n7634;
  assign n11362 = n263 ^ n11685;
  assign n11661 = n11686 ^ n8699;
  assign n11687 = ~n11685;
  assign n11694 = ~n11712;
  assign n11701 = n41 ^ n11733;
  assign n11737 = n11751 & n11752;
  assign n11683 = ~n11753;
  assign n11738 = n11767 ^ n9224;
  assign n11766 = n11774 & n11775;
  assign n11754 = n11786 & n11787;
  assign n7965 = n11793 ^ n11794;
  assign n11795 = ~n11794;
  assign n11639 = n11660 ^ n11661;
  assign n11662 = n11661 & n11671;
  assign n11640 = n7623 & n9786;
  assign n11377 = ~n11362;
  assign n11552 = n11687 & n263;
  assign n11620 = n11694 & n11695;
  assign n11688 = n11700 ^ n11701;
  assign n11702 = ~n11701;
  assign n11705 = ~n11737;
  assign n11724 = n11738 & n11739;
  assign n11655 = n11754 ^ n11755;
  assign n11725 = ~n11738;
  assign n11735 = ~n11766;
  assign n11756 = ~n11754;
  assign n11741 = n7965 & n10401;
  assign n7996 = ~n7965;
  assign n11788 = n11795 & n11796;
  assign n11628 = n11639 & n262;
  assign n11616 = n11640 ^ n8664;
  assign n11626 = ~n11639;
  assign n11641 = ~n11662;
  assign n11680 = n11688 & n8603;
  assign n11663 = ~n11620;
  assign n11681 = ~n11688;
  assign n11664 = n11702 & n11703;
  assign n11689 = n11705 & n11683;
  assign n11715 = n11655 & n55;
  assign n11669 = ~n11724;
  assign n11718 = n11725 & n11726;
  assign n11690 = n11735 & n11736;
  assign n11713 = ~n11655;
  assign n11605 = n11741 ^ n9212;
  assign n11740 = n11756 & n11757;
  assign n11768 = ~n11788;
  assign n11609 = n11616 & n11617;
  assign n11618 = n11626 & n11627;
  assign n11567 = ~n11628;
  assign n11610 = ~n11616;
  assign n11530 = n11641 & n11642;
  assign n11653 = ~n11680;
  assign n11672 = n11681 & n8613;
  assign n11665 = n11689 ^ n11690;
  assign n11667 = ~n11664;
  assign n11706 = n11713 & n11714;
  assign n11624 = ~n11715;
  assign n11707 = n11605 & n11635;
  assign n11692 = ~n11718;
  assign n11704 = ~n11690;
  assign n11708 = ~n11605;
  assign n11716 = ~n11740;
  assign n11727 = n11768 & n11769;
  assign n11544 = ~n11609;
  assign n11601 = n11610 & n11611;
  assign n11600 = ~n11618;
  assign n11581 = ~n11530;
  assign n11652 = n11653 & n11663;
  assign n11643 = n11664 ^ n11665;
  assign n11630 = ~n11672;
  assign n11666 = ~n11665;
  assign n11673 = n11692 & n11669;
  assign n11696 = n11704 & n11705;
  assign n11657 = ~n11706;
  assign n11637 = ~n11707;
  assign n11697 = n11708 & n11709;
  assign n11674 = n11716 & n11717;
  assign n7986 = n11727 ^ n11728;
  assign n11729 = ~n11727;
  assign n11587 = n11600 & n11552;
  assign n11588 = n11600 & n11567;
  assign n11580 = ~n11601;
  assign n11631 = n11643 & n8517;
  assign n11629 = ~n11652;
  assign n11619 = n11630 & n11653;
  assign n11632 = ~n11643;
  assign n11590 = n11666 & n11667;
  assign n11595 = n11673 ^ n11674;
  assign n11682 = ~n11696;
  assign n11607 = ~n11697;
  assign n11691 = ~n11674;
  assign n7976 = ~n7986;
  assign n11719 = n11729 & n11730;
  assign n11565 = n11580 & n11581;
  assign n11568 = n11544 & n11580;
  assign n11566 = ~n11587;
  assign n11553 = ~n11588;
  assign n7553 = n11619 ^ n11620;
  assign n11556 = n11629 & n11630;
  assign n11571 = ~n11631;
  assign n11621 = n11632 & n8543;
  assign n11645 = n11595 & n11658;
  assign n11646 = ~n11595;
  assign n11654 = n11682 & n11683;
  assign n11684 = n11691 & n11692;
  assign n11675 = n7976 & n10366;
  assign n11698 = ~n11719;
  assign n11521 = n11552 ^ n11553;
  assign n11543 = ~n11565;
  assign n11422 = n11566 & n11567;
  assign n11531 = ~n11568;
  assign n11569 = n7553 & n9742;
  assign n7568 = ~n7553;
  assign n11602 = ~n11556;
  assign n11603 = ~n11621;
  assign n11597 = ~n11645;
  assign n11633 = n11646 & n54;
  assign n11622 = n11654 ^ n11655;
  assign n11656 = ~n11654;
  assign n11539 = n11675 ^ n9173;
  assign n11668 = ~n11684;
  assign n11676 = n11698 & n11699;
  assign n11297 = n11521 ^ n11362;
  assign n11370 = n11521 & n11362;
  assign n11507 = n11530 ^ n11531;
  assign n11508 = n11543 & n11544;
  assign n11462 = ~n11422;
  assign n11509 = n11569 ^ n8613;
  assign n11589 = n11602 & n11603;
  assign n11593 = n11603 & n11571;
  assign n11591 = n55 ^ n11622;
  assign n11560 = ~n11633;
  assign n11644 = n11656 & n11657;
  assign n11647 = n11539 & n11659;
  assign n11634 = n11668 & n11669;
  assign n11648 = ~n11539;
  assign n11649 = n11676 ^ n11677;
  assign n11678 = ~n11676;
  assign n11493 = n11507 & n261;
  assign n9682 = ~n11297;
  assign n11470 = n11508 ^ n11509;
  assign n11491 = ~n11507;
  assign n11511 = ~n11508;
  assign n11532 = n11509 & n11545;
  assign n11533 = ~n11509;
  assign n11570 = ~n11589;
  assign n11535 = n11590 ^ n11591;
  assign n11557 = ~n11593;
  assign n11592 = ~n11591;
  assign n11604 = n11634 ^ n11635;
  assign n11623 = ~n11644;
  assign n11541 = ~n11647;
  assign n11638 = n11648 & n11576;
  assign n7909 = n11649 ^ n9101;
  assign n11636 = ~n11634;
  assign n11670 = n11678 & n11679;
  assign n11375 = n11470 ^ n11471;
  assign n11481 = n11491 & n11492;
  assign n11424 = ~n11493;
  assign n11510 = ~n11532;
  assign n11522 = n11533 & n11471;
  assign n7477 = n11556 ^ n11557;
  assign n11534 = n11570 & n11571;
  assign n11555 = n11535 & n8500;
  assign n11554 = ~n11535;
  assign n11524 = n11592 & n11590;
  assign n11527 = n11604 ^ n11605;
  assign n11594 = n11623 & n11624;
  assign n11598 = n7909 & n10289;
  assign n11625 = n11636 & n11637;
  assign n11578 = ~n11638;
  assign n7923 = ~n7909;
  assign n11650 = ~n11670;
  assign n11438 = n11375 & n260;
  assign n11436 = ~n11375;
  assign n11461 = ~n11481;
  assign n11494 = n11510 & n11511;
  assign n11473 = ~n11522;
  assign n11495 = n11534 ^ n11535;
  assign n7463 = ~n7477;
  assign n11536 = ~n11534;
  assign n11546 = n11554 & n8505;
  assign n11537 = ~n11555;
  assign n11572 = n11527 & n11582;
  assign n11558 = n11594 ^ n11595;
  assign n11573 = ~n11527;
  assign n11465 = n11598 ^ n9101;
  assign n11596 = ~n11594;
  assign n11606 = ~n11625;
  assign n11612 = n11650 & n11651;
  assign n11420 = n11436 & n11437;
  assign n11334 = ~n11438;
  assign n11449 = n11461 & n11462;
  assign n11421 = n11461 & n11424;
  assign n11472 = ~n11494;
  assign n7347 = n8500 ^ n11495;
  assign n11482 = n7463 & n9732;
  assign n11523 = n11536 & n11537;
  assign n11497 = ~n11546;
  assign n11525 = n54 ^ n11558;
  assign n11528 = ~n11572;
  assign n11561 = n11573 & n53;
  assign n11562 = n11465 & n11574;
  assign n11563 = ~n11465;
  assign n11583 = n11596 & n11597;
  assign n11575 = n11606 & n11607;
  assign n7808 = n11612 ^ n11613;
  assign n11614 = ~n11612;
  assign n11372 = ~n11420;
  assign n11371 = n11421 ^ n11422;
  assign n11423 = ~n11449;
  assign n11440 = n11472 & n11473;
  assign n11439 = n7347 & n9729;
  assign n7427 = ~n7347;
  assign n11388 = n11482 ^ n8543;
  assign n11496 = ~n11523;
  assign n11498 = n11524 ^ n11525;
  assign n11454 = n11525 & n11524;
  assign n11487 = ~n11561;
  assign n11467 = ~n11562;
  assign n11547 = n11563 & n11503;
  assign n11538 = n11575 ^ n11576;
  assign n11559 = ~n11583;
  assign n11577 = ~n11575;
  assign n11584 = n7808 & n11599;
  assign n7888 = ~n7808;
  assign n11608 = n11614 & n11615;
  assign n11200 = n11370 ^ n11371;
  assign n11288 = n11371 & n11370;
  assign n11374 = n11423 & n11424;
  assign n11402 = n11439 ^ n8500;
  assign n11389 = n11440 ^ n11441;
  assign n11404 = ~n11440;
  assign n11450 = n11388 & n11463;
  assign n11451 = ~n11388;
  assign n11407 = n11496 & n11497;
  assign n11483 = n11498 & n8410;
  assign n11484 = ~n11498;
  assign n11457 = ~n11454;
  assign n11512 = n11538 ^ n11539;
  assign n11505 = ~n11547;
  assign n11526 = n11559 & n11560;
  assign n11564 = n11577 & n11578;
  assign n11548 = n7888 & n10315;
  assign n10371 = ~n11584;
  assign n11579 = n7888 & n10387;
  assign n11585 = ~n11608;
  assign n11220 = ~n11200;
  assign n11332 = n11374 ^ n11375;
  assign n11291 = n11388 ^ n11389;
  assign n11390 = n11402 & n11403;
  assign n11373 = ~n11374;
  assign n11391 = ~n11402;
  assign n11361 = ~n11450;
  assign n11442 = n11451 & n11441;
  assign n11452 = ~n11407;
  assign n11409 = ~n11483;
  assign n11474 = n11484 & n8475;
  assign n11501 = n11512 & n52;
  assign n11485 = n11526 ^ n11527;
  assign n11499 = ~n11512;
  assign n11529 = ~n11526;
  assign n11383 = n11548 ^ n9094;
  assign n11540 = ~n11564;
  assign n10389 = ~n11579;
  assign n11549 = n11585 & n11586;
  assign n11289 = n260 ^ n11332;
  assign n11348 = n11291 & n259;
  assign n11359 = n11372 & n11373;
  assign n11346 = ~n11291;
  assign n11272 = ~n11390;
  assign n11376 = n11391 & n11392;
  assign n11405 = ~n11442;
  assign n11453 = ~n11474;
  assign n11455 = n53 ^ n11485;
  assign n11488 = n11499 & n11500;
  assign n11413 = ~n11501;
  assign n11513 = n11528 & n11529;
  assign n11514 = n11383 & n11432;
  assign n11502 = n11540 & n11541;
  assign n11515 = ~n11383;
  assign n11518 = n11549 ^ n9067;
  assign n11550 = ~n11549;
  assign n11130 = n11288 ^ n11289;
  assign n11210 = n11289 & n11288;
  assign n11335 = n11346 & n11347;
  assign n11251 = ~n11348;
  assign n11333 = ~n11359;
  assign n11317 = ~n11376;
  assign n11393 = n11404 & n11405;
  assign n11443 = n11452 & n11453;
  assign n11406 = n11453 & n11409;
  assign n11425 = n11454 ^ n11455;
  assign n11456 = ~n11455;
  assign n11459 = ~n11488;
  assign n11464 = n11502 ^ n11503;
  assign n11486 = ~n11513;
  assign n11434 = ~n11514;
  assign n11506 = n11515 & n11516;
  assign n7821 = n11517 ^ n11518;
  assign n11504 = ~n11502;
  assign n11542 = n11550 & n11551;
  assign n11111 = ~n11130;
  assign n11213 = ~n11210;
  assign n11290 = n11333 & n11334;
  assign n11292 = ~n11335;
  assign n11306 = n11272 & n11317;
  assign n11360 = ~n11393;
  assign n7352 = n11406 ^ n11407;
  assign n11411 = n11425 & n8429;
  assign n11408 = ~n11443;
  assign n11410 = ~n11425;
  assign n11378 = n11456 & n11457;
  assign n11426 = n11459 & n11413;
  assign n11444 = n11464 ^ n11465;
  assign n11427 = n11486 & n11487;
  assign n11460 = n7821 & n10298;
  assign n11475 = n7821 & n11490;
  assign n11489 = n11504 & n11505;
  assign n11385 = ~n11506;
  assign n7827 = ~n7821;
  assign n11519 = ~n11542;
  assign n11249 = n11290 ^ n11291;
  assign n11293 = ~n11290;
  assign n11307 = n11360 & n11361;
  assign n9735 = n7352 ^ n11362;
  assign n11363 = n7352 & n11377;
  assign n11336 = n7352 & n9639;
  assign n7367 = ~n7352;
  assign n11320 = n11408 & n11409;
  assign n11394 = n11410 & n8438;
  assign n11364 = ~n11411;
  assign n11379 = n11426 ^ n11427;
  assign n11381 = ~n11378;
  assign n11430 = n11444 & n51;
  assign n11428 = ~n11444;
  assign n11299 = n11460 ^ n9067;
  assign n11458 = ~n11427;
  assign n10351 = ~n11475;
  assign n11468 = n7827 & n11476;
  assign n11466 = ~n11489;
  assign n11477 = n11519 & n11520;
  assign n11211 = n259 ^ n11249;
  assign n11270 = n11292 & n11293;
  assign n11169 = n11306 ^ n11307;
  assign n11309 = n11336 ^ n8475;
  assign n11318 = ~n11307;
  assign n9737 = ~n11363;
  assign n11349 = n7367 & n11362;
  assign n11351 = n11378 ^ n11379;
  assign n11365 = ~n11320;
  assign n11322 = ~n11394;
  assign n11380 = ~n11379;
  assign n11414 = n11428 & n11429;
  assign n11327 = ~n11430;
  assign n11415 = n11299 & n11342;
  assign n11416 = ~n11299;
  assign n11445 = n11458 & n11459;
  assign n11431 = n11466 & n11467;
  assign n10332 = ~n11468;
  assign n11446 = n11477 ^ n11478;
  assign n11479 = ~n11477;
  assign n9591 = n11210 ^ n11211;
  assign n11212 = ~n11211;
  assign n11250 = ~n11270;
  assign n11182 = ~n11169;
  assign n11294 = n11309 & n11310;
  assign n11308 = n11317 & n11318;
  assign n11295 = ~n11309;
  assign n9713 = ~n11349;
  assign n11337 = n11351 & n8389;
  assign n11350 = n11364 & n11365;
  assign n11319 = n11322 & n11364;
  assign n11338 = ~n11351;
  assign n11278 = n11380 & n11381;
  assign n11367 = ~n11414;
  assign n11301 = ~n11415;
  assign n11395 = n11416 & n11417;
  assign n11382 = n11431 ^ n11432;
  assign n11412 = ~n11445;
  assign n11435 = n10351 & n10332;
  assign n7708 = n11446 ^ n9006;
  assign n11433 = ~n11431;
  assign n11469 = n11479 & n11480;
  assign n11043 = ~n9591;
  assign n11128 = n11212 & n11213;
  assign n11214 = n11250 & n11251;
  assign n11195 = ~n11294;
  assign n11273 = n11295 & n11296;
  assign n11271 = ~n11308;
  assign n7235 = n11319 ^ n11320;
  assign n11239 = ~n11337;
  assign n11323 = n11338 & n8376;
  assign n11321 = ~n11350;
  assign n11368 = n11367 & n11327;
  assign n11281 = n11382 ^ n11383;
  assign n11344 = ~n11395;
  assign n11324 = n11412 & n11413;
  assign n11396 = n7708 & n11419;
  assign n11418 = n11433 & n11434;
  assign n10349 = ~n11435;
  assign n7814 = ~n7708;
  assign n11447 = ~n11469;
  assign n11168 = n258 ^ n11214;
  assign n11216 = n11214 & n11226;
  assign n11215 = ~n11214;
  assign n11196 = n11271 & n11272;
  assign n11236 = ~n11273;
  assign n11252 = n7235 & n9644;
  assign n11274 = n7235 & n11297;
  assign n7247 = ~n7235;
  assign n11240 = n11321 & n11322;
  assign n11276 = ~n11323;
  assign n11339 = n11281 & n11352;
  assign n11325 = ~n11368;
  assign n11340 = ~n11281;
  assign n11366 = ~n11324;
  assign n11354 = n7814 & n10261;
  assign n10294 = ~n11396;
  assign n11386 = n7814 & n11397;
  assign n11384 = ~n11418;
  assign n11399 = n11447 & n11448;
  assign n11129 = n11168 ^ n11169;
  assign n11193 = n11215 & n258;
  assign n11181 = ~n11216;
  assign n11237 = n11195 & n11236;
  assign n11150 = n11252 ^ n8438;
  assign n11235 = ~n11196;
  assign n9702 = ~n11274;
  assign n11261 = n7247 & n9682;
  assign n11277 = n11276 & n11239;
  assign n11275 = ~n11240;
  assign n11279 = n11324 ^ n11325;
  assign n11283 = ~n11339;
  assign n11328 = n11340 & n50;
  assign n11221 = n11354 ^ n8999;
  assign n11353 = n11366 & n11367;
  assign n11341 = n11384 & n11385;
  assign n10314 = ~n11386;
  assign n7689 = n11398 ^ n11399;
  assign n11400 = ~n11399;
  assign n10941 = n11128 ^ n11129;
  assign n11006 = n11129 & n11128;
  assign n11170 = n11181 & n11182;
  assign n11140 = ~n11193;
  assign n11219 = n11150 & n11108;
  assign n11227 = n11235 & n11236;
  assign n11197 = ~n11237;
  assign n11217 = ~n11150;
  assign n9685 = ~n11261;
  assign n11262 = n11275 & n11276;
  assign n11241 = ~n11277;
  assign n11253 = n11278 ^ n11279;
  assign n11203 = n11279 & n11278;
  assign n11246 = ~n11328;
  assign n11311 = n11221 & n11329;
  assign n11298 = n11341 ^ n11342;
  assign n11312 = ~n11221;
  assign n11326 = ~n11353;
  assign n10311 = n10314 & n10294;
  assign n11343 = ~n11341;
  assign n11331 = n7689 & n10224;
  assign n11356 = n7689 & n11369;
  assign n7725 = ~n7689;
  assign n11387 = n11400 & n11401;
  assign n10959 = ~n10941;
  assign n11013 = ~n11006;
  assign n11139 = ~n11170;
  assign n11171 = n11196 ^ n11197;
  assign n11198 = n11217 & n11218;
  assign n11151 = ~n11219;
  assign n11194 = ~n11227;
  assign n7216 = n11240 ^ n11241;
  assign n11242 = n11253 & n8298;
  assign n11238 = ~n11262;
  assign n11243 = ~n11253;
  assign n11206 = n11298 ^ n11299;
  assign n11224 = ~n11311;
  assign n11304 = n11312 & n11257;
  assign n11280 = n11326 & n11327;
  assign n11302 = n11331 ^ n8935;
  assign n11330 = n11343 & n11344;
  assign n11345 = n7725 & n11355;
  assign n10274 = ~n11356;
  assign n11357 = ~n11387;
  assign n11058 = n11139 & n11140;
  assign n11155 = n11171 & n257;
  assign n11153 = ~n11171;
  assign n11149 = n11194 & n11195;
  assign n11110 = ~n11198;
  assign n11199 = n7216 & n11220;
  assign n7202 = ~n7216;
  assign n11162 = n11238 & n11239;
  assign n11158 = ~n11242;
  assign n11228 = n11243 & n8360;
  assign n11254 = n11206 & n11263;
  assign n11244 = n11280 ^ n11281;
  assign n11255 = ~n11206;
  assign n11286 = n11302 & n11303;
  assign n11259 = ~n11304;
  assign n11282 = ~n11280;
  assign n11284 = ~n11302;
  assign n11300 = ~n11330;
  assign n10251 = ~n11345;
  assign n11313 = n11357 & n11358;
  assign n11094 = ~n11058;
  assign n11107 = n11149 ^ n11150;
  assign n11142 = n11153 & n11154;
  assign n11056 = ~n11155;
  assign n11152 = ~n11149;
  assign n9651 = ~n11199;
  assign n11183 = n7202 & n11200;
  assign n11156 = n7202 & n9565;
  assign n11201 = ~n11162;
  assign n11202 = ~n11228;
  assign n11204 = n50 ^ n11244;
  assign n11208 = ~n11254;
  assign n11247 = n11255 & n49;
  assign n11264 = n11282 & n11283;
  assign n11265 = n11284 & n11285;
  assign n11137 = ~n11286;
  assign n11256 = n11300 & n11301;
  assign n10271 = n10274 & n10251;
  assign n7673 = n11313 ^ n11314;
  assign n11315 = ~n11313;
  assign n11009 = n11107 ^ n11108;
  assign n11095 = ~n11142;
  assign n11141 = n11151 & n11152;
  assign n11131 = n11156 ^ n8376;
  assign n9668 = ~n11183;
  assign n11184 = n11201 & n11202;
  assign n11117 = n11203 ^ n11204;
  assign n11161 = n11202 & n11158;
  assign n11120 = n11204 & n11203;
  assign n11165 = ~n11247;
  assign n11222 = n11256 ^ n11257;
  assign n11245 = ~n11264;
  assign n11178 = ~n11265;
  assign n11258 = ~n11256;
  assign n11266 = n7673 & n11287;
  assign n7616 = ~n7673;
  assign n11305 = n11315 & n11316;
  assign n11070 = n11009 & n11085;
  assign n11086 = n11094 & n11095;
  assign n11071 = ~n11009;
  assign n11096 = n11095 & n11056;
  assign n11113 = n11131 & n11132;
  assign n11109 = ~n11141;
  assign n11114 = ~n11131;
  assign n9665 = n9668 & n9651;
  assign n7099 = n11161 ^ n11162;
  assign n11160 = n11117 & n8337;
  assign n11157 = ~n11184;
  assign n11159 = ~n11117;
  assign n11185 = n11221 ^ n11222;
  assign n11205 = n11245 & n11246;
  assign n11229 = n11178 & n11137;
  assign n11248 = n11258 & n11259;
  assign n11230 = n7616 & n10177;
  assign n10208 = ~n11266;
  assign n11260 = n7616 & n11267;
  assign n11268 = ~n11305;
  assign n11011 = ~n11070;
  assign n11057 = n11071 & n256;
  assign n11055 = ~n11086;
  assign n11059 = ~n11096;
  assign n11015 = n11109 & n11110;
  assign n11025 = ~n11113;
  assign n11098 = n11114 & n11115;
  assign n11112 = n7099 & n11130;
  assign n11087 = n7099 & n9523;
  assign n7120 = ~n7099;
  assign n11116 = n11157 & n11158;
  assign n11143 = n11159 & n8283;
  assign n11076 = ~n11160;
  assign n11174 = n11185 & n48;
  assign n11163 = n11205 ^ n11206;
  assign n11172 = ~n11185;
  assign n11207 = ~n11205;
  assign n11176 = ~n11229;
  assign n11048 = n11230 ^ n8898;
  assign n11223 = ~n11248;
  assign n10232 = ~n11260;
  assign n11231 = n11268 & n11269;
  assign n11008 = n11055 & n11056;
  assign n10971 = ~n11057;
  assign n11007 = n11058 ^ n11059;
  assign n11062 = n11087 ^ n8360;
  assign n11072 = ~n11015;
  assign n11073 = ~n11098;
  assign n11097 = n7120 & n11111;
  assign n9637 = ~n11112;
  assign n11074 = n11116 ^ n11117;
  assign n11118 = ~n11116;
  assign n11119 = ~n11143;
  assign n11121 = n49 ^ n11163;
  assign n11166 = n11172 & n11173;
  assign n11082 = ~n11174;
  assign n11186 = n11207 & n11208;
  assign n11187 = n11048 & n11209;
  assign n11175 = n11223 & n11224;
  assign n11188 = ~n11048;
  assign n10229 = n10232 & n10208;
  assign n7640 = n11231 ^ n11232;
  assign n11233 = ~n11231;
  assign n10869 = n11006 ^ n11007;
  assign n10969 = n11008 ^ n11009;
  assign n11010 = ~n11008;
  assign n11012 = ~n11007;
  assign n11046 = n11062 & n11063;
  assign n11060 = n11072 & n11073;
  assign n7067 = n11074 ^ n8337;
  assign n11064 = n11025 & n11073;
  assign n11044 = ~n11062;
  assign n9617 = ~n11097;
  assign n11099 = n11118 & n11119;
  assign n11028 = n11120 ^ n11121;
  assign n11031 = n11121 & n11120;
  assign n11123 = ~n11166;
  assign n11036 = n11175 ^ n11176;
  assign n11164 = ~n11186;
  assign n11050 = ~n11187;
  assign n11179 = n11188 & n11089;
  assign n11177 = ~n11175;
  assign n11189 = n7640 & n10169;
  assign n7628 = ~n7640;
  assign n11225 = n11233 & n11234;
  assign n10926 = n256 ^ n10969;
  assign n10853 = ~n10869;
  assign n10996 = n11010 & n11011;
  assign n10925 = n11012 & n11013;
  assign n11023 = n7067 & n11043;
  assign n10997 = n7067 & n9534;
  assign n11026 = n11044 & n11045;
  assign n10943 = ~n11046;
  assign n11024 = ~n11060;
  assign n7076 = ~n7067;
  assign n11016 = ~n11064;
  assign n11061 = n9637 & n9617;
  assign n11078 = n11028 & n8304;
  assign n11075 = ~n11099;
  assign n11077 = ~n11028;
  assign n11034 = ~n11031;
  assign n11124 = n11123 & n11082;
  assign n11135 = n11036 & n63;
  assign n11079 = n11164 & n11165;
  assign n11133 = ~n11036;
  assign n11167 = n11177 & n11178;
  assign n11091 = ~n11179;
  assign n11144 = n7628 & n10127;
  assign n10171 = ~n11189;
  assign n11180 = n7628 & n11190;
  assign n11191 = ~n11225;
  assign n9490 = n10925 ^ n10926;
  assign n10970 = ~n10996;
  assign n10939 = ~n10925;
  assign n10972 = n10997 ^ n8283;
  assign n10986 = n11015 ^ n11016;
  assign n11014 = n7076 & n9591;
  assign n9607 = ~n11023;
  assign n10945 = n11024 & n11025;
  assign n10985 = ~n11026;
  assign n9635 = ~n11061;
  assign n11027 = n11075 & n11076;
  assign n11065 = n11077 & n8294;
  assign n10990 = ~n11078;
  assign n11080 = ~n11124;
  assign n11125 = n11133 & n11134;
  assign n10993 = ~n11135;
  assign n11122 = ~n11079;
  assign n10965 = n11144 ^ n8854;
  assign n11136 = ~n11167;
  assign n10188 = ~n11180;
  assign n11146 = n11191 & n11192;
  assign n10767 = ~n9490;
  assign n10823 = n10926 & n10939;
  assign n10864 = n10970 & n10971;
  assign n10962 = n10972 & n10973;
  assign n10977 = n10986 & n271;
  assign n10960 = ~n10972;
  assign n10975 = ~n10986;
  assign n10988 = n10943 & n10985;
  assign n9594 = ~n11014;
  assign n10984 = ~n10945;
  assign n10987 = n11027 ^ n11028;
  assign n11029 = ~n11027;
  assign n11030 = ~n11065;
  assign n11032 = n11079 ^ n11080;
  assign n11100 = n11122 & n11123;
  assign n11038 = ~n11125;
  assign n11101 = n10965 & n11126;
  assign n11088 = n11136 & n11137;
  assign n11102 = ~n10965;
  assign n7469 = n11145 ^ n11146;
  assign n11147 = ~n11146;
  assign n10927 = ~n10864;
  assign n10944 = n10960 & n10961;
  assign n10850 = ~n10962;
  assign n10963 = n10975 & n10976;
  assign n10880 = ~n10977;
  assign n10974 = n10984 & n10985;
  assign n7007 = n10987 ^ n8304;
  assign n10946 = ~n10988;
  assign n11017 = n11029 & n11030;
  assign n10899 = n11031 ^ n11032;
  assign n11033 = ~n11032;
  assign n11047 = n11088 ^ n11089;
  assign n11081 = ~n11100;
  assign n10967 = ~n11101;
  assign n11092 = n11102 & n11002;
  assign n11090 = ~n11088;
  assign n11084 = n7469 & n10093;
  assign n11104 = n7469 & n11127;
  assign n7530 = ~n7469;
  assign n11138 = n11147 & n11148;
  assign n10893 = ~n10944;
  assign n10910 = n10945 ^ n10946;
  assign n10940 = n7007 & n10959;
  assign n10928 = ~n10963;
  assign n10911 = n7007 & n9520;
  assign n10942 = ~n10974;
  assign n7017 = ~n7007;
  assign n10989 = ~n11017;
  assign n10914 = ~n10899;
  assign n10950 = n11033 & n11034;
  assign n10953 = n11047 ^ n11048;
  assign n11035 = n11081 & n11082;
  assign n11051 = n11084 ^ n8800;
  assign n11083 = n11090 & n11091;
  assign n11004 = ~n11092;
  assign n11093 = n7530 & n11103;
  assign n10154 = ~n11104;
  assign n11105 = ~n11138;
  assign n10897 = n10850 & n10893;
  assign n10898 = n10910 & n270;
  assign n10881 = n10911 ^ n8294;
  assign n10909 = n10927 & n10928;
  assign n10912 = n10928 & n10880;
  assign n10895 = ~n10910;
  assign n9573 = ~n10940;
  assign n10929 = n7017 & n10941;
  assign n10847 = n10942 & n10943;
  assign n10947 = n10989 & n10990;
  assign n11000 = n10953 & n62;
  assign n10991 = n11035 ^ n11036;
  assign n10998 = ~n10953;
  assign n11039 = n11051 & n11052;
  assign n11037 = ~n11035;
  assign n11040 = ~n11051;
  assign n11049 = ~n11083;
  assign n10131 = ~n11093;
  assign n11066 = n11105 & n11106;
  assign n10868 = n10881 & n10882;
  assign n10884 = n10895 & n10896;
  assign n10848 = ~n10897;
  assign n10795 = ~n10898;
  assign n10866 = ~n10881;
  assign n10879 = ~n10909;
  assign n10865 = ~n10912;
  assign n9554 = ~n10929;
  assign n10894 = ~n10847;
  assign n10900 = n10947 ^ n8229;
  assign n10949 = n10947 & n8229;
  assign n10948 = ~n10947;
  assign n10951 = n63 ^ n10991;
  assign n10994 = n10998 & n10999;
  assign n10906 = ~n11000;
  assign n11018 = n11037 & n11038;
  assign n10876 = ~n11039;
  assign n11019 = n11040 & n11041;
  assign n11001 = n11049 & n11050;
  assign n11053 = n10154 & n10131;
  assign n7357 = n11066 ^ n11067;
  assign n11068 = ~n11066;
  assign n10826 = n10847 ^ n10848;
  assign n10824 = n10864 ^ n10865;
  assign n10851 = n10866 & n10867;
  assign n10772 = ~n10868;
  assign n10796 = n10879 & n10880;
  assign n10838 = ~n10884;
  assign n9570 = n9573 & n9554;
  assign n10883 = n10893 & n10894;
  assign n6951 = n10899 ^ n10900;
  assign n10930 = n10948 & n8211;
  assign n10913 = ~n10949;
  assign n10915 = n10950 ^ n10951;
  assign n10854 = n10951 & n10950;
  assign n10955 = ~n10994;
  assign n10964 = n11001 ^ n11002;
  assign n10992 = ~n11018;
  assign n10922 = ~n11019;
  assign n11003 = ~n11001;
  assign n11020 = n7357 & n11042;
  assign n10152 = ~n11053;
  assign n7492 = ~n7357;
  assign n11054 = n11068 & n11069;
  assign n10684 = n10823 ^ n10824;
  assign n10807 = n10826 & n269;
  assign n10755 = n10824 & n10823;
  assign n10805 = ~n10826;
  assign n10839 = n10838 & n10795;
  assign n10809 = ~n10851;
  assign n10837 = ~n10796;
  assign n10852 = n6951 & n10869;
  assign n10827 = n6951 & n9481;
  assign n10849 = ~n10883;
  assign n6995 = ~n6951;
  assign n10901 = n10913 & n10914;
  assign n10903 = n10915 & n8198;
  assign n10871 = ~n10930;
  assign n10902 = ~n10915;
  assign n10857 = ~n10854;
  assign n10931 = n10964 ^ n10965;
  assign n10952 = n10992 & n10993;
  assign n10978 = n10922 & n10876;
  assign n10995 = n11003 & n11004;
  assign n10979 = n7492 & n10033;
  assign n10088 = ~n11020;
  assign n11005 = n7492 & n10107;
  assign n11021 = ~n11054;
  assign n10676 = ~n10684;
  assign n10798 = n10805 & n10806;
  assign n10708 = ~n10807;
  assign n10760 = ~n10755;
  assign n10810 = n10772 & n10809;
  assign n10683 = n10827 ^ n8229;
  assign n10825 = n10837 & n10838;
  assign n10797 = ~n10839;
  assign n10769 = n10849 & n10850;
  assign n9532 = ~n10852;
  assign n10840 = n6995 & n10853;
  assign n10870 = ~n10901;
  assign n10885 = n10902 & n8209;
  assign n10829 = ~n10903;
  assign n10918 = n10931 & n61;
  assign n10904 = n10952 ^ n10953;
  assign n10916 = ~n10931;
  assign n10954 = ~n10952;
  assign n10920 = ~n10978;
  assign n10956 = n10979 ^ n8818;
  assign n10966 = ~n10995;
  assign n10109 = ~n11005;
  assign n10980 = n11021 & n11022;
  assign n10756 = n10796 ^ n10797;
  assign n10758 = ~n10798;
  assign n10770 = ~n10810;
  assign n10794 = ~n10825;
  assign n10808 = ~n10769;
  assign n9509 = ~n10840;
  assign n10812 = n10870 & n10871;
  assign n10786 = ~n10885;
  assign n10855 = n62 ^ n10904;
  assign n10907 = n10916 & n10917;
  assign n10819 = ~n10918;
  assign n10932 = n10954 & n10955;
  assign n10935 = n10956 & n10957;
  assign n10919 = n10966 & n10967;
  assign n10933 = ~n10956;
  assign n7289 = n10980 ^ n10981;
  assign n10982 = ~n10980;
  assign n10601 = n10755 ^ n10756;
  assign n10720 = n10758 & n10708;
  assign n10646 = n10769 ^ n10770;
  assign n10759 = ~n10756;
  assign n10721 = n10794 & n10795;
  assign n10799 = n10808 & n10809;
  assign n9529 = n9532 & n9509;
  assign n10828 = ~n10812;
  assign n10811 = n10786 & n10829;
  assign n10830 = n10854 ^ n10855;
  assign n10856 = ~n10855;
  assign n10859 = ~n10907;
  assign n10886 = n10919 ^ n10920;
  assign n10905 = ~n10932;
  assign n10923 = n10933 & n10934;
  assign n10791 = ~n10935;
  assign n10921 = ~n10919;
  assign n10936 = n7289 & n10958;
  assign n7421 = ~n7289;
  assign n10968 = n10982 & n10983;
  assign n10681 = n10720 ^ n10721;
  assign n10616 = ~n10601;
  assign n10724 = n10646 & n268;
  assign n10680 = n10759 & n10760;
  assign n10722 = ~n10646;
  assign n10757 = ~n10721;
  assign n10771 = ~n10799;
  assign n6925 = n10811 ^ n10812;
  assign n10813 = n10828 & n10829;
  assign n10815 = n10830 & n8189;
  assign n10814 = ~n10830;
  assign n10773 = n10856 & n10857;
  assign n10860 = n10859 & n10819;
  assign n10874 = n10886 & n60;
  assign n10816 = n10905 & n10906;
  assign n10872 = ~n10886;
  assign n10908 = n10921 & n10922;
  assign n10834 = ~n10923;
  assign n10887 = n7421 & n9923;
  assign n10048 = ~n10936;
  assign n10924 = n7421 & n10067;
  assign n10937 = ~n10968;
  assign n9368 = n10680 ^ n10681;
  assign n10611 = n10681 & n10680;
  assign n10709 = n10722 & n10723;
  assign n10648 = ~n10724;
  assign n10744 = n10757 & n10758;
  assign n10725 = n10771 & n10772;
  assign n10768 = n6925 & n9490;
  assign n10745 = n6925 & n9417;
  assign n6968 = ~n6925;
  assign n10785 = ~n10813;
  assign n10800 = n10814 & n8176;
  assign n10700 = ~n10815;
  assign n10776 = ~n10773;
  assign n10817 = ~n10860;
  assign n10861 = n10872 & n10873;
  assign n10738 = ~n10874;
  assign n10858 = ~n10816;
  assign n10877 = n10834 & n10791;
  assign n10862 = n10887 ^ n8718;
  assign n10875 = ~n10908;
  assign n10069 = ~n10924;
  assign n10888 = n10937 & n10938;
  assign n10574 = ~n9368;
  assign n10674 = ~n10709;
  assign n10682 = n10725 ^ n10726;
  assign n10707 = ~n10744;
  assign n10729 = n10725 & n10726;
  assign n10711 = n10745 ^ n8198;
  assign n10727 = ~n10725;
  assign n10761 = n6968 & n10767;
  assign n9492 = ~n10768;
  assign n10713 = n10785 & n10786;
  assign n10747 = ~n10800;
  assign n10774 = n10816 ^ n10817;
  assign n10841 = n10858 & n10859;
  assign n10780 = ~n10861;
  assign n10844 = n10862 & n10863;
  assign n10831 = n10875 & n10876;
  assign n10832 = ~n10877;
  assign n10842 = ~n10862;
  assign n10845 = n10888 ^ n10889;
  assign n10892 = n10888 & n10889;
  assign n10890 = ~n10888;
  assign n10584 = n10682 ^ n10683;
  assign n10672 = n10707 & n10708;
  assign n10698 = n10711 & n10712;
  assign n10710 = n10727 & n10728;
  assign n10695 = ~n10729;
  assign n10696 = ~n10711;
  assign n9469 = ~n10761;
  assign n10746 = ~n10713;
  assign n10762 = n10747 & n10700;
  assign n10666 = n10773 ^ n10774;
  assign n10775 = ~n10774;
  assign n10777 = n10780 & n10738;
  assign n10801 = n10831 ^ n10832;
  assign n10818 = ~n10841;
  assign n10835 = n10842 & n10843;
  assign n10706 = ~n10844;
  assign n7255 = n8709 ^ n10845;
  assign n10833 = ~n10831;
  assign n10878 = n10890 & n10891;
  assign n10804 = ~n10892;
  assign n10645 = n268 ^ n10672;
  assign n10673 = ~n10672;
  assign n10685 = n10695 & n10683;
  assign n10686 = n10696 & n10697;
  assign n10600 = ~n10698;
  assign n10663 = ~n10710;
  assign n10730 = n10746 & n10747;
  assign n10731 = n10666 & n8137;
  assign n10714 = ~n10762;
  assign n10732 = ~n10666;
  assign n10733 = n10775 & n10776;
  assign n10789 = n10801 & n59;
  assign n10778 = n10818 & n10819;
  assign n10787 = ~n10801;
  assign n10782 = n7255 & n9951;
  assign n10820 = n10833 & n10834;
  assign n10753 = ~n10835;
  assign n7307 = ~n7255;
  assign n10846 = n10804 & n8607;
  assign n10822 = ~n10878;
  assign n10612 = n10645 ^ n10646;
  assign n10661 = n10673 & n10674;
  assign n10662 = ~n10685;
  assign n10639 = ~n10686;
  assign n6922 = n10713 ^ n10714;
  assign n10699 = ~n10730;
  assign n10668 = ~n10731;
  assign n10715 = n10732 & n8146;
  assign n10736 = ~n10733;
  assign n10734 = n10777 ^ n10778;
  assign n10748 = n10782 ^ n8709;
  assign n10781 = n10787 & n10788;
  assign n10657 = ~n10789;
  assign n10779 = ~n10778;
  assign n10792 = n10753 & n10706;
  assign n10790 = ~n10820;
  assign n10821 = ~n10846;
  assign n10836 = n10822 & n8709;
  assign n9329 = n10611 ^ n10612;
  assign n10556 = n10612 & n10611;
  assign n10647 = ~n10661;
  assign n10628 = n10662 & n10663;
  assign n10652 = n10600 & n10639;
  assign n10675 = n6922 & n10684;
  assign n10665 = n10699 & n10700;
  assign n6915 = ~n6922;
  assign n10642 = ~n10715;
  assign n10701 = n10733 ^ n10734;
  assign n10740 = n10748 & n10749;
  assign n10735 = ~n10734;
  assign n10741 = ~n10748;
  assign n10763 = n10779 & n10780;
  assign n10692 = ~n10781;
  assign n10750 = n10790 & n10791;
  assign n10751 = ~n10792;
  assign n10802 = n10821 & n10822;
  assign n10803 = ~n10836;
  assign n10506 = ~n9329;
  assign n10613 = n10647 & n10648;
  assign n10638 = ~n10628;
  assign n10629 = ~n10652;
  assign n10640 = n10665 ^ n10666;
  assign n9430 = ~n10675;
  assign n10664 = n6915 & n10676;
  assign n10649 = n6915 & n9323;
  assign n10667 = ~n10665;
  assign n10687 = n10701 & n8095;
  assign n10688 = ~n10701;
  assign n10654 = n10735 & n10736;
  assign n10644 = ~n10740;
  assign n10717 = n10741 & n10742;
  assign n10739 = n10692 & n10657;
  assign n10716 = n10750 ^ n10751;
  assign n10737 = ~n10763;
  assign n10752 = ~n10750;
  assign n10783 = ~n10802;
  assign n10793 = n10803 & n10804;
  assign n10583 = n267 ^ n10613;
  assign n10615 = n10613 & n10627;
  assign n10598 = n10628 ^ n10629;
  assign n10614 = ~n10613;
  assign n10630 = n10638 & n10639;
  assign n6898 = n10640 ^ n8146;
  assign n10625 = n10649 ^ n8176;
  assign n9453 = ~n10664;
  assign n10653 = n10667 & n10668;
  assign n10578 = ~n10687;
  assign n10677 = n10688 & n8048;
  assign n10704 = n10716 & n58;
  assign n10670 = ~n10717;
  assign n10689 = n10737 & n10738;
  assign n10690 = ~n10739;
  assign n10702 = ~n10716;
  assign n10743 = n10752 & n10753;
  assign n10764 = n10783 & n10784;
  assign n10765 = ~n10793;
  assign n10557 = n10583 ^ n10584;
  assign n10590 = n10598 & n266;
  assign n10597 = n10614 & n267;
  assign n10587 = ~n10615;
  assign n10588 = ~n10598;
  assign n10602 = n6898 & n10616;
  assign n10617 = n10625 & n10626;
  assign n10599 = ~n10630;
  assign n6888 = ~n6898;
  assign n10618 = ~n10625;
  assign n9450 = n9453 & n9430;
  assign n10641 = ~n10653;
  assign n10607 = ~n10677;
  assign n10655 = n10689 ^ n10690;
  assign n10679 = n10670 & n10644;
  assign n10693 = n10702 & n10703;
  assign n10596 = ~n10704;
  assign n10691 = ~n10689;
  assign n10705 = ~n10743;
  assign n10719 = ~n10764;
  assign n10754 = n10765 & n10766;
  assign n10485 = n10556 ^ n10557;
  assign n10508 = n10557 & n10556;
  assign n10585 = n10587 & n10584;
  assign n10586 = n10588 & n10589;
  assign n10511 = ~n10590;
  assign n10564 = ~n10597;
  assign n10548 = n10599 & n10600;
  assign n10575 = n6888 & n9283;
  assign n10591 = n6888 & n10601;
  assign n9385 = ~n10602;
  assign n10544 = ~n10617;
  assign n10603 = n10618 & n10619;
  assign n10605 = n10641 & n10642;
  assign n10604 = n10607 & n10578;
  assign n10526 = n10654 ^ n10655;
  assign n10593 = n10655 & n10654;
  assign n10651 = ~n10679;
  assign n10678 = n10691 & n10692;
  assign n10636 = ~n10693;
  assign n10650 = n10705 & n10706;
  assign n10718 = ~n10754;
  assign n9267 = ~n10485;
  assign n10558 = n10575 ^ n8137;
  assign n10563 = ~n10585;
  assign n10536 = ~n10586;
  assign n10571 = ~n10548;
  assign n9406 = ~n10591;
  assign n10572 = ~n10603;
  assign n6789 = n10604 ^ n10605;
  assign n10606 = ~n10605;
  assign n10631 = n10526 & n8061;
  assign n10632 = ~n10526;
  assign n10637 = n10650 ^ n10651;
  assign n10658 = n10636 & n10596;
  assign n10656 = ~n10678;
  assign n10669 = ~n10650;
  assign n7209 = n10718 & n10719;
  assign n10547 = n10558 & n10559;
  assign n10534 = n10563 & n10564;
  assign n10533 = n10536 & n10511;
  assign n10545 = ~n10558;
  assign n10565 = n10571 & n10572;
  assign n9403 = n9406 & n9385;
  assign n10573 = n6789 & n9368;
  assign n10560 = n6789 & n9295;
  assign n10576 = n10572 & n10544;
  assign n6861 = ~n6789;
  assign n10592 = n10606 & n10607;
  assign n10528 = ~n10631;
  assign n10620 = n10632 & n8054;
  assign n10624 = n10637 & n57;
  assign n10622 = ~n10637;
  assign n10633 = n10656 & n10657;
  assign n10634 = ~n10658;
  assign n10659 = n10669 & n10670;
  assign n10660 = n7209 & n10694;
  assign n8673 = ~n7209;
  assign n10509 = n10533 ^ n10534;
  assign n10537 = n10545 & n10546;
  assign n10499 = ~n10547;
  assign n10535 = ~n10534;
  assign n10538 = n10560 ^ n8048;
  assign n10543 = ~n10565;
  assign n9370 = ~n10573;
  assign n10566 = n6861 & n10574;
  assign n10549 = ~n10576;
  assign n10577 = ~n10592;
  assign n10552 = ~n10620;
  assign n10608 = n10622 & n10623;
  assign n10542 = ~n10624;
  assign n10594 = n10633 ^ n10634;
  assign n10635 = ~n10633;
  assign n10643 = ~n10659;
  assign n10581 = n10660 ^ n8586;
  assign n9969 = n10671 ^ n8673;
  assign n10432 = n10508 ^ n10509;
  assign n10446 = n10509 & n10508;
  assign n10529 = n10535 & n10536;
  assign n10520 = ~n10537;
  assign n10532 = n10538 & n10539;
  assign n10491 = n10543 & n10544;
  assign n10465 = n10548 ^ n10549;
  assign n10530 = ~n10538;
  assign n9349 = ~n10566;
  assign n10550 = n10577 & n10578;
  assign n10579 = n10593 ^ n10594;
  assign n10517 = n10594 & n10593;
  assign n10570 = ~n10608;
  assign n10621 = n10635 & n10636;
  assign n10609 = n10643 & n10644;
  assign n9965 = ~n9969;
  assign n9229 = ~n10432;
  assign n10514 = n10520 & n10499;
  assign n10510 = ~n10529;
  assign n10523 = n10465 & n265;
  assign n10524 = n10530 & n10531;
  assign n10455 = ~n10532;
  assign n10519 = ~n10491;
  assign n10521 = ~n10465;
  assign n10525 = n10550 ^ n8054;
  assign n10551 = ~n10550;
  assign n10568 = n10579 & n7996;
  assign n10567 = ~n10579;
  assign n10582 = n10570 & n10542;
  assign n10580 = n10609 ^ n10610;
  assign n10595 = ~n10621;
  assign n10487 = n10510 & n10511;
  assign n10492 = ~n10514;
  assign n10512 = n10519 & n10520;
  assign n10513 = n10521 & n10522;
  assign n10467 = ~n10523;
  assign n10481 = ~n10524;
  assign n6707 = n10525 ^ n10526;
  assign n10540 = n10551 & n10552;
  assign n10561 = n10567 & n7965;
  assign n10484 = ~n10568;
  assign n10553 = n10580 ^ n10581;
  assign n10555 = ~n10582;
  assign n10554 = n10595 & n10596;
  assign n10464 = n265 ^ n10487;
  assign n10477 = n10491 ^ n10492;
  assign n10488 = ~n10487;
  assign n10497 = n6707 & n10506;
  assign n10478 = n10481 & n10455;
  assign n10498 = ~n10512;
  assign n10489 = ~n10513;
  assign n6809 = ~n6707;
  assign n10527 = ~n10540;
  assign n10516 = n56 ^ n10553;
  assign n10518 = n10554 ^ n10555;
  assign n10503 = ~n10561;
  assign n10569 = ~n10554;
  assign n10447 = n10464 ^ n10465;
  assign n10471 = n10477 & n264;
  assign n10469 = ~n10477;
  assign n10486 = n10488 & n10489;
  assign n9313 = ~n10497;
  assign n10490 = n6809 & n9329;
  assign n10479 = n10498 & n10499;
  assign n10482 = n6809 & n9246;
  assign n10507 = n10517 ^ n10518;
  assign n10501 = n10527 & n10528;
  assign n10494 = n10518 & n10517;
  assign n10500 = n10503 & n10484;
  assign n10562 = n10569 & n10570;
  assign n10381 = n10446 ^ n10447;
  assign n10409 = n10447 & n10446;
  assign n10460 = n10469 & n10470;
  assign n10429 = ~n10471;
  assign n10391 = n10478 ^ n10479;
  assign n10436 = n10482 ^ n8061;
  assign n10466 = ~n10486;
  assign n9331 = ~n10490;
  assign n10480 = ~n10479;
  assign n6731 = n10500 ^ n10501;
  assign n10504 = n10507 & n7986;
  assign n10502 = ~n10501;
  assign n10505 = ~n10507;
  assign n10541 = ~n10562;
  assign n9208 = ~n10381;
  assign n10412 = ~n10409;
  assign n10449 = ~n10460;
  assign n10457 = n10436 & n10461;
  assign n10431 = n10466 & n10467;
  assign n10396 = ~n10391;
  assign n10456 = ~n10436;
  assign n10472 = n10480 & n10481;
  assign n10476 = n6731 & n10485;
  assign n10462 = n6731 & n9212;
  assign n6741 = ~n6731;
  assign n10493 = n10502 & n10503;
  assign n10441 = ~n10504;
  assign n10496 = n10505 & n7976;
  assign n10515 = n10541 & n10542;
  assign n10430 = n10449 & n10429;
  assign n10450 = n10456 & n10420;
  assign n10438 = ~n10457;
  assign n10448 = ~n10431;
  assign n10383 = n10462 ^ n7965;
  assign n10454 = ~n10472;
  assign n10468 = n6741 & n9267;
  assign n9293 = ~n10476;
  assign n10483 = ~n10493;
  assign n10459 = ~n10496;
  assign n10495 = n10515 ^ n10516;
  assign n10410 = n10430 ^ n10431;
  assign n10442 = n10448 & n10449;
  assign n10422 = ~n10450;
  assign n10445 = n10383 & n10401;
  assign n10435 = n10454 & n10455;
  assign n10443 = ~n10383;
  assign n9270 = ~n10468;
  assign n10451 = n10483 & n10484;
  assign n10475 = n10459 & n10441;
  assign n10424 = n10494 ^ n10495;
  assign n9170 = n10409 ^ n10410;
  assign n10411 = ~n10410;
  assign n10419 = n10435 ^ n10436;
  assign n10428 = ~n10442;
  assign n10439 = n10443 & n10444;
  assign n10385 = ~n10445;
  assign n10437 = ~n10435;
  assign n10458 = ~n10451;
  assign n10452 = ~n10475;
  assign n10474 = n10424 & n7923;
  assign n10473 = ~n10424;
  assign n10345 = ~n9170;
  assign n10373 = n10411 & n10412;
  assign n10407 = n10419 ^ n10420;
  assign n10413 = n10428 & n10429;
  assign n10434 = n10437 & n10438;
  assign n10403 = ~n10439;
  assign n6713 = n10451 ^ n10452;
  assign n10453 = n10458 & n10459;
  assign n10463 = n10473 & n7909;
  assign n10406 = ~n10474;
  assign n10399 = n10407 & n278;
  assign n10390 = n279 ^ n10413;
  assign n10397 = ~n10407;
  assign n10415 = n10413 & n10418;
  assign n10414 = ~n10413;
  assign n10421 = ~n10434;
  assign n10433 = n6713 & n9229;
  assign n6700 = ~n6713;
  assign n10440 = ~n10453;
  assign n10426 = ~n10463;
  assign n10374 = n10390 ^ n10391;
  assign n10393 = n10397 & n10398;
  assign n10342 = ~n10399;
  assign n10408 = n10414 & n279;
  assign n10395 = ~n10415;
  assign n10400 = n10421 & n10422;
  assign n10427 = n6700 & n10432;
  assign n9231 = ~n10433;
  assign n10416 = n6700 & n9118;
  assign n10423 = n10440 & n10441;
  assign n10333 = n10373 ^ n10374;
  assign n10337 = n10374 & n10373;
  assign n10360 = ~n10393;
  assign n10392 = n10395 & n10396;
  assign n10382 = n10400 ^ n10401;
  assign n10379 = ~n10408;
  assign n10402 = ~n10400;
  assign n10343 = n10416 ^ n7986;
  assign n10404 = n10423 ^ n10424;
  assign n9252 = ~n10427;
  assign n10425 = ~n10423;
  assign n10322 = ~n10333;
  assign n10375 = n10360 & n10342;
  assign n10325 = n10382 ^ n10383;
  assign n10378 = ~n10392;
  assign n10394 = n10402 & n10403;
  assign n6641 = n10404 ^ n7909;
  assign n10353 = ~n10343;
  assign n10417 = n10425 & n10426;
  assign n10361 = n10325 & n10372;
  assign n10355 = ~n10375;
  assign n10362 = ~n10325;
  assign n10354 = n10378 & n10379;
  assign n10380 = n6641 & n9208;
  assign n10384 = ~n10394;
  assign n6629 = ~n6641;
  assign n10405 = ~n10417;
  assign n10338 = n10354 ^ n10355;
  assign n10327 = ~n10361;
  assign n10357 = n10362 & n277;
  assign n10359 = ~n10354;
  assign n9189 = ~n10380;
  assign n10376 = n6629 & n10381;
  assign n10363 = n10384 & n10385;
  assign n10368 = n6629 & n9135;
  assign n10386 = n10405 & n10406;
  assign n9059 = n10337 ^ n10338;
  assign n10282 = n10338 & n10337;
  assign n10305 = ~n10357;
  assign n10356 = n10359 & n10360;
  assign n10344 = n10363 ^ n10364;
  assign n10300 = n10368 ^ n7909;
  assign n10367 = n10363 & n10364;
  assign n9210 = ~n10376;
  assign n10365 = ~n10363;
  assign n10369 = n10386 ^ n10387;
  assign n10388 = ~n10386;
  assign n10295 = ~n9059;
  assign n10265 = n10343 ^ n10344;
  assign n10341 = ~n10356;
  assign n10358 = n10365 & n10366;
  assign n10352 = ~n10367;
  assign n6568 = n10369 ^ n7808;
  assign n10377 = n10388 & n10389;
  assign n10328 = n10265 & n10334;
  assign n10329 = ~n10265;
  assign n10324 = n10341 & n10342;
  assign n10346 = n6568 & n9170;
  assign n10347 = n10352 & n10353;
  assign n10336 = ~n10358;
  assign n6553 = ~n6568;
  assign n10370 = ~n10377;
  assign n10303 = n10324 ^ n10325;
  assign n10286 = ~n10328;
  assign n10319 = n10329 & n276;
  assign n10326 = ~n10324;
  assign n10339 = n6553 & n10345;
  assign n9146 = ~n10346;
  assign n10335 = ~n10347;
  assign n10330 = n6553 & n9094;
  assign n10348 = n10370 & n10371;
  assign n10283 = n277 ^ n10303;
  assign n10267 = ~n10319;
  assign n10318 = n10326 & n10327;
  assign n10236 = n10330 ^ n7888;
  assign n10320 = n10335 & n10336;
  assign n9172 = ~n10339;
  assign n6356 = n10348 ^ n10349;
  assign n10350 = ~n10348;
  assign n10245 = n10282 ^ n10283;
  assign n10241 = n10283 & n10282;
  assign n10308 = n10236 & n10315;
  assign n10304 = ~n10318;
  assign n10316 = n10320 & n10321;
  assign n10309 = ~n10236;
  assign n10306 = ~n10320;
  assign n10323 = n6356 & n10333;
  assign n6476 = ~n6356;
  assign n10340 = n10350 & n10351;
  assign n10252 = ~n10245;
  assign n10244 = ~n10241;
  assign n10284 = n10304 & n10305;
  assign n10288 = n10306 ^ n10300;
  assign n10240 = ~n10308;
  assign n10301 = n10309 & n10258;
  assign n10307 = n10306 & n10289;
  assign n10299 = ~n10316;
  assign n10317 = n6476 & n10322;
  assign n9106 = ~n10323;
  assign n10310 = n6476 & n8994;
  assign n10331 = ~n10340;
  assign n10264 = n276 ^ n10284;
  assign n10275 = n10288 ^ n10289;
  assign n10285 = ~n10284;
  assign n10296 = n10299 & n10300;
  assign n10260 = ~n10301;
  assign n10280 = ~n10307;
  assign n10297 = n10310 ^ n7821;
  assign n9127 = ~n10317;
  assign n10312 = n10331 & n10332;
  assign n10242 = n10264 ^ n10265;
  assign n10270 = n10275 & n275;
  assign n10268 = ~n10275;
  assign n10277 = n10285 & n10286;
  assign n10279 = ~n10296;
  assign n10292 = n10297 & n10298;
  assign n10290 = ~n10297;
  assign n9124 = n9127 & n9106;
  assign n6419 = n10311 ^ n10312;
  assign n10313 = ~n10312;
  assign n10209 = n10241 ^ n10242;
  assign n10243 = ~n10242;
  assign n10256 = n10268 & n10269;
  assign n10228 = ~n10270;
  assign n10266 = ~n10277;
  assign n10257 = n10279 & n10280;
  assign n10281 = n10290 & n10291;
  assign n10202 = ~n10292;
  assign n10287 = n6419 & n10295;
  assign n10276 = n6419 & n9006;
  assign n6437 = ~n6419;
  assign n10302 = n10313 & n10314;
  assign n10204 = ~n10209;
  assign n10194 = n10243 & n10244;
  assign n10248 = ~n10256;
  assign n10235 = n10257 ^ n10258;
  assign n10218 = n10266 & n10267;
  assign n10259 = ~n10257;
  assign n10163 = n10276 ^ n7814;
  assign n10223 = ~n10281;
  assign n9083 = ~n10287;
  assign n10278 = n6437 & n9059;
  assign n10293 = ~n10302;
  assign n10205 = ~n10194;
  assign n10226 = n10235 ^ n10236;
  assign n10238 = n10248 & n10228;
  assign n10247 = ~n10218;
  assign n10253 = n10259 & n10260;
  assign n10254 = n10163 & n10261;
  assign n10262 = n10223 & n10202;
  assign n10255 = ~n10163;
  assign n9062 = ~n10278;
  assign n10272 = n10293 & n10294;
  assign n10217 = n10226 & n274;
  assign n10215 = ~n10226;
  assign n10219 = ~n10238;
  assign n10237 = n10247 & n10248;
  assign n10239 = ~n10253;
  assign n10166 = ~n10254;
  assign n10249 = n10255 & n10182;
  assign n10221 = ~n10262;
  assign n6204 = n10271 ^ n10272;
  assign n10273 = ~n10272;
  assign n10210 = n10215 & n10216;
  assign n10180 = ~n10217;
  assign n10195 = n10218 ^ n10219;
  assign n10227 = ~n10237;
  assign n10220 = n10239 & n10240;
  assign n10184 = ~n10249;
  assign n10246 = n6204 & n10252;
  assign n10233 = n6204 & n8983;
  assign n6361 = ~n6204;
  assign n10263 = n10273 & n10274;
  assign n8961 = n10194 ^ n10195;
  assign n10155 = n10195 & n10205;
  assign n10196 = ~n10210;
  assign n10136 = n10220 ^ n10221;
  assign n10172 = n10227 & n10228;
  assign n10222 = ~n10220;
  assign n10144 = n10233 ^ n7689;
  assign n10234 = n6361 & n10245;
  assign n9044 = ~n10246;
  assign n10250 = ~n10263;
  assign n10150 = ~n8961;
  assign n10158 = ~n10155;
  assign n10190 = n10196 & n10180;
  assign n10200 = n10136 & n273;
  assign n10198 = ~n10136;
  assign n10197 = ~n10172;
  assign n10211 = n10222 & n10223;
  assign n10213 = n10144 & n10224;
  assign n10212 = ~n10144;
  assign n9025 = ~n10234;
  assign n10230 = n10250 & n10251;
  assign n10173 = ~n10190;
  assign n10189 = n10196 & n10197;
  assign n10191 = n10198 & n10199;
  assign n10138 = ~n10200;
  assign n10201 = ~n10211;
  assign n10206 = n10212 & n10123;
  assign n10125 = ~n10213;
  assign n10214 = n9044 & n9025;
  assign n6252 = n10229 ^ n10230;
  assign n10231 = ~n10230;
  assign n10156 = n10172 ^ n10173;
  assign n10179 = ~n10189;
  assign n10162 = ~n10191;
  assign n10181 = n10201 & n10202;
  assign n10146 = ~n10206;
  assign n10203 = n6252 & n10209;
  assign n10192 = n6252 & n8945;
  assign n9042 = ~n10214;
  assign n6268 = ~n6252;
  assign n10225 = n10231 & n10232;
  assign n10129 = n10155 ^ n10156;
  assign n10157 = ~n10156;
  assign n10160 = n10179 & n10180;
  assign n10164 = n10181 ^ n10182;
  assign n10183 = ~n10181;
  assign n10100 = n10192 ^ n7673;
  assign n9004 = ~n10203;
  assign n10193 = n6268 & n10204;
  assign n10207 = ~n10225;
  assign n8922 = ~n10129;
  assign n10115 = n10157 & n10158;
  assign n10135 = n273 ^ n10160;
  assign n10148 = n10163 ^ n10164;
  assign n10161 = ~n10160;
  assign n10174 = n10183 & n10184;
  assign n10175 = n10100 & n10080;
  assign n10176 = ~n10100;
  assign n8980 = ~n10193;
  assign n10186 = n10207 & n10208;
  assign n10116 = n10135 ^ n10136;
  assign n10118 = ~n10115;
  assign n10141 = n10148 & n272;
  assign n10139 = ~n10148;
  assign n10159 = n10161 & n10162;
  assign n10165 = ~n10174;
  assign n10102 = ~n10175;
  assign n10167 = n10176 & n10177;
  assign n10178 = n9004 & n8980;
  assign n10168 = n10186 ^ n7640;
  assign n10187 = ~n10186;
  assign n10070 = n10115 ^ n10116;
  assign n10117 = ~n10116;
  assign n10132 = n10139 & n10140;
  assign n10095 = ~n10141;
  assign n10137 = ~n10159;
  assign n10143 = n10165 & n10166;
  assign n10082 = ~n10167;
  assign n6174 = n10168 ^ n10169;
  assign n9002 = ~n10178;
  assign n10185 = n10187 & n10188;
  assign n10063 = ~n10070;
  assign n10071 = n10117 & n10118;
  assign n10120 = ~n10132;
  assign n10089 = n10137 & n10138;
  assign n10122 = n10143 ^ n10144;
  assign n10149 = n6174 & n8961;
  assign n10145 = ~n10143;
  assign n10134 = n6174 & n8891;
  assign n6054 = ~n6174;
  assign n10170 = ~n10185;
  assign n10074 = ~n10071;
  assign n10111 = n10120 & n10095;
  assign n10052 = n10122 ^ n10123;
  assign n10121 = ~n10089;
  assign n10126 = n10134 ^ n7628;
  assign n10133 = n10145 & n10146;
  assign n8963 = ~n10149;
  assign n10142 = n6054 & n10150;
  assign n10151 = n10170 & n10171;
  assign n10098 = n10052 & n287;
  assign n10090 = ~n10111;
  assign n10096 = ~n10052;
  assign n10110 = n10120 & n10121;
  assign n10112 = n10126 & n10127;
  assign n10113 = ~n10126;
  assign n10124 = ~n10133;
  assign n8942 = ~n10142;
  assign n5972 = n10151 ^ n10152;
  assign n10153 = ~n10151;
  assign n10072 = n10089 ^ n10090;
  assign n10091 = n10096 & n10097;
  assign n10055 = ~n10098;
  assign n10094 = ~n10110;
  assign n10043 = ~n10112;
  assign n10104 = n10113 & n10114;
  assign n10099 = n10124 & n10125;
  assign n10128 = n5972 & n8922;
  assign n6133 = ~n5972;
  assign n10147 = n10153 & n10154;
  assign n8827 = n10071 ^ n10072;
  assign n10073 = ~n10072;
  assign n10077 = ~n10091;
  assign n10076 = n10094 & n10095;
  assign n10079 = n10099 ^ n10100;
  assign n10061 = ~n10104;
  assign n10101 = ~n10099;
  assign n8903 = ~n10128;
  assign n10119 = n6133 & n10129;
  assign n10105 = n6133 & n8843;
  assign n10130 = ~n10147;
  assign n10022 = ~n8827;
  assign n10034 = n10073 & n10074;
  assign n10051 = n287 ^ n10076;
  assign n10037 = n10079 ^ n10080;
  assign n10078 = ~n10076;
  assign n10058 = n10061 & n10043;
  assign n10092 = n10101 & n10102;
  assign n10003 = n10105 ^ n7469;
  assign n8924 = ~n10119;
  assign n10106 = n10130 & n10131;
  assign n10035 = n10051 ^ n10052;
  assign n10056 = n10037 & n10065;
  assign n10057 = ~n10037;
  assign n10075 = n10077 & n10078;
  assign n10081 = ~n10092;
  assign n10085 = n10003 & n10093;
  assign n10084 = ~n10003;
  assign n10086 = n10106 ^ n10107;
  assign n10108 = ~n10106;
  assign n9983 = n10034 ^ n10035;
  assign n9996 = n10035 & n10034;
  assign n10039 = ~n10056;
  assign n10049 = n10057 & n286;
  assign n10054 = ~n10075;
  assign n10059 = n10081 & n10082;
  assign n10083 = n10084 & n10017;
  assign n10005 = ~n10085;
  assign n6024 = n10086 ^ n7357;
  assign n10103 = n10108 & n10109;
  assign n9990 = ~n9983;
  assign n10014 = ~n10049;
  assign n10036 = n10054 & n10055;
  assign n9971 = n10058 ^ n10059;
  assign n10064 = n6024 & n10070;
  assign n10060 = ~n10059;
  assign n10019 = ~n10083;
  assign n6001 = ~n6024;
  assign n10087 = ~n10103;
  assign n10012 = n10036 ^ n10037;
  assign n10040 = n9971 & n10044;
  assign n10038 = ~n10036;
  assign n10041 = ~n9971;
  assign n10050 = n10060 & n10061;
  assign n10053 = n6001 & n10063;
  assign n8860 = ~n10064;
  assign n10045 = n6001 & n8714;
  assign n10066 = n10087 & n10088;
  assign n9997 = n286 ^ n10012;
  assign n10031 = n10038 & n10039;
  assign n10001 = ~n10040;
  assign n10032 = n10041 & n285;
  assign n9957 = n10045 ^ n7492;
  assign n10042 = ~n10050;
  assign n8881 = ~n10053;
  assign n10046 = n10066 ^ n10067;
  assign n10068 = ~n10066;
  assign n9926 = n9996 ^ n9997;
  assign n9998 = ~n9997;
  assign n10013 = ~n10031;
  assign n9974 = ~n10032;
  assign n10025 = n9957 & n10033;
  assign n10016 = n10042 & n10043;
  assign n10024 = ~n9957;
  assign n8878 = n8881 & n8860;
  assign n5847 = n10046 ^ n7421;
  assign n10062 = n10068 & n10069;
  assign n9952 = n9998 & n9996;
  assign n9999 = n10013 & n10014;
  assign n10002 = n10016 ^ n10017;
  assign n10020 = n10024 & n9979;
  assign n9960 = ~n10025;
  assign n10023 = n5847 & n8827;
  assign n10018 = ~n10016;
  assign n10011 = n5847 & n8725;
  assign n5905 = ~n5847;
  assign n10047 = ~n10062;
  assign n9970 = n285 ^ n9999;
  assign n9985 = n10002 ^ n10003;
  assign n10000 = ~n9999;
  assign n9939 = n10011 ^ n7289;
  assign n10010 = n10018 & n10019;
  assign n9981 = ~n10020;
  assign n10015 = n5905 & n10022;
  assign n8829 = ~n10023;
  assign n10026 = n10047 & n10048;
  assign n9953 = n9970 ^ n9971;
  assign n9977 = n9985 & n284;
  assign n9975 = ~n9985;
  assign n9991 = n10000 & n10001;
  assign n9992 = n9939 & n10006;
  assign n9993 = ~n9939;
  assign n10004 = ~n10010;
  assign n8806 = ~n10015;
  assign n10008 = n10026 ^ n10027;
  assign n10030 = n10026 & n10027;
  assign n10028 = ~n10026;
  assign n8885 = n9952 ^ n9953;
  assign n9954 = ~n9953;
  assign n9966 = n9975 & n9976;
  assign n9934 = ~n9977;
  assign n9973 = ~n9991;
  assign n9941 = ~n9992;
  assign n9986 = n9993 & n9923;
  assign n9978 = n10004 & n10005;
  assign n5738 = n10008 ^ n7307;
  assign n10021 = n10028 & n10029;
  assign n9989 = ~n10030;
  assign n6735 = n8885 ^ n7817;
  assign n8848 = n8885 ^ n9930;
  assign n9869 = n8885 & n7817;
  assign n9918 = n9954 & n9952;
  assign n9956 = ~n9966;
  assign n9932 = n9973 & n9974;
  assign n9958 = n9978 ^ n9979;
  assign n9925 = ~n9986;
  assign n9984 = n5738 & n9990;
  assign n9980 = ~n9978;
  assign n5831 = ~n5738;
  assign n10009 = n9989 & n7307;
  assign n9995 = ~n10021;
  assign n8847 = ~n6735;
  assign n9931 = n9956 & n9934;
  assign n9943 = n9957 ^ n9958;
  assign n9955 = ~n9932;
  assign n9967 = n9980 & n9981;
  assign n9972 = n5831 & n9983;
  assign n8753 = ~n9984;
  assign n9962 = n5831 & n8607;
  assign n10007 = n9995 & n7255;
  assign n9994 = ~n10009;
  assign n9898 = n8847 & n8831;
  assign n9919 = n9931 ^ n9932;
  assign n9937 = n9943 & n283;
  assign n9935 = ~n9943;
  assign n9949 = n9955 & n9956;
  assign n9950 = n9962 ^ n7255;
  assign n9959 = ~n9967;
  assign n8758 = ~n9972;
  assign n9987 = n9994 & n9995;
  assign n9988 = ~n10007;
  assign n9892 = n9898 ^ n9899;
  assign n9879 = n9898 ^ n9900;
  assign n9914 = n9918 ^ n9919;
  assign n9882 = n9919 & n9918;
  assign n9927 = n9935 & n9936;
  assign n9906 = ~n9937;
  assign n9933 = ~n9949;
  assign n9944 = n9950 & n9951;
  assign n9938 = n9959 & n9960;
  assign n9945 = ~n9950;
  assign n8777 = n8758 & n8753;
  assign n9968 = ~n9987;
  assign n9982 = n9988 & n9989;
  assign n9575 = n487 ^ n9879;
  assign n9803 = n9892 & n9893;
  assign n9761 = n9879 & n487;
  assign n9901 = n9914 & n7792;
  assign n9902 = ~n9914;
  assign n9885 = ~n9882;
  assign n9921 = ~n9927;
  assign n9904 = n9933 & n9934;
  assign n9922 = n9938 ^ n9939;
  assign n9891 = ~n9944;
  assign n9942 = n9945 & n9946;
  assign n9940 = ~n9938;
  assign n9963 = n9968 & n9969;
  assign n9964 = ~n9982;
  assign n9568 = ~n9575;
  assign n9881 = ~n9901;
  assign n9895 = n9902 & n7642;
  assign n9903 = n9921 & n9906;
  assign n9915 = n9922 ^ n9923;
  assign n9920 = ~n9904;
  assign n9928 = n9940 & n9941;
  assign n9913 = ~n9942;
  assign n9948 = ~n9963;
  assign n9961 = n9964 & n9965;
  assign n9880 = n9881 & n9869;
  assign n9875 = ~n9895;
  assign n9883 = n9903 ^ n9904;
  assign n9909 = n9915 & n282;
  assign n9907 = ~n9915;
  assign n9916 = n9920 & n9921;
  assign n9910 = n9913 & n9891;
  assign n9924 = ~n9928;
  assign n9947 = ~n9961;
  assign n9874 = ~n9880;
  assign n9868 = n9875 & n9881;
  assign n9847 = n9882 ^ n9883;
  assign n9884 = ~n9883;
  assign n9896 = n9907 & n9908;
  assign n9871 = ~n9909;
  assign n9905 = ~n9916;
  assign n9911 = n9924 & n9925;
  assign n5715 = n9947 & n9948;
  assign n6665 = n9868 ^ n9869;
  assign n9863 = n9874 & n9875;
  assign n9851 = n9884 & n9885;
  assign n9887 = ~n9896;
  assign n9866 = n9905 & n9906;
  assign n9858 = n9910 ^ n9911;
  assign n9912 = ~n9911;
  assign n8722 = n9926 ^ n5715;
  assign n9917 = n5715 & n9929;
  assign n7271 = ~n5715;
  assign n9848 = n9863 ^ n7634;
  assign n9865 = n9863 & n7623;
  assign n6702 = ~n6665;
  assign n9864 = ~n9863;
  assign n9854 = ~n9851;
  assign n9877 = n9887 & n9871;
  assign n9888 = n9858 & n9894;
  assign n9886 = ~n9866;
  assign n9889 = ~n9858;
  assign n9897 = n9912 & n9913;
  assign n9861 = n9917 ^ n7209;
  assign n8728 = ~n8722;
  assign n6636 = n9847 ^ n9848;
  assign n9842 = n6702 & n8712;
  assign n9856 = n9864 & n7634;
  assign n9850 = ~n9865;
  assign n9867 = ~n9877;
  assign n9876 = n9886 & n9887;
  assign n9860 = ~n9888;
  assign n9878 = n9889 & n281;
  assign n9890 = ~n9897;
  assign n9821 = n6636 & n8670;
  assign n6646 = ~n6636;
  assign n9835 = n9842 ^ n7792;
  assign n9849 = n9850 & n9847;
  assign n9839 = ~n9856;
  assign n9852 = n9866 ^ n9867;
  assign n9870 = ~n9876;
  assign n9846 = ~n9878;
  assign n9872 = n9890 & n9891;
  assign n9770 = n9821 ^ n7623;
  assign n9829 = n9835 & n9836;
  assign n9827 = ~n9835;
  assign n9838 = ~n9849;
  assign n9824 = n9851 ^ n9852;
  assign n9853 = ~n9852;
  assign n9857 = n9870 & n9871;
  assign n9862 = n9872 ^ n9873;
  assign n9812 = n9770 & n9786;
  assign n9810 = ~n9770;
  assign n9822 = n9827 & n9828;
  assign n9805 = ~n9829;
  assign n9823 = n9838 & n9839;
  assign n9841 = n9824 & n7553;
  assign n9840 = ~n9824;
  assign n9830 = n9853 & n9854;
  assign n9843 = n9857 ^ n9858;
  assign n9844 = n9861 ^ n9862;
  assign n9859 = ~n9857;
  assign n9808 = n9810 & n9811;
  assign n9778 = ~n9812;
  assign n9817 = ~n9822;
  assign n9813 = n9823 ^ n9824;
  assign n9825 = ~n9823;
  assign n9837 = n9840 & n7568;
  assign n9826 = ~n9841;
  assign n9831 = n281 ^ n9843;
  assign n9834 = n280 ^ n9844;
  assign n9855 = n9859 & n9860;
  assign n9789 = ~n9808;
  assign n6588 = n9813 ^ n7553;
  assign n9814 = n9817 & n9803;
  assign n9802 = n9805 & n9817;
  assign n9820 = n9825 & n9826;
  assign n9794 = n9830 ^ n9831;
  assign n9816 = ~n9837;
  assign n9832 = ~n9831;
  assign n9845 = ~n9855;
  assign n9788 = n6588 & n8613;
  assign n9795 = n9802 ^ n9803;
  assign n6601 = ~n6588;
  assign n9804 = ~n9814;
  assign n9815 = ~n9820;
  assign n9818 = n9832 & n9830;
  assign n9833 = n9845 & n9846;
  assign n9756 = n9788 ^ n7553;
  assign n9792 = n9795 & n486;
  assign n9790 = ~n9795;
  assign n9797 = n9804 & n9805;
  assign n9798 = n9815 & n9816;
  assign n9819 = n9833 ^ n9834;
  assign n9776 = n9756 & n9742;
  assign n9774 = ~n9756;
  assign n9783 = n9790 & n9791;
  assign n9764 = ~n9792;
  assign n9785 = ~n9797;
  assign n9784 = n9798 ^ n9794;
  assign n9801 = n9798 & n7463;
  assign n9799 = ~n9798;
  assign n9809 = n9818 ^ n9819;
  assign n9769 = n9774 & n9775;
  assign n9747 = ~n9776;
  assign n9779 = ~n9783;
  assign n6517 = n7477 ^ n9784;
  assign n9771 = n9785 ^ n9786;
  assign n9782 = n9789 & n9785;
  assign n9796 = n9799 & n7477;
  assign n9793 = ~n9801;
  assign n9807 = n9809 & n7427;
  assign n9806 = ~n9809;
  assign n9759 = ~n9769;
  assign n9745 = n9770 ^ n9771;
  assign n9773 = n9779 & n9761;
  assign n9760 = n9779 & n9764;
  assign n9762 = n6517 & n8517;
  assign n6407 = ~n6517;
  assign n9777 = ~n9782;
  assign n9787 = n9793 & n9794;
  assign n9781 = ~n9796;
  assign n9800 = n9806 & n7347;
  assign n9749 = ~n9807;
  assign n9754 = n9745 & n485;
  assign n9551 = n9760 ^ n9761;
  assign n9715 = n9762 ^ n7463;
  assign n9752 = ~n9745;
  assign n9763 = ~n9773;
  assign n9772 = n9777 & n9778;
  assign n9780 = ~n9787;
  assign n9768 = ~n9800;
  assign n9750 = n9752 & n9753;
  assign n9726 = ~n9754;
  assign n9557 = ~n9551;
  assign n9757 = n9763 & n9764;
  assign n9755 = ~n9772;
  assign n9766 = n9780 & n9781;
  assign n9765 = n9768 & n9749;
  assign n9743 = ~n9750;
  assign n9741 = n9755 ^ n9756;
  assign n9744 = ~n9757;
  assign n9751 = n9759 & n9755;
  assign n6413 = n9765 ^ n9766;
  assign n9767 = ~n9766;
  assign n9731 = n9741 ^ n9742;
  assign n9739 = n9743 & n9744;
  assign n9723 = n9744 ^ n9745;
  assign n9740 = n6413 & n8505;
  assign n9746 = ~n9751;
  assign n6424 = ~n6413;
  assign n9758 = n9767 & n9768;
  assign n8287 = n485 ^ n9723;
  assign n9722 = n9731 & n484;
  assign n9720 = ~n9731;
  assign n9725 = ~n9739;
  assign n9728 = n9740 ^ n7347;
  assign n9738 = n9746 & n9747;
  assign n9748 = ~n9758;
  assign n9514 = ~n8287;
  assign n9716 = n9720 & n9721;
  assign n9695 = ~n9722;
  assign n9693 = n9725 & n9726;
  assign n9717 = n9728 & n9729;
  assign n9718 = ~n9728;
  assign n9733 = n9738 & n9707;
  assign n9724 = ~n9738;
  assign n9734 = n9748 & n9749;
  assign n9708 = ~n9716;
  assign n9709 = ~n9693;
  assign n9672 = ~n9717;
  assign n9711 = n9718 & n9719;
  assign n9706 = n9724 ^ n9715;
  assign n9727 = n9724 & n9732;
  assign n9714 = ~n9733;
  assign n6250 = n9734 ^ n9735;
  assign n9736 = ~n9734;
  assign n9657 = n9706 ^ n9707;
  assign n9703 = n9708 & n9709;
  assign n9692 = n9708 & n9695;
  assign n9688 = ~n9711;
  assign n9710 = n9714 & n9715;
  assign n9705 = ~n9727;
  assign n6344 = ~n6250;
  assign n9730 = n9736 & n9737;
  assign n8266 = n9692 ^ n9693;
  assign n9690 = n9657 & n9697;
  assign n9691 = ~n9657;
  assign n9694 = ~n9703;
  assign n9698 = n9672 & n9688;
  assign n9704 = ~n9710;
  assign n9699 = n6344 & n8410;
  assign n9712 = ~n9730;
  assign n9448 = ~n8266;
  assign n9673 = ~n9690;
  assign n9686 = n9691 & n483;
  assign n9675 = n9694 & n9695;
  assign n9678 = ~n9698;
  assign n9653 = n9699 ^ n7367;
  assign n9677 = n9704 & n9705;
  assign n9700 = n9712 & n9713;
  assign n9656 = n483 ^ n9675;
  assign n9670 = n9677 ^ n9678;
  assign n9659 = ~n9686;
  assign n9674 = ~n9675;
  assign n9680 = n9653 & n9689;
  assign n9681 = ~n9653;
  assign n9687 = ~n9677;
  assign n9683 = n9700 ^ n7235;
  assign n9701 = ~n9700;
  assign n9428 = n9656 ^ n9657;
  assign n9664 = n9670 & n482;
  assign n9669 = n9673 & n9674;
  assign n9662 = ~n9670;
  assign n9655 = ~n9680;
  assign n9676 = n9681 & n9639;
  assign n6181 = n9682 ^ n9683;
  assign n9679 = n9687 & n9688;
  assign n9696 = n9701 & n9702;
  assign n9433 = ~n9428;
  assign n9660 = n9662 & n9663;
  assign n9625 = ~n9664;
  assign n9658 = ~n9669;
  assign n9642 = ~n9676;
  assign n6235 = ~n6181;
  assign n9671 = ~n9679;
  assign n9684 = ~n9696;
  assign n9630 = n9658 & n9659;
  assign n9647 = ~n9660;
  assign n9649 = n6235 & n8438;
  assign n9652 = n9671 & n9672;
  assign n9666 = n9684 & n9685;
  assign n9629 = n9647 & n9625;
  assign n9643 = n9649 ^ n7235;
  assign n9646 = ~n9630;
  assign n9638 = n9652 ^ n9653;
  assign n9654 = ~n9652;
  assign n6118 = n9665 ^ n9666;
  assign n9667 = ~n9666;
  assign n9377 = n9629 ^ n9630;
  assign n9623 = n9638 ^ n9639;
  assign n9631 = n9643 & n9644;
  assign n9640 = n9646 & n9647;
  assign n9632 = ~n9643;
  assign n9648 = n9654 & n9655;
  assign n9645 = n6118 & n8389;
  assign n6120 = ~n6118;
  assign n9661 = n9667 & n9668;
  assign n9620 = n9623 & n481;
  assign n9389 = ~n9377;
  assign n9618 = ~n9623;
  assign n9603 = ~n9631;
  assign n9627 = n9632 & n9633;
  assign n9624 = ~n9640;
  assign n9585 = n9645 ^ n7216;
  assign n9641 = ~n9648;
  assign n9650 = ~n9661;
  assign n9612 = n9618 & n9619;
  assign n9596 = ~n9620;
  assign n9581 = n9624 & n9625;
  assign n9621 = n9585 & n9626;
  assign n9614 = ~n9627;
  assign n9622 = ~n9585;
  assign n9597 = n9641 & n9642;
  assign n9634 = n9650 & n9651;
  assign n9608 = ~n9612;
  assign n9611 = n9603 & n9614;
  assign n9609 = ~n9581;
  assign n9587 = ~n9621;
  assign n9615 = n9622 & n9565;
  assign n9613 = ~n9597;
  assign n6076 = n9634 ^ n9635;
  assign n9636 = ~n9634;
  assign n9600 = n9608 & n9609;
  assign n9601 = n9608 & n9596;
  assign n9598 = ~n9611;
  assign n9610 = n9613 & n9614;
  assign n9567 = ~n9615;
  assign n5982 = ~n6076;
  assign n9628 = n9636 & n9637;
  assign n9583 = n9597 ^ n9598;
  assign n9595 = ~n9600;
  assign n9582 = ~n9601;
  assign n9602 = ~n9610;
  assign n9604 = n5982 & n8298;
  assign n9616 = ~n9628;
  assign n9562 = n9581 ^ n9582;
  assign n9578 = n9583 & n480;
  assign n9540 = n9595 & n9596;
  assign n9576 = ~n9583;
  assign n9584 = n9602 & n9603;
  assign n9547 = n9604 ^ n7099;
  assign n9605 = n9616 & n9617;
  assign n9327 = n9562 ^ n9389;
  assign n9332 = n9562 ^ n9377;
  assign n9563 = ~n9562;
  assign n9574 = n9576 & n9577;
  assign n9537 = ~n9578;
  assign n9558 = ~n9540;
  assign n9564 = n9584 ^ n9585;
  assign n9588 = n9547 & n9523;
  assign n9586 = ~n9584;
  assign n9589 = ~n9547;
  assign n9592 = n9605 ^ n7067;
  assign n9606 = ~n9605;
  assign n9515 = n9563 & n9377;
  assign n9555 = n9564 ^ n9565;
  assign n9559 = ~n9574;
  assign n9579 = n9586 & n9587;
  assign n9525 = ~n9588;
  assign n9580 = n9589 & n9590;
  assign n5894 = n9591 ^ n9592;
  assign n9599 = n9606 & n9607;
  assign n9545 = n9555 & n495;
  assign n9556 = n9558 & n9559;
  assign n9543 = ~n9555;
  assign n9539 = n9559 & n9537;
  assign n9569 = n5894 & n9575;
  assign n9566 = ~n9579;
  assign n9549 = ~n9580;
  assign n5985 = ~n5894;
  assign n9593 = ~n9599;
  assign n9516 = n9539 ^ n9540;
  assign n9538 = n9543 & n9544;
  assign n9495 = ~n9545;
  assign n9536 = ~n9556;
  assign n9546 = n9566 & n9567;
  assign n9550 = n5985 & n8337;
  assign n9560 = n5985 & n9568;
  assign n8362 = ~n9569;
  assign n9571 = n9593 & n9594;
  assign n9290 = n9515 ^ n9516;
  assign n9483 = n9516 & n9515;
  assign n9501 = n9536 & n9537;
  assign n9517 = ~n9538;
  assign n9522 = n9546 ^ n9547;
  assign n9533 = n9550 ^ n7067;
  assign n9548 = ~n9546;
  assign n8383 = ~n9560;
  assign n5870 = n9570 ^ n9571;
  assign n9572 = ~n9571;
  assign n9296 = ~n9290;
  assign n9486 = ~n9483;
  assign n9500 = n9517 & n9495;
  assign n9475 = n9522 ^ n9523;
  assign n9518 = ~n9501;
  assign n9526 = n9533 & n9534;
  assign n9527 = ~n9533;
  assign n9541 = n9548 & n9549;
  assign n8380 = n8383 & n8362;
  assign n9535 = n5870 & n8304;
  assign n9552 = n5870 & n9557;
  assign n5879 = ~n5870;
  assign n9561 = n9572 & n9573;
  assign n9484 = n9500 ^ n9501;
  assign n9502 = n9475 & n9510;
  assign n9511 = n9517 & n9518;
  assign n9503 = ~n9475;
  assign n9488 = ~n9526;
  assign n9519 = n9527 & n9528;
  assign n9445 = n9535 ^ n7007;
  assign n9524 = ~n9541;
  assign n9542 = n5879 & n9551;
  assign n8342 = ~n9552;
  assign n9553 = ~n9561;
  assign n8055 = n9483 ^ n9484;
  assign n9485 = ~n9484;
  assign n9477 = ~n9502;
  assign n9496 = n9503 & n494;
  assign n9494 = ~n9511;
  assign n9505 = ~n9519;
  assign n9513 = n9445 & n9520;
  assign n9478 = n9524 & n9525;
  assign n9512 = ~n9445;
  assign n8326 = ~n9542;
  assign n9530 = n9553 & n9554;
  assign n9248 = ~n8055;
  assign n9434 = n9485 & n9486;
  assign n9474 = n9494 & n9495;
  assign n9457 = ~n9496;
  assign n9498 = n9505 & n9488;
  assign n9506 = n9512 & n9463;
  assign n9447 = ~n9513;
  assign n9504 = ~n9478;
  assign n8339 = n8342 & n8326;
  assign n5757 = n9529 ^ n9530;
  assign n9531 = ~n9530;
  assign n9437 = ~n9434;
  assign n9455 = n9474 ^ n9475;
  assign n9476 = ~n9474;
  assign n9479 = ~n9498;
  assign n9497 = n9504 & n9505;
  assign n9465 = ~n9506;
  assign n9507 = n5757 & n9514;
  assign n9493 = n5757 & n8211;
  assign n5829 = ~n5757;
  assign n9521 = n9531 & n9532;
  assign n9435 = n494 ^ n9455;
  assign n9470 = n9476 & n9477;
  assign n9439 = n9478 ^ n9479;
  assign n9480 = n9493 ^ n6951;
  assign n9487 = ~n9497;
  assign n8308 = ~n9507;
  assign n9499 = n5829 & n8287;
  assign n9508 = ~n9521;
  assign n9206 = n9434 ^ n9435;
  assign n9436 = ~n9435;
  assign n9460 = n9439 & n493;
  assign n9456 = ~n9470;
  assign n9458 = ~n9439;
  assign n9473 = n9480 & n9481;
  assign n9462 = n9487 & n9488;
  assign n9471 = ~n9480;
  assign n8290 = ~n9499;
  assign n9489 = n9508 & n9509;
  assign n9213 = ~n9206;
  assign n9390 = n9436 & n9437;
  assign n9438 = n9456 & n9457;
  assign n9454 = n9458 & n9459;
  assign n9414 = ~n9460;
  assign n9444 = n9462 ^ n9463;
  assign n9466 = n9471 & n9472;
  assign n9401 = ~n9473;
  assign n9464 = ~n9462;
  assign n9467 = n9489 ^ n9490;
  assign n9491 = ~n9489;
  assign n9412 = n9438 ^ n9439;
  assign n9373 = n9444 ^ n9445;
  assign n9440 = ~n9438;
  assign n9441 = ~n9454;
  assign n9461 = n9464 & n9465;
  assign n9426 = ~n9466;
  assign n5733 = n6925 ^ n9467;
  assign n9482 = n9491 & n9492;
  assign n9391 = n493 ^ n9412;
  assign n9422 = n9373 & n492;
  assign n9431 = n9440 & n9441;
  assign n9420 = ~n9373;
  assign n9423 = n9426 & n9401;
  assign n9432 = n5733 & n8209;
  assign n9449 = n5733 & n8266;
  assign n9446 = ~n9461;
  assign n5675 = ~n5733;
  assign n9468 = ~n9482;
  assign n7969 = n9390 ^ n9391;
  assign n9354 = n9391 & n9390;
  assign n9415 = n9420 & n9421;
  assign n9375 = ~n9422;
  assign n9413 = ~n9431;
  assign n9416 = n9432 ^ n6925;
  assign n9424 = n9446 & n9447;
  assign n9442 = n5675 & n9448;
  assign n8268 = ~n9449;
  assign n9451 = n9468 & n9469;
  assign n9168 = ~n7969;
  assign n9357 = ~n9354;
  assign n9392 = n9413 & n9414;
  assign n9393 = ~n9415;
  assign n9410 = n9416 & n9417;
  assign n9334 = n9423 ^ n9424;
  assign n9408 = ~n9416;
  assign n9425 = ~n9424;
  assign n8253 = ~n9442;
  assign n5649 = n9450 ^ n9451;
  assign n9452 = ~n9451;
  assign n9372 = n492 ^ n9392;
  assign n9394 = ~n9392;
  assign n9398 = n9334 & n9407;
  assign n9402 = n9408 & n9409;
  assign n9366 = ~n9410;
  assign n9399 = ~n9334;
  assign n9418 = n9425 & n9426;
  assign n9411 = n5649 & n8189;
  assign n9427 = n5649 & n9433;
  assign n5651 = ~n5649;
  assign n9443 = n9452 & n9453;
  assign n9355 = n9372 ^ n9373;
  assign n9386 = n9393 & n9394;
  assign n9360 = ~n9398;
  assign n9395 = n9399 & n491;
  assign n9380 = ~n9402;
  assign n9343 = n9411 ^ n6922;
  assign n9400 = ~n9418;
  assign n8234 = ~n9427;
  assign n9419 = n5651 & n9428;
  assign n9429 = ~n9443;
  assign n9123 = n9354 ^ n9355;
  assign n9356 = ~n9355;
  assign n9374 = ~n9386;
  assign n9381 = n9380 & n9366;
  assign n9336 = ~n9395;
  assign n9387 = n9343 & n9396;
  assign n9363 = n9400 & n9401;
  assign n9388 = ~n9343;
  assign n8215 = ~n9419;
  assign n9404 = n9429 & n9430;
  assign n9130 = ~n9123;
  assign n9315 = n9356 & n9357;
  assign n9358 = n9374 & n9375;
  assign n9364 = ~n9381;
  assign n9345 = ~n9387;
  assign n9382 = n9388 & n9323;
  assign n9379 = ~n9363;
  assign n8231 = n8234 & n8215;
  assign n5586 = n9403 ^ n9404;
  assign n9405 = ~n9404;
  assign n9333 = n491 ^ n9358;
  assign n9351 = n9363 ^ n9364;
  assign n9359 = ~n9358;
  assign n9376 = n9379 & n9380;
  assign n9325 = ~n9382;
  assign n9371 = n5586 & n8146;
  assign n9383 = n5586 & n9389;
  assign n5634 = ~n5586;
  assign n9397 = n9405 & n9406;
  assign n9316 = n9333 ^ n9334;
  assign n9341 = n9351 & n490;
  assign n9350 = n9359 & n9360;
  assign n9339 = ~n9351;
  assign n9307 = n9371 ^ n6898;
  assign n9365 = ~n9376;
  assign n8193 = n9377 ^ n5634;
  assign n9378 = n5634 & n9377;
  assign n8195 = ~n9383;
  assign n9384 = ~n9397;
  assign n7881 = n9315 ^ n9316;
  assign n9272 = n9316 & n9315;
  assign n9337 = n9339 & n9340;
  assign n9298 = ~n9341;
  assign n9335 = ~n9350;
  assign n9353 = n9307 & n9361;
  assign n9342 = n9365 & n9366;
  assign n9352 = ~n9307;
  assign n8173 = ~n9378;
  assign n9367 = n9384 & n9385;
  assign n9109 = ~n7881;
  assign n9275 = ~n9272;
  assign n9300 = n9335 & n9336;
  assign n9318 = ~n9337;
  assign n9322 = n9342 ^ n9343;
  assign n9346 = n9352 & n9283;
  assign n9309 = ~n9353;
  assign n9344 = ~n9342;
  assign n9347 = n9367 ^ n9368;
  assign n9369 = ~n9367;
  assign n9254 = n9322 ^ n9323;
  assign n9319 = n9318 & n9298;
  assign n9317 = ~n9300;
  assign n9338 = n9344 & n9345;
  assign n9285 = ~n9346;
  assign n5547 = n9347 ^ n6861;
  assign n9362 = n9369 & n9370;
  assign n9305 = n9254 & n489;
  assign n9314 = n9317 & n9318;
  assign n9303 = ~n9254;
  assign n9301 = ~n9319;
  assign n9326 = n5547 & n9332;
  assign n9324 = ~n9338;
  assign n5574 = ~n5547;
  assign n9348 = ~n9362;
  assign n9273 = n9300 ^ n9301;
  assign n9299 = n9303 & n9304;
  assign n9256 = ~n9305;
  assign n9297 = ~n9314;
  assign n9306 = n9324 & n9325;
  assign n9310 = n5574 & n8095;
  assign n8134 = ~n9326;
  assign n9320 = n5574 & n9327;
  assign n9328 = n9348 & n9349;
  assign n9040 = n9272 ^ n9273;
  assign n9274 = ~n9273;
  assign n9276 = n9297 & n9298;
  assign n9278 = ~n9299;
  assign n9282 = n9306 ^ n9307;
  assign n9294 = n9310 ^ n6789;
  assign n9308 = ~n9306;
  assign n8154 = ~n9320;
  assign n9311 = n9328 ^ n9329;
  assign n9330 = ~n9328;
  assign n9045 = ~n9040;
  assign n9233 = n9274 & n9275;
  assign n9253 = n489 ^ n9276;
  assign n9215 = n9282 ^ n9283;
  assign n9277 = ~n9276;
  assign n9286 = n9294 & n9295;
  assign n9287 = ~n9294;
  assign n9302 = n9308 & n9309;
  assign n8151 = n8154 & n8134;
  assign n5484 = n9311 ^ n6707;
  assign n9321 = n9330 & n9331;
  assign n9234 = n9253 ^ n9254;
  assign n9263 = n9215 & n488;
  assign n9271 = n9277 & n9278;
  assign n9261 = ~n9215;
  assign n9244 = ~n9286;
  assign n9279 = n9287 & n9288;
  assign n9289 = n5484 & n9296;
  assign n9284 = ~n9302;
  assign n5541 = ~n5484;
  assign n9312 = ~n9321;
  assign n9023 = n9233 ^ n9234;
  assign n9192 = n9234 & n9233;
  assign n9257 = n9261 & n9262;
  assign n9217 = ~n9263;
  assign n9255 = ~n9271;
  assign n9265 = ~n9279;
  assign n9238 = n9284 & n9285;
  assign n9266 = n5541 & n8061;
  assign n8092 = ~n9289;
  assign n9280 = n5541 & n9290;
  assign n9291 = n9312 & n9313;
  assign n7796 = ~n9023;
  assign n9235 = n9255 & n9256;
  assign n9237 = ~n9257;
  assign n9259 = n9265 & n9244;
  assign n9200 = n9266 ^ n6707;
  assign n9264 = ~n9238;
  assign n8112 = ~n9280;
  assign n9268 = n9291 ^ n6731;
  assign n9292 = ~n9291;
  assign n9214 = n488 ^ n9235;
  assign n9236 = ~n9235;
  assign n9247 = n9200 & n9224;
  assign n9239 = ~n9259;
  assign n9245 = ~n9200;
  assign n9258 = n9264 & n9265;
  assign n9260 = n8112 & n8092;
  assign n5508 = n9267 ^ n9268;
  assign n9281 = n9292 & n9293;
  assign n9193 = n9214 ^ n9215;
  assign n9232 = n9236 & n9237;
  assign n9222 = n9238 ^ n9239;
  assign n9240 = n9245 & n9246;
  assign n9226 = ~n9247;
  assign n9249 = n5508 & n8055;
  assign n9243 = ~n9258;
  assign n8110 = ~n9260;
  assign n5467 = ~n5508;
  assign n9269 = ~n9281;
  assign n7770 = n9192 ^ n9193;
  assign n9150 = n9193 & n9192;
  assign n9220 = n9222 & n503;
  assign n9216 = ~n9232;
  assign n9218 = ~n9222;
  assign n9202 = ~n9240;
  assign n9223 = n9243 & n9244;
  assign n9227 = n5467 & n7996;
  assign n9241 = n5467 & n9248;
  assign n8058 = ~n9249;
  assign n9250 = n9269 & n9270;
  assign n8984 = ~n7770;
  assign n9153 = ~n9150;
  assign n9178 = n9216 & n9217;
  assign n9211 = n9218 & n9219;
  assign n9175 = ~n9220;
  assign n9199 = n9223 ^ n9224;
  assign n9162 = n9227 ^ n6731;
  assign n9225 = ~n9223;
  assign n8075 = ~n9241;
  assign n9228 = n9250 ^ n6700;
  assign n9251 = ~n9250;
  assign n9155 = n9199 ^ n9200;
  assign n9194 = ~n9178;
  assign n9195 = ~n9211;
  assign n9204 = n9162 & n9212;
  assign n9203 = ~n9162;
  assign n9221 = n9225 & n9226;
  assign n5426 = n9228 ^ n9229;
  assign n9242 = n9251 & n9252;
  assign n9180 = n9155 & n9190;
  assign n9191 = n9194 & n9195;
  assign n9181 = ~n9155;
  assign n9177 = n9195 & n9175;
  assign n9196 = n9203 & n9183;
  assign n9164 = ~n9204;
  assign n9205 = n5426 & n9213;
  assign n9201 = ~n9221;
  assign n5451 = ~n5426;
  assign n9230 = ~n9242;
  assign n9151 = n9177 ^ n9178;
  assign n9157 = ~n9180;
  assign n9176 = n9181 & n502;
  assign n9174 = ~n9191;
  assign n9185 = ~n9196;
  assign n9182 = n9201 & n9202;
  assign n9186 = n5451 & n7986;
  assign n8019 = ~n9205;
  assign n9197 = n5451 & n9206;
  assign n9207 = n9230 & n9231;
  assign n8919 = n9150 ^ n9151;
  assign n9152 = ~n9151;
  assign n9154 = n9174 & n9175;
  assign n9133 = ~n9176;
  assign n9161 = n9182 ^ n9183;
  assign n9141 = n9186 ^ n6713;
  assign n9184 = ~n9182;
  assign n8037 = ~n9197;
  assign n9187 = n9207 ^ n9208;
  assign n9209 = ~n9207;
  assign n8925 = ~n8919;
  assign n9110 = n9152 & n9153;
  assign n9131 = n9154 ^ n9155;
  assign n9147 = n9161 ^ n9162;
  assign n9156 = ~n9154;
  assign n9166 = n9141 & n9173;
  assign n9165 = ~n9141;
  assign n9179 = n9184 & n9185;
  assign n8034 = n8037 & n8019;
  assign n5388 = n6641 ^ n9187;
  assign n9198 = n9209 & n9210;
  assign n9111 = n502 ^ n9131;
  assign n9139 = n9147 & n501;
  assign n9148 = n9156 & n9157;
  assign n9137 = ~n9147;
  assign n9158 = n9165 & n9118;
  assign n9143 = ~n9166;
  assign n9149 = n5388 & n7923;
  assign n9167 = n5388 & n7969;
  assign n9163 = ~n9179;
  assign n5412 = ~n5388;
  assign n9188 = ~n9198;
  assign n7629 = n9110 ^ n9111;
  assign n9068 = n9111 & n9110;
  assign n9134 = n9137 & n9138;
  assign n9091 = ~n9139;
  assign n9132 = ~n9148;
  assign n9076 = n9149 ^ n6629;
  assign n9120 = ~n9158;
  assign n9140 = n9163 & n9164;
  assign n7992 = ~n9167;
  assign n9159 = n5412 & n9168;
  assign n9169 = n9188 & n9189;
  assign n8884 = ~n7629;
  assign n9071 = ~n9068;
  assign n9088 = n9132 & n9133;
  assign n9113 = ~n9134;
  assign n9128 = n9076 & n9135;
  assign n9117 = n9140 ^ n9141;
  assign n9129 = ~n9076;
  assign n9142 = ~n9140;
  assign n7972 = ~n9159;
  assign n9144 = n9169 ^ n9170;
  assign n9171 = ~n9169;
  assign n9114 = n9113 & n9091;
  assign n9047 = n9117 ^ n9118;
  assign n9112 = ~n9088;
  assign n9079 = ~n9128;
  assign n9121 = n9129 & n9101;
  assign n9136 = n9142 & n9143;
  assign n5348 = n6568 ^ n9144;
  assign n9160 = n9171 & n9172;
  assign n9099 = n9047 & n500;
  assign n9107 = n9112 & n9113;
  assign n9089 = ~n9114;
  assign n9097 = ~n9047;
  assign n9103 = ~n9121;
  assign n9108 = n5348 & n7808;
  assign n9122 = n5348 & n9130;
  assign n9119 = ~n9136;
  assign n5350 = ~n5348;
  assign n9145 = ~n9160;
  assign n9069 = n9088 ^ n9089;
  assign n9092 = n9097 & n9098;
  assign n9049 = ~n9099;
  assign n9090 = ~n9107;
  assign n9093 = n9108 ^ n6553;
  assign n9100 = n9119 & n9120;
  assign n7951 = ~n9122;
  assign n9115 = n5350 & n9123;
  assign n9125 = n9145 & n9146;
  assign n8864 = n9068 ^ n9069;
  assign n9070 = ~n9069;
  assign n9072 = n9090 & n9091;
  assign n9074 = ~n9092;
  assign n9084 = n9093 & n9094;
  assign n9077 = n9100 ^ n9101;
  assign n9085 = ~n9093;
  assign n9102 = ~n9100;
  assign n7934 = ~n9115;
  assign n5298 = n9124 ^ n9125;
  assign n9126 = ~n9125;
  assign n8857 = ~n8864;
  assign n9028 = n9070 & n9071;
  assign n9046 = n500 ^ n9072;
  assign n9063 = n9076 ^ n9077;
  assign n9073 = ~n9072;
  assign n9038 = ~n9084;
  assign n9080 = n9085 & n9086;
  assign n9095 = n9102 & n9103;
  assign n7948 = n7951 & n7934;
  assign n9087 = n5298 & n7827;
  assign n9104 = n5298 & n9109;
  assign n5300 = ~n5298;
  assign n9116 = n9126 & n9127;
  assign n9029 = n9046 ^ n9047;
  assign n9054 = n9063 & n499;
  assign n9064 = n9073 & n9074;
  assign n9052 = ~n9063;
  assign n9056 = ~n9080;
  assign n9018 = n9087 ^ n6476;
  assign n9078 = ~n9095;
  assign n7904 = ~n9104;
  assign n9096 = n5300 & n7881;
  assign n9105 = ~n9116;
  assign n8776 = n9028 ^ n9029;
  assign n8985 = n9029 & n9028;
  assign n9050 = n9052 & n9053;
  assign n9010 = ~n9054;
  assign n9048 = ~n9064;
  assign n9057 = n9056 & n9038;
  assign n9065 = n9018 & n8994;
  assign n9035 = n9078 & n9079;
  assign n9066 = ~n9018;
  assign n7884 = ~n9096;
  assign n9081 = n9105 & n9106;
  assign n8782 = ~n8776;
  assign n8992 = ~n8985;
  assign n9007 = n9048 & n9049;
  assign n9031 = ~n9050;
  assign n9036 = ~n9057;
  assign n8996 = ~n9065;
  assign n9058 = n9066 & n9067;
  assign n9055 = ~n9035;
  assign n9060 = n9081 ^ n6419;
  assign n9082 = ~n9081;
  assign n9032 = n9031 & n9010;
  assign n9027 = n9035 ^ n9036;
  assign n9030 = ~n9007;
  assign n9051 = n9055 & n9056;
  assign n9020 = ~n9058;
  assign n5295 = n9059 ^ n9060;
  assign n9075 = n9082 & n9083;
  assign n9016 = n9027 & n498;
  assign n9026 = n9030 & n9031;
  assign n9008 = ~n9032;
  assign n9014 = ~n9027;
  assign n9039 = n5295 & n9045;
  assign n9037 = ~n9051;
  assign n5249 = ~n5295;
  assign n9061 = ~n9075;
  assign n8986 = n9007 ^ n9008;
  assign n9011 = n9014 & n9015;
  assign n8965 = ~n9016;
  assign n9009 = ~n9026;
  assign n9017 = n9037 & n9038;
  assign n9021 = n5249 & n7708;
  assign n7851 = ~n9039;
  assign n9033 = n5249 & n9040;
  assign n9041 = n9061 & n9062;
  assign n7446 = n8985 ^ n8986;
  assign n8946 = n8986 & n8992;
  assign n8967 = n9009 & n9010;
  assign n8988 = ~n9011;
  assign n8993 = n9017 ^ n9018;
  assign n9005 = n9021 ^ n6419;
  assign n9019 = ~n9017;
  assign n7869 = ~n9033;
  assign n5213 = n9041 ^ n9042;
  assign n9043 = ~n9041;
  assign n7448 = ~n7446;
  assign n8953 = ~n8946;
  assign n8949 = n8993 ^ n8994;
  assign n8989 = n8988 & n8965;
  assign n8987 = ~n8967;
  assign n8997 = n9005 & n9006;
  assign n8998 = ~n9005;
  assign n9012 = n9019 & n9020;
  assign n7866 = n7869 & n7851;
  assign n9022 = n5213 & n7796;
  assign n5253 = ~n5213;
  assign n9034 = n9043 & n9044;
  assign n8972 = n8949 & n8981;
  assign n8982 = n8987 & n8988;
  assign n8973 = ~n8949;
  assign n8968 = ~n8989;
  assign n8958 = ~n8997;
  assign n8990 = n8998 & n8999;
  assign n8995 = ~n9012;
  assign n9000 = n5253 & n7725;
  assign n7799 = ~n9022;
  assign n9013 = n5253 & n9023;
  assign n9024 = ~n9034;
  assign n8947 = n8967 ^ n8968;
  assign n8951 = ~n8972;
  assign n8966 = n8973 & n497;
  assign n8964 = ~n8982;
  assign n8975 = ~n8990;
  assign n8956 = n8995 & n8996;
  assign n8916 = n9000 ^ n6204;
  assign n7824 = ~n9013;
  assign n9001 = n9024 & n9025;
  assign n8668 = n8946 ^ n8947;
  assign n8952 = ~n8947;
  assign n8948 = n8964 & n8965;
  assign n8928 = ~n8966;
  assign n8955 = n8975 & n8958;
  assign n8977 = n8916 & n8983;
  assign n8974 = ~n8956;
  assign n8976 = ~n8916;
  assign n5150 = n9001 ^ n9002;
  assign n9003 = ~n9001;
  assign n8926 = n8948 ^ n8949;
  assign n8906 = n8952 & n8953;
  assign n8909 = n8955 ^ n8956;
  assign n8950 = ~n8948;
  assign n8969 = n8974 & n8975;
  assign n8970 = n8976 & n8935;
  assign n8918 = ~n8977;
  assign n8978 = n5150 & n8984;
  assign n5225 = ~n5150;
  assign n8991 = n9003 & n9004;
  assign n8907 = n497 ^ n8926;
  assign n8914 = ~n8906;
  assign n8932 = n8909 & n8944;
  assign n8943 = n8950 & n8951;
  assign n8933 = ~n8909;
  assign n8957 = ~n8969;
  assign n8937 = ~n8970;
  assign n8959 = n5225 & n7673;
  assign n7748 = ~n8978;
  assign n8971 = n5225 & n7770;
  assign n8979 = ~n8991;
  assign n6752 = n8906 ^ n8907;
  assign n8865 = n8907 & n8914;
  assign n8911 = ~n8932;
  assign n8929 = n8933 & n496;
  assign n8927 = ~n8943;
  assign n8934 = n8957 & n8958;
  assign n8873 = n8959 ^ n6252;
  assign n7772 = ~n8971;
  assign n8960 = n8979 & n8980;
  assign n6751 = n6735 ^ n6752;
  assign n7831 = n8885 ^ n6752;
  assign n8886 = ~n6752;
  assign n8908 = n8927 & n8928;
  assign n8889 = ~n8929;
  assign n8915 = n8934 ^ n8935;
  assign n8938 = n8873 & n8945;
  assign n8936 = ~n8934;
  assign n8939 = ~n8873;
  assign n8940 = n8960 ^ n8961;
  assign n8962 = ~n8960;
  assign n8846 = n6751 & n7817;
  assign n4953 = ~n6751;
  assign n8784 = n8886 & n6735;
  assign n8887 = n8908 ^ n8909;
  assign n8839 = n8915 ^ n8916;
  assign n8910 = ~n8908;
  assign n8930 = n8936 & n8937;
  assign n8875 = ~n8938;
  assign n8931 = n8939 & n8898;
  assign n5134 = n6174 ^ n8940;
  assign n8954 = n8962 & n8963;
  assign n8830 = n8846 ^ n8847;
  assign n8820 = n8846 ^ n8848;
  assign n8866 = n496 ^ n8887;
  assign n8896 = n8839 & n511;
  assign n8904 = n8910 & n8911;
  assign n8894 = ~n8839;
  assign n8905 = n5134 & n7640;
  assign n8920 = n5134 & n8925;
  assign n8917 = ~n8930;
  assign n8900 = ~n8931;
  assign n5185 = ~n5134;
  assign n8941 = ~n8954;
  assign n8170 = n199 ^ n8820;
  assign n8648 = n8830 & n8831;
  assign n8566 = n8820 & n199;
  assign n8849 = n8865 ^ n8866;
  assign n8812 = n8866 & n8865;
  assign n8890 = n8894 & n8895;
  assign n8841 = ~n8896;
  assign n8888 = ~n8904;
  assign n8822 = n8905 ^ n6174;
  assign n8897 = n8917 & n8918;
  assign n8912 = n5185 & n8919;
  assign n7721 = ~n8920;
  assign n8921 = n8941 & n8942;
  assign n8177 = ~n8170;
  assign n8836 = n8849 & n6665;
  assign n8837 = ~n8849;
  assign n8867 = n8888 & n8889;
  assign n8869 = ~n8890;
  assign n8882 = n8822 & n8891;
  assign n8872 = n8897 ^ n8898;
  assign n8883 = ~n8822;
  assign n8899 = ~n8897;
  assign n7700 = ~n8912;
  assign n8901 = n8921 ^ n8922;
  assign n8923 = ~n8921;
  assign n8786 = ~n8836;
  assign n8832 = n8837 & n6702;
  assign n8838 = n511 ^ n8867;
  assign n8861 = n8872 ^ n8873;
  assign n8868 = ~n8867;
  assign n8824 = ~n8882;
  assign n8876 = n8883 & n8854;
  assign n8892 = n8899 & n8900;
  assign n8893 = n7721 & n7700;
  assign n5093 = n5972 ^ n8901;
  assign n8913 = n8923 & n8924;
  assign n8811 = ~n8832;
  assign n8813 = n8838 ^ n8839;
  assign n8852 = n8861 & n510;
  assign n8862 = n8868 & n8869;
  assign n8850 = ~n8861;
  assign n8856 = ~n8876;
  assign n8863 = n5093 & n7530;
  assign n8877 = n5093 & n8884;
  assign n8874 = ~n8892;
  assign n7719 = ~n8893;
  assign n5145 = ~n5093;
  assign n8902 = ~n8913;
  assign n8807 = n8811 & n8784;
  assign n8783 = n8811 & n8786;
  assign n8795 = n8812 ^ n8813;
  assign n8814 = ~n8813;
  assign n8842 = n8850 & n8851;
  assign n8792 = ~n8852;
  assign n8840 = ~n8862;
  assign n8771 = n8863 ^ n6133;
  assign n8853 = n8874 & n8875;
  assign n8870 = n5145 & n7629;
  assign n7667 = ~n8877;
  assign n8879 = n8902 & n8903;
  assign n4934 = n8783 ^ n8784;
  assign n8788 = n8795 & n6636;
  assign n8785 = ~n8807;
  assign n8787 = ~n8795;
  assign n8761 = n8814 & n8812;
  assign n8789 = n8840 & n8841;
  assign n8816 = ~n8842;
  assign n8833 = n8771 & n8843;
  assign n8821 = n8853 ^ n8854;
  assign n8834 = ~n8771;
  assign n8855 = ~n8853;
  assign n7632 = ~n8870;
  assign n5046 = n8878 ^ n8879;
  assign n8880 = ~n8879;
  assign n4936 = ~n4934;
  assign n8731 = n8785 & n8786;
  assign n8781 = n8787 & n6646;
  assign n8760 = ~n8788;
  assign n8764 = ~n8761;
  assign n8817 = n8816 & n8792;
  assign n8766 = n8821 ^ n8822;
  assign n8815 = ~n8789;
  assign n8774 = ~n8833;
  assign n8825 = n8834 & n8800;
  assign n8844 = n8855 & n8856;
  assign n8835 = n5046 & n7357;
  assign n8858 = n5046 & n8864;
  assign n5102 = ~n5046;
  assign n8871 = n8880 & n8881;
  assign n8729 = n4936 & n7642;
  assign n8759 = ~n8731;
  assign n8733 = ~n8781;
  assign n8798 = n8766 & n509;
  assign n8808 = n8815 & n8816;
  assign n8790 = ~n8817;
  assign n8796 = ~n8766;
  assign n8802 = ~n8825;
  assign n8748 = n8835 ^ n6024;
  assign n8823 = ~n8844;
  assign n8845 = n5102 & n8857;
  assign n7598 = ~n8858;
  assign n8859 = ~n8871;
  assign n8711 = n8729 ^ n6702;
  assign n8755 = n8759 & n8760;
  assign n8730 = n8760 & n8733;
  assign n8762 = n8789 ^ n8790;
  assign n8793 = n8796 & n8797;
  assign n8738 = ~n8798;
  assign n8791 = ~n8808;
  assign n8810 = n8748 & n8818;
  assign n8799 = n8823 & n8824;
  assign n8809 = ~n8748;
  assign n7564 = ~n8845;
  assign n8826 = n8859 & n8860;
  assign n8700 = n8711 & n8712;
  assign n8698 = ~n8711;
  assign n4879 = n8730 ^ n8731;
  assign n8732 = ~n8755;
  assign n8743 = n8761 ^ n8762;
  assign n8763 = ~n8762;
  assign n8765 = n8791 & n8792;
  assign n8768 = ~n8793;
  assign n8772 = n8799 ^ n8800;
  assign n8803 = n8809 & n8714;
  assign n8750 = ~n8810;
  assign n8801 = ~n8799;
  assign n7595 = n7598 & n7564;
  assign n8804 = n8826 ^ n8827;
  assign n8828 = ~n8826;
  assign n8693 = n8698 & n8699;
  assign n8650 = ~n8700;
  assign n8686 = n4879 & n7634;
  assign n4881 = ~n4879;
  assign n8679 = n8732 & n8733;
  assign n8734 = n8743 & n6588;
  assign n8735 = ~n8743;
  assign n8703 = n8763 & n8764;
  assign n8736 = n8765 ^ n8766;
  assign n8681 = n8771 ^ n8772;
  assign n8767 = ~n8765;
  assign n8794 = n8801 & n8802;
  assign n8716 = ~n8803;
  assign n5050 = n8804 ^ n5905;
  assign n8819 = n8828 & n8829;
  assign n8669 = n8686 ^ n6636;
  assign n8674 = ~n8693;
  assign n8702 = ~n8679;
  assign n8701 = ~n8734;
  assign n8723 = n8735 & n6601;
  assign n8704 = n509 ^ n8736;
  assign n8746 = n8681 & n508;
  assign n8756 = n8767 & n8768;
  assign n8744 = ~n8681;
  assign n8775 = n5050 & n8782;
  assign n8773 = ~n8794;
  assign n5013 = ~n5050;
  assign n8805 = ~n8819;
  assign n8662 = n8669 & n8670;
  assign n8671 = n8674 & n8648;
  assign n8647 = n8674 & n8650;
  assign n8663 = ~n8669;
  assign n8694 = n8701 & n8702;
  assign n8687 = n8703 ^ n8704;
  assign n8655 = n8704 & n8703;
  assign n8676 = ~n8723;
  assign n8739 = n8744 & n8745;
  assign n8683 = ~n8746;
  assign n8737 = ~n8756;
  assign n8747 = n8773 & n8774;
  assign n8751 = n5013 & n7289;
  assign n7485 = ~n8775;
  assign n8769 = n5013 & n8776;
  assign n8778 = n8805 & n8806;
  assign n8635 = n8647 ^ n8648;
  assign n8595 = ~n8662;
  assign n8651 = n8663 & n8664;
  assign n8649 = ~n8671;
  assign n8677 = n8687 & n6517;
  assign n8675 = ~n8694;
  assign n8622 = ~n8687;
  assign n8678 = n8701 & n8676;
  assign n8705 = n8737 & n8738;
  assign n8707 = ~n8739;
  assign n8713 = n8747 ^ n8748;
  assign n8724 = n8751 ^ n5847;
  assign n8749 = ~n8747;
  assign n7521 = ~n8769;
  assign n4983 = n8777 ^ n8778;
  assign n8780 = n8778 & n8753;
  assign n8779 = ~n8778;
  assign n8618 = n8635 & n198;
  assign n8616 = ~n8635;
  assign n8592 = n8649 & n8650;
  assign n8619 = ~n8651;
  assign n8652 = n8675 & n8676;
  assign n8672 = n8622 & n6407;
  assign n8653 = ~n8677;
  assign n4830 = n8678 ^ n8679;
  assign n8680 = n508 ^ n8705;
  assign n8629 = n8713 ^ n8714;
  assign n8706 = ~n8705;
  assign n8719 = n8724 & n8725;
  assign n8717 = ~n8724;
  assign n8740 = n8749 & n8750;
  assign n8741 = n7521 & n7485;
  assign n8726 = n4983 & n7307;
  assign n4985 = ~n4983;
  assign n8770 = n8779 & n8758;
  assign n8757 = ~n8780;
  assign n8610 = n8616 & n8617;
  assign n8568 = ~n8618;
  assign n8621 = n8619 & n8595;
  assign n8620 = ~n8592;
  assign n8623 = n8652 ^ n6517;
  assign n8636 = n4830 & n7568;
  assign n8654 = ~n8652;
  assign n8625 = ~n8672;
  assign n4834 = ~n4830;
  assign n8656 = n8680 ^ n8681;
  assign n8695 = n8706 & n8707;
  assign n8708 = n8717 & n8718;
  assign n8667 = ~n8719;
  assign n8641 = n8726 ^ n5738;
  assign n8715 = ~n8740;
  assign n7519 = ~n8741;
  assign n8754 = n8757 & n8758;
  assign n8752 = ~n8770;
  assign n8591 = ~n8610;
  assign n8611 = n8619 & n8620;
  assign n8593 = ~n8621;
  assign n4783 = n8622 ^ n8623;
  assign n8612 = n8636 ^ n6588;
  assign n8644 = n8653 & n8654;
  assign n8637 = n8655 ^ n8656;
  assign n8599 = n8656 & n8655;
  assign n8682 = ~n8695;
  assign n8689 = ~n8708;
  assign n8697 = n8641 & n8709;
  assign n8660 = n8715 & n8716;
  assign n8696 = ~n8641;
  assign n8742 = n8752 & n8753;
  assign n8727 = ~n8754;
  assign n8587 = n8591 & n8566;
  assign n8565 = n8591 & n8568;
  assign n8529 = n8592 ^ n8593;
  assign n8594 = ~n8611;
  assign n8601 = n8612 & n8613;
  assign n4794 = ~n4783;
  assign n8602 = ~n8612;
  assign n8627 = n8637 & n6413;
  assign n8624 = ~n8644;
  assign n8626 = ~n8637;
  assign n8657 = n8682 & n8683;
  assign n8685 = n8689 & n8667;
  assign n8690 = n8696 & n8607;
  assign n8643 = ~n8697;
  assign n8688 = ~n8660;
  assign n8720 = n8727 & n8728;
  assign n8721 = ~n8742;
  assign n8131 = n8565 ^ n8566;
  assign n8567 = ~n8587;
  assign n8556 = n8594 & n8595;
  assign n8569 = n4794 & n7477;
  assign n8546 = ~n8601;
  assign n8596 = n8602 & n8603;
  assign n8562 = n8624 & n8625;
  assign n8614 = n8626 & n6424;
  assign n8598 = ~n8627;
  assign n8628 = n507 ^ n8657;
  assign n8659 = n8657 & n8665;
  assign n8658 = ~n8657;
  assign n8661 = ~n8685;
  assign n8684 = n8688 & n8689;
  assign n8609 = ~n8690;
  assign n8692 = ~n8720;
  assign n8710 = n8721 & n8722;
  assign n8138 = ~n8131;
  assign n8553 = n8567 & n8568;
  assign n8497 = n8569 ^ n6517;
  assign n8571 = ~n8556;
  assign n8570 = ~n8596;
  assign n8597 = ~n8562;
  assign n8573 = ~n8614;
  assign n8600 = n8628 ^ n8629;
  assign n8645 = n8658 & n507;
  assign n8638 = ~n8659;
  assign n8639 = n8660 ^ n8661;
  assign n8666 = ~n8684;
  assign n8691 = ~n8710;
  assign n8541 = n8553 & n8554;
  assign n8544 = n8497 & n8517;
  assign n8536 = ~n8553;
  assign n8542 = ~n8497;
  assign n8561 = n8570 & n8571;
  assign n8555 = n8570 & n8546;
  assign n8588 = n8597 & n8598;
  assign n8589 = n8598 & n8573;
  assign n8579 = n8599 ^ n8600;
  assign n8551 = n8600 & n8599;
  assign n8630 = n8638 & n8629;
  assign n8633 = n8639 & n506;
  assign n8605 = ~n8645;
  assign n8631 = ~n8639;
  assign n8640 = n8666 & n8667;
  assign n4926 = n8691 & n8692;
  assign n8514 = n8536 ^ n8529;
  assign n8537 = n8536 & n197;
  assign n8528 = ~n8541;
  assign n8538 = n8542 & n8543;
  assign n8503 = ~n8544;
  assign n8462 = n8555 ^ n8556;
  assign n8545 = ~n8561;
  assign n8574 = n8579 & n6344;
  assign n8572 = ~n8588;
  assign n8563 = ~n8589;
  assign n8548 = ~n8579;
  assign n8604 = ~n8630;
  assign n8615 = n8631 & n8632;
  assign n8558 = ~n8633;
  assign n8606 = n8640 ^ n8641;
  assign n8642 = ~n8640;
  assign n7330 = n8668 ^ n4926;
  assign n8646 = n4926 & n8673;
  assign n5798 = ~n4926;
  assign n8089 = n197 ^ n8514;
  assign n8521 = n8528 & n8529;
  assign n8509 = ~n8537;
  assign n8520 = ~n8538;
  assign n8539 = n8545 & n8546;
  assign n8472 = ~n8462;
  assign n4750 = n8562 ^ n8563;
  assign n8547 = n8572 & n8573;
  assign n8564 = n8548 & n6250;
  assign n8550 = ~n8574;
  assign n8576 = n8604 & n8605;
  assign n8590 = n8606 ^ n8607;
  assign n8581 = ~n8615;
  assign n8634 = n8642 & n8643;
  assign n8560 = n8646 ^ n5715;
  assign n7345 = ~n7330;
  assign n8097 = ~n8089;
  assign n8508 = ~n8521;
  assign n8516 = ~n8539;
  assign n8522 = n8547 ^ n8548;
  assign n4763 = ~n4750;
  assign n8549 = ~n8547;
  assign n8524 = ~n8564;
  assign n8584 = n8590 & n505;
  assign n8580 = ~n8576;
  assign n8582 = ~n8590;
  assign n8575 = n8581 & n8558;
  assign n8608 = ~n8634;
  assign n8486 = n8508 & n8509;
  assign n8496 = n8516 ^ n8517;
  assign n8515 = n8520 & n8516;
  assign n4712 = n6250 ^ n8522;
  assign n8518 = n4763 & n7427;
  assign n8540 = n8549 & n8550;
  assign n8552 = n8575 ^ n8576;
  assign n8577 = n8580 & n8581;
  assign n8578 = n8582 & n8583;
  assign n8513 = ~n8584;
  assign n8585 = n8608 & n8609;
  assign n8461 = n196 ^ n8486;
  assign n8488 = n8486 & n8495;
  assign n8479 = n8496 ^ n8497;
  assign n8487 = ~n8486;
  assign n8489 = n4712 & n7367;
  assign n8502 = ~n8515;
  assign n4714 = ~n4712;
  assign n8504 = n8518 ^ n6413;
  assign n8523 = ~n8540;
  assign n8530 = n8551 ^ n8552;
  assign n8510 = n8552 & n8551;
  assign n8557 = ~n8577;
  assign n8535 = ~n8578;
  assign n8559 = n8585 ^ n8586;
  assign n8443 = n8461 ^ n8462;
  assign n8476 = n8479 & n195;
  assign n8480 = n8487 & n196;
  assign n8471 = ~n8488;
  assign n8473 = ~n8479;
  assign n8433 = n8489 ^ n6250;
  assign n8445 = n8502 & n8503;
  assign n8498 = n8504 & n8505;
  assign n8499 = ~n8504;
  assign n8484 = n8523 & n8524;
  assign n8525 = n8530 & n6235;
  assign n8526 = ~n8530;
  assign n8533 = n8557 & n8558;
  assign n8532 = n8535 & n8513;
  assign n8531 = n8559 ^ n8560;
  assign n6799 = n8443 ^ n8089;
  assign n8403 = n8443 & n8089;
  assign n8463 = n8471 & n8472;
  assign n8464 = n8473 & n8474;
  assign n8466 = n8433 & n8475;
  assign n8412 = ~n8476;
  assign n8451 = ~n8480;
  assign n8465 = ~n8433;
  assign n8478 = ~n8445;
  assign n8453 = ~n8498;
  assign n8490 = n8499 & n8500;
  assign n8506 = ~n8484;
  assign n8507 = ~n8525;
  assign n8519 = n8526 & n6181;
  assign n8494 = n504 ^ n8531;
  assign n8511 = n8532 ^ n8533;
  assign n8534 = ~n8533;
  assign n8040 = ~n6799;
  assign n8406 = ~n8403;
  assign n8450 = ~n8463;
  assign n8431 = ~n8464;
  assign n8456 = n8465 & n8410;
  assign n8434 = ~n8466;
  assign n8477 = ~n8490;
  assign n8501 = n8506 & n8507;
  assign n8458 = n8510 ^ n8511;
  assign n8469 = n8511 & n8510;
  assign n8482 = ~n8519;
  assign n8527 = n8534 & n8535;
  assign n8420 = n8450 & n8451;
  assign n8444 = n8431 & n8412;
  assign n8414 = ~n8456;
  assign n8467 = n8477 & n8478;
  assign n8468 = n8477 & n8453;
  assign n8481 = ~n8501;
  assign n8491 = n8458 & n6118;
  assign n8483 = n8507 & n8482;
  assign n8492 = ~n8458;
  assign n8512 = ~n8527;
  assign n8430 = ~n8420;
  assign n8421 = ~n8444;
  assign n8452 = ~n8467;
  assign n8446 = ~n8468;
  assign n8457 = n8481 & n8482;
  assign n4671 = n8483 ^ n8484;
  assign n8460 = ~n8491;
  assign n8485 = n8492 & n6120;
  assign n8493 = n8512 & n8513;
  assign n8404 = n8420 ^ n8421;
  assign n8422 = n8430 & n8431;
  assign n8436 = n8445 ^ n8446;
  assign n8432 = n8452 & n8453;
  assign n8439 = n8457 ^ n8458;
  assign n8447 = n4671 & n7247;
  assign n8459 = ~n8457;
  assign n4673 = ~n4671;
  assign n8441 = ~n8485;
  assign n8470 = n8493 ^ n8494;
  assign n8021 = n8403 ^ n8404;
  assign n8405 = ~n8404;
  assign n8411 = ~n8422;
  assign n8409 = n8432 ^ n8433;
  assign n8426 = n8436 & n194;
  assign n4626 = n8439 ^ n6120;
  assign n8424 = ~n8436;
  assign n8435 = ~n8432;
  assign n8437 = n8447 ^ n6235;
  assign n8454 = n8459 & n8460;
  assign n8455 = n8469 ^ n8470;
  assign n8016 = ~n8021;
  assign n8363 = n8405 & n8406;
  assign n8398 = n8409 ^ n8410;
  assign n8386 = n8411 & n8412;
  assign n8416 = n8424 & n8425;
  assign n8369 = ~n8426;
  assign n8423 = n8434 & n8435;
  assign n8427 = n8437 & n8438;
  assign n4649 = ~n4626;
  assign n8428 = ~n8437;
  assign n8440 = ~n8454;
  assign n8449 = n8455 & n5982;
  assign n8448 = ~n8455;
  assign n8393 = n8398 & n193;
  assign n8366 = ~n8363;
  assign n8391 = ~n8398;
  assign n8394 = ~n8386;
  assign n8395 = ~n8416;
  assign n8399 = n4649 & n7216;
  assign n8413 = ~n8423;
  assign n8371 = ~n8427;
  assign n8417 = n8428 & n8429;
  assign n8408 = n8440 & n8441;
  assign n8442 = n8448 & n6076;
  assign n8419 = ~n8449;
  assign n8384 = n8391 & n8392;
  assign n8332 = ~n8393;
  assign n8387 = n8394 & n8395;
  assign n8388 = n8399 ^ n6118;
  assign n8385 = n8395 & n8369;
  assign n8378 = n8413 & n8414;
  assign n8397 = ~n8417;
  assign n8418 = ~n8408;
  assign n8402 = ~n8442;
  assign n8349 = ~n8384;
  assign n8364 = n8385 ^ n8386;
  assign n8368 = ~n8387;
  assign n8377 = n8388 & n8389;
  assign n8375 = ~n8388;
  assign n8396 = ~n8378;
  assign n8400 = n8397 & n8371;
  assign n8415 = n8418 & n8419;
  assign n8407 = n8419 & n8402;
  assign n7947 = n8363 ^ n8364;
  assign n8367 = n8349 & n8332;
  assign n8343 = n8368 & n8369;
  assign n8365 = ~n8364;
  assign n8372 = n8375 & n8376;
  assign n8336 = ~n8377;
  assign n8390 = n8396 & n8397;
  assign n8379 = ~n8400;
  assign n4589 = n8407 ^ n8408;
  assign n8401 = ~n8415;
  assign n7955 = ~n7947;
  assign n8327 = n8365 & n8366;
  assign n8344 = ~n8367;
  assign n8350 = ~n8343;
  assign n8352 = ~n8372;
  assign n8296 = n8378 ^ n8379;
  assign n8370 = ~n8390;
  assign n8373 = n4589 & n7120;
  assign n8381 = n8401 & n8402;
  assign n4613 = ~n4589;
  assign n8328 = n8343 ^ n8344;
  assign n8345 = n8349 & n8350;
  assign n8354 = n8352 & n8336;
  assign n8359 = n8296 & n192;
  assign n8333 = n8370 & n8371;
  assign n8357 = ~n8296;
  assign n8320 = n8373 ^ n6076;
  assign n4550 = n8380 ^ n8381;
  assign n8382 = ~n8381;
  assign n7931 = n8327 ^ n8328;
  assign n8274 = n8328 & n8327;
  assign n8331 = ~n8345;
  assign n8334 = ~n8354;
  assign n8353 = n8357 & n8358;
  assign n8300 = ~n8359;
  assign n8356 = n8320 & n8360;
  assign n8351 = ~n8333;
  assign n8347 = n4550 & n7076;
  assign n8355 = ~n8320;
  assign n4582 = ~n4550;
  assign n8374 = n8382 & n8383;
  assign n7936 = ~n7931;
  assign n8313 = n8331 & n8332;
  assign n8323 = n8333 ^ n8334;
  assign n8258 = n8347 ^ n5985;
  assign n8346 = n8351 & n8352;
  assign n8315 = ~n8353;
  assign n8348 = n8355 & n8298;
  assign n8322 = ~n8356;
  assign n8361 = ~n8374;
  assign n8295 = n192 ^ n8313;
  assign n8318 = n8323 & n207;
  assign n8314 = ~n8313;
  assign n8316 = ~n8323;
  assign n8330 = n8258 & n8337;
  assign n8329 = ~n8258;
  assign n8335 = ~n8346;
  assign n8302 = ~n8348;
  assign n8340 = n8361 & n8362;
  assign n8275 = n8295 ^ n8296;
  assign n8309 = n8314 & n8315;
  assign n8310 = n8316 & n8317;
  assign n8261 = ~n8318;
  assign n8324 = n8329 & n8283;
  assign n8263 = ~n8330;
  assign n8319 = n8335 & n8336;
  assign n4509 = n8339 ^ n8340;
  assign n8341 = ~n8340;
  assign n6556 = n8274 ^ n8275;
  assign n8276 = ~n8275;
  assign n8299 = ~n8309;
  assign n8280 = ~n8310;
  assign n8297 = n8319 ^ n8320;
  assign n8285 = ~n8324;
  assign n8321 = ~n8319;
  assign n8312 = n4509 & n7017;
  assign n4536 = ~n4509;
  assign n8338 = n8341 & n8342;
  assign n7872 = ~n6556;
  assign n8254 = n8276 & n8274;
  assign n8242 = n8297 ^ n8298;
  assign n8270 = n8299 & n8300;
  assign n8291 = n8280 & n8261;
  assign n8303 = n8312 ^ n5870;
  assign n8311 = n8321 & n8322;
  assign n8325 = ~n8338;
  assign n8257 = ~n8254;
  assign n8279 = n8242 & n206;
  assign n8277 = ~n8242;
  assign n8281 = ~n8270;
  assign n8271 = ~n8291;
  assign n8292 = n8303 & n8304;
  assign n8293 = ~n8303;
  assign n8301 = ~n8311;
  assign n8306 = n8325 & n8326;
  assign n8255 = n8270 ^ n8271;
  assign n8269 = n8277 & n8278;
  assign n8220 = ~n8279;
  assign n8272 = n8280 & n8281;
  assign n8224 = ~n8292;
  assign n8286 = n8293 & n8294;
  assign n8282 = n8301 & n8302;
  assign n8288 = n8306 ^ n5757;
  assign n8307 = ~n8306;
  assign n7853 = n8254 ^ n8255;
  assign n8256 = ~n8255;
  assign n8243 = ~n8269;
  assign n8260 = ~n8272;
  assign n8259 = n8282 ^ n8283;
  assign n8248 = ~n8286;
  assign n4466 = n8287 ^ n8288;
  assign n8284 = ~n8282;
  assign n8305 = n8307 & n8308;
  assign n7848 = ~n7853;
  assign n8202 = n8256 & n8257;
  assign n8249 = n8258 ^ n8259;
  assign n8241 = n8260 & n8261;
  assign n8245 = n8248 & n8224;
  assign n8273 = n8284 & n8285;
  assign n4495 = ~n4466;
  assign n8289 = ~n8305;
  assign n8218 = n8241 ^ n8242;
  assign n8240 = n8249 & n205;
  assign n8238 = ~n8249;
  assign n8244 = ~n8241;
  assign n8250 = n4495 & n6995;
  assign n8262 = ~n8273;
  assign n8265 = n8289 & n8290;
  assign n8203 = n206 ^ n8218;
  assign n8235 = n8238 & n8239;
  assign n8185 = ~n8240;
  assign n8236 = n8243 & n8244;
  assign n8183 = n8250 ^ n5757;
  assign n8246 = n8262 & n8263;
  assign n8251 = n8265 ^ n8266;
  assign n8267 = ~n8265;
  assign n7777 = n8202 ^ n8203;
  assign n8178 = n8203 & n8202;
  assign n8207 = ~n8235;
  assign n8219 = ~n8236;
  assign n8230 = n8183 & n8211;
  assign n8140 = n8245 ^ n8246;
  assign n8228 = ~n8183;
  assign n4424 = n8251 ^ n5733;
  assign n8247 = ~n8246;
  assign n8264 = n8267 & n8268;
  assign n7767 = ~n7777;
  assign n8181 = ~n8178;
  assign n8204 = n8207 & n8185;
  assign n8205 = n8219 & n8220;
  assign n8221 = n8140 & n8227;
  assign n8225 = n8228 & n8229;
  assign n8187 = ~n8230;
  assign n8222 = ~n8140;
  assign n8217 = n4424 & n6968;
  assign n8237 = n8247 & n8248;
  assign n4469 = ~n4424;
  assign n8252 = ~n8264;
  assign n8179 = n8204 ^ n8205;
  assign n8206 = ~n8205;
  assign n8208 = n8217 ^ n5733;
  assign n8163 = ~n8221;
  assign n8216 = n8222 & n204;
  assign n8212 = ~n8225;
  assign n8223 = ~n8237;
  assign n8232 = n8252 & n8253;
  assign n7729 = n8178 ^ n8179;
  assign n8180 = ~n8179;
  assign n8196 = n8206 & n8207;
  assign n8199 = n8208 & n8209;
  assign n8197 = ~n8208;
  assign n8142 = ~n8216;
  assign n8210 = n8223 & n8224;
  assign n4379 = n8231 ^ n8232;
  assign n8233 = ~n8232;
  assign n7717 = ~n7729;
  assign n8116 = n8180 & n8181;
  assign n8184 = ~n8196;
  assign n8191 = n8197 & n8198;
  assign n8144 = ~n8199;
  assign n8182 = n8210 ^ n8211;
  assign n8213 = ~n8210;
  assign n8201 = n4379 & n6922;
  assign n4416 = ~n4379;
  assign n8226 = n8233 & n8234;
  assign n8099 = n8182 ^ n8183;
  assign n8161 = n8184 & n8185;
  assign n8165 = ~n8191;
  assign n8188 = n8201 ^ n5649;
  assign n8200 = n8212 & n8213;
  assign n8214 = ~n8226;
  assign n8139 = n204 ^ n8161;
  assign n8159 = n8099 & n8167;
  assign n8160 = ~n8099;
  assign n8162 = ~n8161;
  assign n8168 = n8165 & n8144;
  assign n8174 = n8188 & n8189;
  assign n8175 = ~n8188;
  assign n8186 = ~n8200;
  assign n8192 = n8214 & n8215;
  assign n8117 = n8139 ^ n8140;
  assign n8120 = ~n8159;
  assign n8155 = n8160 & n203;
  assign n8156 = n8162 & n8163;
  assign n8150 = ~n8168;
  assign n8105 = ~n8174;
  assign n8169 = n8175 & n8176;
  assign n8149 = n8186 & n8187;
  assign n4337 = n8192 ^ n8193;
  assign n8194 = ~n8192;
  assign n6295 = n8116 ^ n8117;
  assign n8078 = n8117 & n8116;
  assign n8063 = n8149 ^ n8150;
  assign n8101 = ~n8155;
  assign n8141 = ~n8156;
  assign n8125 = ~n8169;
  assign n8164 = ~n8149;
  assign n8158 = n4337 & n6898;
  assign n8171 = n4337 & n8177;
  assign n4370 = ~n4337;
  assign n8190 = n8194 & n8195;
  assign n7697 = ~n6295;
  assign n8129 = n8063 & n202;
  assign n8118 = n8141 & n8142;
  assign n8127 = ~n8063;
  assign n8122 = n8125 & n8105;
  assign n8145 = n8158 ^ n5586;
  assign n8157 = n8164 & n8165;
  assign n8166 = n4370 & n8170;
  assign n6944 = ~n8171;
  assign n8172 = ~n8190;
  assign n8098 = n203 ^ n8118;
  assign n8121 = n8127 & n8128;
  assign n8065 = ~n8129;
  assign n8119 = ~n8118;
  assign n8135 = n8145 & n8146;
  assign n8136 = ~n8145;
  assign n8143 = ~n8157;
  assign n6931 = ~n8166;
  assign n8152 = n8172 & n8173;
  assign n8079 = n8098 ^ n8099;
  assign n8113 = n8119 & n8120;
  assign n8082 = ~n8121;
  assign n8070 = ~n8135;
  assign n8130 = n8136 & n8137;
  assign n8123 = n8143 & n8144;
  assign n8147 = n6944 & n6931;
  assign n4298 = n8151 ^ n8152;
  assign n8153 = ~n8152;
  assign n7607 = n8078 ^ n8079;
  assign n8041 = n8079 & n8078;
  assign n8100 = ~n8113;
  assign n8023 = n8122 ^ n8123;
  assign n8086 = ~n8130;
  assign n8124 = ~n8123;
  assign n8115 = n4298 & n6861;
  assign n8132 = n4298 & n8138;
  assign n6942 = ~n8147;
  assign n4359 = ~n4298;
  assign n8148 = n8153 & n8154;
  assign n7593 = ~n7607;
  assign n8080 = n8100 & n8101;
  assign n8102 = n8023 & n8107;
  assign n8103 = ~n8023;
  assign n8108 = n8086 & n8070;
  assign n8025 = n8115 ^ n5547;
  assign n8114 = n8124 & n8125;
  assign n8126 = n4359 & n8131;
  assign n6909 = ~n8132;
  assign n8133 = ~n8148;
  assign n8062 = n202 ^ n8080;
  assign n8081 = ~n8080;
  assign n8046 = ~n8102;
  assign n8093 = n8103 & n201;
  assign n8096 = n8025 & n8048;
  assign n8084 = ~n8108;
  assign n8094 = ~n8025;
  assign n8104 = ~n8114;
  assign n6890 = ~n8126;
  assign n8109 = n8133 & n8134;
  assign n8042 = n8062 ^ n8063;
  assign n8076 = n8081 & n8082;
  assign n8027 = ~n8093;
  assign n8088 = n8094 & n8095;
  assign n8050 = ~n8096;
  assign n8083 = n8104 & n8105;
  assign n6906 = n6909 & n6890;
  assign n4235 = n8109 ^ n8110;
  assign n8111 = ~n8109;
  assign n6147 = n8041 ^ n8042;
  assign n8043 = ~n8042;
  assign n8064 = ~n8076;
  assign n8007 = n8083 ^ n8084;
  assign n8029 = ~n8088;
  assign n6867 = n8089 ^ n4235;
  assign n8085 = ~n8083;
  assign n8090 = n4235 & n8097;
  assign n4262 = ~n4235;
  assign n8106 = n8111 & n8112;
  assign n7562 = ~n6147;
  assign n8000 = n8043 & n8041;
  assign n8044 = n8064 & n8065;
  assign n8068 = n8007 & n200;
  assign n8066 = ~n8007;
  assign n8077 = n8085 & n8086;
  assign n8072 = n4262 & n6707;
  assign n8087 = n4262 & n8089;
  assign n6849 = ~n8090;
  assign n8091 = ~n8106;
  assign n8003 = ~n8000;
  assign n8022 = n201 ^ n8044;
  assign n8045 = ~n8044;
  assign n8059 = n8066 & n8067;
  assign n7979 = ~n8068;
  assign n8060 = n8072 ^ n5541;
  assign n8069 = ~n8077;
  assign n6869 = ~n8087;
  assign n8073 = n8091 & n8092;
  assign n8001 = n8022 ^ n8023;
  assign n8038 = n8045 & n8046;
  assign n8009 = ~n8059;
  assign n8052 = n8060 & n8061;
  assign n8047 = n8069 & n8070;
  assign n8053 = ~n8060;
  assign n8056 = n8073 ^ n5508;
  assign n8074 = ~n8073;
  assign n6072 = n8000 ^ n8001;
  assign n8002 = ~n8001;
  assign n8026 = ~n8038;
  assign n8024 = n8047 ^ n8048;
  assign n7984 = ~n8052;
  assign n8051 = n8053 & n8054;
  assign n4198 = n8055 ^ n8056;
  assign n8049 = ~n8047;
  assign n8071 = n8074 & n8075;
  assign n7494 = ~n6072;
  assign n7956 = n8002 & n8003;
  assign n7961 = n8024 ^ n8025;
  assign n8006 = n8026 & n8027;
  assign n8020 = n4198 & n6741;
  assign n8033 = n4198 & n8040;
  assign n8039 = n8049 & n8050;
  assign n8013 = ~n8051;
  assign n4249 = ~n4198;
  assign n8057 = ~n8071;
  assign n7959 = ~n7956;
  assign n7977 = n8006 ^ n8007;
  assign n8004 = n7961 & n8015;
  assign n8005 = ~n7961;
  assign n8008 = ~n8006;
  assign n7939 = n8020 ^ n5508;
  assign n8030 = n8013 & n7984;
  assign n6828 = ~n8033;
  assign n8031 = n4249 & n6799;
  assign n8028 = ~n8039;
  assign n8035 = n8057 & n8058;
  assign n7957 = n200 ^ n7977;
  assign n7962 = ~n8004;
  assign n7993 = n8005 & n215;
  assign n7994 = n8008 & n8009;
  assign n7997 = n7939 & n7965;
  assign n7995 = ~n7939;
  assign n8010 = n8028 & n8029;
  assign n8011 = ~n8030;
  assign n6801 = ~n8031;
  assign n4156 = n8034 ^ n8035;
  assign n8036 = ~n8035;
  assign n5957 = n7956 ^ n7957;
  assign n7958 = ~n7957;
  assign n7941 = ~n7993;
  assign n7978 = ~n7994;
  assign n7989 = n7995 & n7996;
  assign n7967 = ~n7997;
  assign n7988 = n8010 ^ n8011;
  assign n8012 = ~n8010;
  assign n7999 = n4156 & n6713;
  assign n8017 = n4156 & n8021;
  assign n4202 = ~n4156;
  assign n8032 = n8036 & n8037;
  assign n6004 = ~n5957;
  assign n7912 = n7958 & n7959;
  assign n7960 = n7978 & n7979;
  assign n7982 = n7988 & n214;
  assign n7943 = ~n7989;
  assign n7980 = ~n7988;
  assign n7985 = n7999 ^ n5451;
  assign n7998 = n8012 & n8013;
  assign n8014 = n4202 & n8016;
  assign n6772 = ~n8017;
  assign n8018 = ~n8032;
  assign n7915 = ~n7912;
  assign n7937 = n7960 ^ n7961;
  assign n7963 = ~n7960;
  assign n7973 = n7980 & n7981;
  assign n7893 = ~n7982;
  assign n7974 = n7985 & n7986;
  assign n7975 = ~n7985;
  assign n7983 = ~n7998;
  assign n6749 = ~n8014;
  assign n7990 = n8018 & n8019;
  assign n7913 = n215 ^ n7937;
  assign n7952 = n7962 & n7963;
  assign n7921 = ~n7973;
  assign n7897 = ~n7974;
  assign n7968 = n7975 & n7976;
  assign n7964 = n7983 & n7984;
  assign n6769 = n6772 & n6749;
  assign n7970 = n7990 ^ n5388;
  assign n7991 = ~n7990;
  assign n7258 = n7912 ^ n7913;
  assign n7914 = ~n7913;
  assign n7940 = ~n7952;
  assign n7953 = n7921 & n7893;
  assign n7938 = n7964 ^ n7965;
  assign n7927 = ~n7968;
  assign n4111 = n7969 ^ n7970;
  assign n7966 = ~n7964;
  assign n7987 = n7991 & n7992;
  assign n7889 = n7914 & n7915;
  assign n7856 = n7938 ^ n7939;
  assign n7918 = n7940 & n7941;
  assign n7919 = ~n7953;
  assign n7924 = n7927 & n7897;
  assign n7935 = n4111 & n6641;
  assign n7946 = n4111 & n7955;
  assign n7954 = n7966 & n7967;
  assign n4171 = ~n4111;
  assign n7971 = ~n7987;
  assign n7891 = ~n7889;
  assign n7890 = n7918 ^ n7919;
  assign n7916 = n7856 & n7930;
  assign n7917 = ~n7856;
  assign n7920 = ~n7918;
  assign n7922 = n7935 ^ n5388;
  assign n6719 = ~n7946;
  assign n7944 = n4171 & n7947;
  assign n7942 = ~n7954;
  assign n7949 = n7971 & n7972;
  assign n6803 = n7889 ^ n7890;
  assign n7832 = n7890 & n7891;
  assign n7875 = ~n7916;
  assign n7905 = n7917 & n213;
  assign n7906 = n7920 & n7921;
  assign n7907 = n7922 & n7923;
  assign n7908 = ~n7922;
  assign n7925 = n7942 & n7943;
  assign n6691 = ~n7944;
  assign n4070 = n7948 ^ n7949;
  assign n7950 = ~n7949;
  assign n3807 = n6803 ^ n6751;
  assign n7873 = ~n6803;
  assign n7858 = ~n7905;
  assign n7892 = ~n7906;
  assign n7860 = ~n7907;
  assign n7901 = n7908 & n7909;
  assign n7835 = n7924 ^ n7925;
  assign n7928 = n6719 & n6691;
  assign n7926 = ~n7925;
  assign n7911 = n4070 & n6568;
  assign n7932 = n4070 & n7936;
  assign n4121 = ~n4070;
  assign n7945 = n7950 & n7951;
  assign n7854 = ~n3807;
  assign n6829 = n7873 & n4953;
  assign n7874 = n7892 & n7893;
  assign n7894 = n7835 & n7900;
  assign n7878 = ~n7901;
  assign n7895 = ~n7835;
  assign n7840 = n7911 ^ n5348;
  assign n7910 = n7926 & n7927;
  assign n6717 = ~n7928;
  assign n7929 = n4121 & n7931;
  assign n6663 = ~n7932;
  assign n7933 = ~n7945;
  assign n7830 = n7854 & n6735;
  assign n7855 = n213 ^ n7874;
  assign n7876 = ~n7874;
  assign n7879 = n7878 & n7860;
  assign n7837 = ~n7894;
  assign n7885 = n7895 & n212;
  assign n7886 = n7840 & n7808;
  assign n7887 = ~n7840;
  assign n7896 = ~n7910;
  assign n6631 = ~n7929;
  assign n7902 = n7933 & n7934;
  assign n7816 = n7830 ^ n6751;
  assign n7803 = n7830 ^ n7831;
  assign n7833 = n7855 ^ n7856;
  assign n7870 = n7875 & n7876;
  assign n7864 = ~n7879;
  assign n7810 = ~n7885;
  assign n7812 = ~n7886;
  assign n7880 = n7887 & n7888;
  assign n7863 = n7896 & n7897;
  assign n7898 = n6663 & n6631;
  assign n7882 = n7902 ^ n5298;
  assign n7903 = ~n7902;
  assign n5413 = n423 ^ n7803;
  assign n7675 = n7816 & n7817;
  assign n7547 = n7803 & n423;
  assign n7818 = n7832 ^ n7833;
  assign n7780 = n7833 & n7832;
  assign n7852 = n7863 ^ n7864;
  assign n7857 = ~n7870;
  assign n7842 = ~n7880;
  assign n4015 = n7881 ^ n7882;
  assign n7877 = ~n7863;
  assign n6661 = ~n7898;
  assign n7899 = n7903 & n7904;
  assign n7793 = n7675 & n7642;
  assign n5441 = ~n5413;
  assign n7791 = ~n7675;
  assign n7805 = n7818 & n4934;
  assign n7804 = ~n7818;
  assign n7846 = n7852 & n211;
  assign n7834 = n7857 & n7858;
  assign n7844 = ~n7852;
  assign n7865 = n4015 & n7872;
  assign n7871 = n7877 & n7878;
  assign n4106 = ~n4015;
  assign n7883 = ~n7899;
  assign n7778 = n7791 & n7792;
  assign n7658 = ~n7793;
  assign n7800 = n7804 & n4936;
  assign n7753 = ~n7805;
  assign n7806 = n7834 ^ n7835;
  assign n7838 = n7844 & n7845;
  assign n7760 = ~n7846;
  assign n7836 = ~n7834;
  assign n7847 = n4106 & n6356;
  assign n6558 = ~n7865;
  assign n7861 = n4106 & n6556;
  assign n7859 = ~n7871;
  assign n7867 = n7883 & n7884;
  assign n7694 = ~n7778;
  assign n7779 = ~n7800;
  assign n7781 = n212 ^ n7806;
  assign n7825 = n7836 & n7837;
  assign n7787 = ~n7838;
  assign n7826 = n7847 ^ n5298;
  assign n7839 = n7859 & n7860;
  assign n6596 = ~n7861;
  assign n4044 = n7866 ^ n7867;
  assign n7868 = ~n7867;
  assign n7773 = n7779 & n6829;
  assign n7751 = n7779 & n7753;
  assign n7731 = n7780 ^ n7781;
  assign n7756 = n7781 & n7780;
  assign n7784 = n7787 & n7760;
  assign n7809 = ~n7825;
  assign n7819 = n7826 & n7827;
  assign n7807 = n7839 ^ n7840;
  assign n7820 = ~n7826;
  assign n7841 = ~n7839;
  assign n7829 = n4044 & n6437;
  assign n7849 = n4044 & n7853;
  assign n4055 = ~n4044;
  assign n7862 = n7868 & n7869;
  assign n3710 = n7751 ^ n6829;
  assign n7755 = n7731 & n4881;
  assign n7752 = ~n7773;
  assign n7754 = ~n7731;
  assign n7735 = n7807 ^ n7808;
  assign n7785 = n7809 & n7810;
  assign n7764 = ~n7819;
  assign n7813 = n7820 & n7821;
  assign n7742 = n7829 ^ n5295;
  assign n7828 = n7841 & n7842;
  assign n7843 = n4055 & n7848;
  assign n6525 = ~n7849;
  assign n7850 = ~n7862;
  assign n3768 = ~n3710;
  assign n7730 = n7752 & n7753;
  assign n7749 = n7754 & n4879;
  assign n7705 = ~n7755;
  assign n7757 = n7784 ^ n7785;
  assign n7782 = n7735 & n7794;
  assign n7783 = ~n7735;
  assign n7786 = ~n7785;
  assign n7788 = ~n7813;
  assign n7802 = n7742 & n7814;
  assign n7801 = ~n7742;
  assign n7811 = ~n7828;
  assign n6489 = ~n7843;
  assign n7822 = n7850 & n7851;
  assign n7703 = n3768 & n6665;
  assign n7702 = n7730 ^ n7731;
  assign n7733 = ~n7730;
  assign n7732 = ~n7749;
  assign n7643 = n7756 ^ n7757;
  assign n7758 = ~n7757;
  assign n7736 = ~n7782;
  assign n7774 = n7783 & n210;
  assign n7775 = n7786 & n7787;
  assign n7790 = n7788 & n7764;
  assign n7795 = n7801 & n7708;
  assign n7744 = ~n7802;
  assign n7761 = n7811 & n7812;
  assign n6522 = n6525 & n6489;
  assign n7797 = n7822 ^ n5213;
  assign n7823 = ~n7822;
  assign n3672 = n7702 ^ n4881;
  assign n7676 = n7703 ^ n4936;
  assign n7722 = n7732 & n7733;
  assign n7660 = ~n7643;
  assign n7681 = n7758 & n7756;
  assign n7710 = ~n7774;
  assign n7759 = ~n7775;
  assign n7762 = ~n7790;
  assign n7712 = ~n7795;
  assign n3946 = n7796 ^ n7797;
  assign n7789 = ~n7761;
  assign n7815 = n7823 & n7824;
  assign n7641 = n7675 ^ n7676;
  assign n7677 = n7676 & n7694;
  assign n7656 = n3672 & n6646;
  assign n3674 = ~n3672;
  assign n7704 = ~n7722;
  assign n7734 = n7759 & n7760;
  assign n7745 = n7761 ^ n7762;
  assign n7750 = n3946 & n6361;
  assign n7768 = n3946 & n7777;
  assign n7776 = n7788 & n7789;
  assign n3971 = ~n3946;
  assign n7798 = ~n7815;
  assign n7620 = n7641 ^ n7642;
  assign n7633 = n7656 ^ n4879;
  assign n7657 = ~n7677;
  assign n7678 = n7704 & n7705;
  assign n7706 = n7734 ^ n7735;
  assign n7740 = n7745 & n209;
  assign n7737 = ~n7734;
  assign n7738 = ~n7745;
  assign n7649 = n7750 ^ n5213;
  assign n7765 = n3971 & n7767;
  assign n6449 = ~n7768;
  assign n7763 = ~n7776;
  assign n7769 = n7798 & n7799;
  assign n7610 = n7620 & n422;
  assign n7621 = n7633 & n7634;
  assign n7608 = ~n7620;
  assign n7622 = ~n7633;
  assign n7550 = n7657 & n7658;
  assign n7644 = n7678 ^ n4830;
  assign n7680 = n7678 & n4830;
  assign n7679 = ~n7678;
  assign n7682 = n210 ^ n7706;
  assign n7723 = n7736 & n7737;
  assign n7726 = n7738 & n7739;
  assign n7651 = ~n7740;
  assign n7727 = n7649 & n7689;
  assign n7724 = ~n7649;
  assign n7741 = n7763 & n7764;
  assign n6404 = ~n7765;
  assign n7746 = n7769 ^ n7770;
  assign n7771 = ~n7769;
  assign n7599 = n7608 & n7609;
  assign n7549 = ~n7610;
  assign n7566 = ~n7621;
  assign n7611 = n7622 & n7623;
  assign n7588 = ~n7550;
  assign n3584 = n7643 ^ n7644;
  assign n7668 = n7679 & n4834;
  assign n7659 = ~n7680;
  assign n7661 = n7681 ^ n7682;
  assign n7636 = n7682 & n7681;
  assign n7709 = ~n7723;
  assign n7715 = n7724 & n7725;
  assign n7687 = ~n7726;
  assign n7691 = ~n7727;
  assign n7707 = n7741 ^ n7742;
  assign n6446 = n6449 & n6404;
  assign n3872 = n7746 ^ n5150;
  assign n7743 = ~n7741;
  assign n7766 = n7771 & n7772;
  assign n7586 = ~n7599;
  assign n7587 = ~n7611;
  assign n7589 = n3584 & n6601;
  assign n3574 = ~n3584;
  assign n7645 = n7659 & n7660;
  assign n7647 = n7661 & n4783;
  assign n7625 = ~n7668;
  assign n7646 = ~n7661;
  assign n7695 = n7707 ^ n7708;
  assign n7670 = n7709 & n7710;
  assign n7701 = n7687 & n7651;
  assign n7653 = ~n7715;
  assign n7716 = n3872 & n7729;
  assign n7728 = n7743 & n7744;
  assign n3913 = ~n3872;
  assign n7747 = ~n7766;
  assign n7573 = n7586 & n7547;
  assign n7546 = n7586 & n7549;
  assign n7574 = n7587 & n7588;
  assign n7575 = n7587 & n7566;
  assign n7567 = n7589 ^ n4830;
  assign n7624 = ~n7645;
  assign n7635 = n7646 & n4794;
  assign n7556 = ~n7647;
  assign n7685 = n7695 & n208;
  assign n7683 = ~n7695;
  assign n7686 = ~n7670;
  assign n7671 = ~n7701;
  assign n7696 = n3913 & n6268;
  assign n6337 = ~n7716;
  assign n7713 = n3913 & n7717;
  assign n7711 = ~n7728;
  assign n7718 = n7747 & n7748;
  assign n7505 = n7546 ^ n7547;
  assign n7554 = n7567 & n7568;
  assign n7548 = ~n7573;
  assign n7565 = ~n7574;
  assign n7551 = ~n7575;
  assign n7552 = ~n7567;
  assign n7569 = n7624 & n7625;
  assign n7591 = ~n7635;
  assign n7637 = n7670 ^ n7671;
  assign n7669 = n7683 & n7684;
  assign n7580 = ~n7685;
  assign n7672 = n7686 & n7687;
  assign n7578 = n7696 ^ n5225;
  assign n7688 = n7711 & n7712;
  assign n6370 = ~n7713;
  assign n3901 = n7718 ^ n7719;
  assign n7720 = ~n7718;
  assign n5380 = n7505 ^ n5413;
  assign n7422 = n7505 & n5413;
  assign n7522 = n7548 & n7549;
  assign n7487 = n7550 ^ n7551;
  assign n7533 = n7552 & n7553;
  assign n7489 = ~n7554;
  assign n7474 = n7565 & n7566;
  assign n7590 = ~n7569;
  assign n7600 = n7591 & n7556;
  assign n7612 = n7636 ^ n7637;
  assign n7571 = n7637 & n7636;
  assign n7614 = ~n7669;
  assign n7650 = ~n7672;
  assign n7663 = n7578 & n7673;
  assign n7648 = n7688 ^ n7689;
  assign n7662 = ~n7578;
  assign n7692 = n6370 & n6337;
  assign n7690 = ~n7688;
  assign n7698 = n3901 & n6295;
  assign n3887 = ~n3901;
  assign n7714 = n7720 & n7721;
  assign n6533 = ~n5380;
  assign n7506 = n7522 & n7523;
  assign n7495 = ~n7522;
  assign n7524 = ~n7533;
  assign n7525 = ~n7474;
  assign n7576 = n7590 & n7591;
  assign n7570 = ~n7600;
  assign n7601 = n7612 & n4750;
  assign n7602 = ~n7612;
  assign n7638 = n7614 & n7580;
  assign n7499 = n7648 ^ n7649;
  assign n7603 = n7650 & n7651;
  assign n7654 = n7662 & n7616;
  assign n7582 = ~n7663;
  assign n7674 = n7690 & n7691;
  assign n6368 = ~n7692;
  assign n7664 = n3887 & n6054;
  assign n7693 = n3887 & n7697;
  assign n6256 = ~n7698;
  assign n7699 = ~n7714;
  assign n7460 = n7495 ^ n7487;
  assign n7496 = n7495 & n421;
  assign n7486 = ~n7506;
  assign n7507 = n7524 & n7525;
  assign n7508 = n7524 & n7489;
  assign n3510 = n7569 ^ n7570;
  assign n7555 = ~n7576;
  assign n7479 = ~n7601;
  assign n7592 = n7602 & n4763;
  assign n7604 = ~n7638;
  assign n7515 = ~n7499;
  assign n7613 = ~n7603;
  assign n7618 = ~n7654;
  assign n7639 = n7664 ^ n5134;
  assign n7652 = ~n7674;
  assign n6297 = ~n7693;
  assign n7665 = n7699 & n7700;
  assign n7423 = n421 ^ n7460;
  assign n7473 = n7486 & n7487;
  assign n7451 = ~n7496;
  assign n7488 = ~n7507;
  assign n7475 = ~n7508;
  assign n7509 = n7555 & n7556;
  assign n3522 = ~n3510;
  assign n7512 = ~n7592;
  assign n7572 = n7603 ^ n7604;
  assign n7605 = n7613 & n7614;
  assign n7626 = n7639 & n7640;
  assign n7615 = n7652 & n7653;
  assign n7627 = ~n7639;
  assign n7630 = n7665 ^ n5093;
  assign n7666 = ~n7665;
  assign n5341 = n7422 ^ n7423;
  assign n7321 = n7423 & n7422;
  assign n7450 = ~n7473;
  assign n7452 = n7474 ^ n7475;
  assign n7376 = n7488 & n7489;
  assign n7490 = n3522 & n6407;
  assign n7511 = ~n7509;
  assign n7557 = n7512 & n7479;
  assign n7534 = n7571 ^ n7572;
  assign n7464 = n7572 & n7571;
  assign n7579 = ~n7605;
  assign n7577 = n7615 ^ n7616;
  assign n7502 = ~n7626;
  assign n7619 = n7627 & n7628;
  assign n3852 = n7629 ^ n7630;
  assign n7617 = ~n7615;
  assign n7655 = n7666 & n7667;
  assign n6496 = ~n5341;
  assign n7363 = n7450 & n7451;
  assign n7438 = n7452 & n420;
  assign n7436 = ~n7452;
  assign n7426 = ~n7376;
  assign n7476 = n7490 ^ n4794;
  assign n7497 = n7511 & n7512;
  assign n7526 = n7534 & n4714;
  assign n7510 = ~n7557;
  assign n7527 = ~n7534;
  assign n7467 = ~n7464;
  assign n7558 = n7577 ^ n7578;
  assign n7538 = n7579 & n7580;
  assign n7594 = n3852 & n7607;
  assign n7606 = n7617 & n7618;
  assign n7544 = ~n7619;
  assign n3837 = ~n3852;
  assign n7631 = ~n7655;
  assign n7403 = ~n7363;
  assign n7424 = n7436 & n7437;
  assign n7365 = ~n7438;
  assign n7461 = n7476 & n7477;
  assign n7462 = ~n7476;
  assign n7478 = ~n7497;
  assign n3450 = n7509 ^ n7510;
  assign n7419 = ~n7526;
  assign n7513 = n7527 & n4712;
  assign n7498 = n223 ^ n7538;
  assign n7537 = n7558 & n222;
  assign n7540 = n7538 & n7559;
  assign n7535 = ~n7558;
  assign n7539 = ~n7538;
  assign n7583 = n7544 & n7502;
  assign n7560 = n3837 & n5972;
  assign n7584 = n3837 & n7593;
  assign n6186 = ~n7594;
  assign n7581 = ~n7606;
  assign n7596 = n7631 & n7632;
  assign n7402 = ~n7424;
  assign n7390 = ~n7461;
  assign n7454 = n7462 & n7463;
  assign n7456 = n7478 & n7479;
  assign n3463 = ~n3450;
  assign n7465 = n7498 ^ n7499;
  assign n7458 = ~n7513;
  assign n7528 = n7535 & n7536;
  assign n7409 = ~n7537;
  assign n7529 = n7539 & n223;
  assign n7514 = ~n7540;
  assign n7431 = n7560 ^ n5093;
  assign n7541 = n7581 & n7582;
  assign n7542 = ~n7583;
  assign n6224 = ~n7584;
  assign n3775 = n7595 ^ n7596;
  assign n7597 = ~n7596;
  assign n7388 = n7402 & n7403;
  assign n7362 = n7402 & n7365;
  assign n7425 = ~n7454;
  assign n7457 = ~n7456;
  assign n7336 = n7464 ^ n7465;
  assign n7453 = n3463 & n6424;
  assign n7455 = n7458 & n7419;
  assign n7466 = ~n7465;
  assign n7500 = n7514 & n7515;
  assign n7443 = ~n7528;
  assign n7481 = ~n7529;
  assign n7517 = n7431 & n7530;
  assign n7341 = n7541 ^ n7542;
  assign n7516 = ~n7431;
  assign n6221 = n6224 & n6186;
  assign n7543 = ~n7541;
  assign n7532 = n3775 & n6024;
  assign n7561 = n3775 & n6147;
  assign n3665 = ~n3775;
  assign n7585 = n7597 & n7598;
  assign n7322 = n7362 ^ n7363;
  assign n7364 = ~n7388;
  assign n7414 = n7425 & n7426;
  assign n7417 = n7425 & n7390;
  assign n7429 = n7336 & n4671;
  assign n7309 = n7453 ^ n4763;
  assign n3410 = n7455 ^ n7456;
  assign n7439 = n7457 & n7458;
  assign n7428 = ~n7336;
  assign n7405 = n7466 & n7467;
  assign n7440 = n7443 & n7409;
  assign n7480 = ~n7500;
  assign n7503 = n7516 & n7469;
  assign n7434 = ~n7517;
  assign n7397 = n7532 ^ n5046;
  assign n7531 = n7543 & n7544;
  assign n6149 = ~n7561;
  assign n7545 = n3665 & n7562;
  assign n7563 = ~n7585;
  assign n5327 = n7321 ^ n7322;
  assign n7323 = ~n7322;
  assign n7248 = n7364 & n7365;
  assign n7389 = ~n7414;
  assign n7377 = ~n7417;
  assign n7415 = n7309 & n7427;
  assign n7391 = n3410 & n6250;
  assign n7420 = n7428 & n4673;
  assign n7379 = ~n7429;
  assign n7416 = ~n7309;
  assign n3401 = ~n3410;
  assign n7418 = ~n7439;
  assign n7441 = n7480 & n7481;
  assign n7471 = ~n7503;
  assign n7493 = n7397 & n7357;
  assign n7491 = ~n7397;
  assign n7501 = ~n7531;
  assign n6109 = ~n7545;
  assign n7518 = n7563 & n7564;
  assign n6402 = ~n5327;
  assign n7212 = n7323 & n7321;
  assign n7297 = ~n7248;
  assign n7353 = n7376 ^ n7377;
  assign n7346 = n7389 & n7390;
  assign n7366 = n7391 ^ n4712;
  assign n7312 = ~n7415;
  assign n7404 = n7416 & n7347;
  assign n7378 = n7418 & n7419;
  assign n7339 = ~n7420;
  assign n7406 = n7440 ^ n7441;
  assign n7442 = ~n7441;
  assign n7482 = n7491 & n7492;
  assign n7360 = ~n7493;
  assign n7468 = n7501 & n7502;
  assign n3639 = n7518 ^ n7519;
  assign n7520 = ~n7518;
  assign n7310 = n7346 ^ n7347;
  assign n7335 = n7353 & n419;
  assign n7350 = n7366 & n7367;
  assign n7332 = ~n7353;
  assign n7348 = ~n7346;
  assign n7351 = ~n7366;
  assign n7337 = n7378 ^ n4671;
  assign n7349 = ~n7404;
  assign n7380 = ~n7378;
  assign n7392 = n7405 ^ n7406;
  assign n7303 = n7406 & n7405;
  assign n7432 = n7442 & n7443;
  assign n7430 = n7468 ^ n7469;
  assign n7399 = ~n7482;
  assign n7470 = ~n7468;
  assign n7483 = n3639 & n7494;
  assign n3637 = ~n3639;
  assign n7504 = n7520 & n7521;
  assign n7284 = n7309 ^ n7310;
  assign n7324 = n7332 & n7333;
  assign n7261 = ~n7335;
  assign n3353 = n7336 ^ n7337;
  assign n7331 = n7348 & n7349;
  assign n7238 = ~n7350;
  assign n7334 = n7351 & n7352;
  assign n7368 = n7379 & n7380;
  assign n7382 = n7392 & n4649;
  assign n7381 = ~n7392;
  assign n7306 = ~n7303;
  assign n7407 = n7430 ^ n7431;
  assign n7408 = ~n7432;
  assign n7459 = n7470 & n7471;
  assign n7444 = n3637 & n5905;
  assign n7472 = n3637 & n6072;
  assign n6039 = ~n7483;
  assign n7484 = ~n7504;
  assign n7274 = n7284 & n418;
  assign n7272 = ~n7284;
  assign n7275 = n3353 & n6181;
  assign n7296 = ~n7324;
  assign n3369 = ~n3353;
  assign n7311 = ~n7331;
  assign n7277 = ~n7334;
  assign n7338 = ~n7368;
  assign n7369 = n7381 & n4626;
  assign n7301 = ~n7382;
  assign n7395 = n7407 & n220;
  assign n7370 = n7408 & n7409;
  assign n7393 = ~n7407;
  assign n7317 = n7444 ^ n5050;
  assign n7433 = ~n7459;
  assign n6074 = ~n7472;
  assign n7445 = n7484 & n7485;
  assign n7259 = n7272 & n7273;
  assign n7190 = ~n7274;
  assign n7246 = n7275 ^ n4671;
  assign n7285 = n7296 & n7297;
  assign n7286 = n7296 & n7261;
  assign n7262 = n7311 & n7312;
  assign n7298 = n7277 & n7238;
  assign n7300 = n7338 & n7339;
  assign n7266 = ~n7369;
  assign n7340 = n221 ^ n7370;
  assign n7372 = n7370 & n7384;
  assign n7383 = n7393 & n7394;
  assign n7243 = ~n7395;
  assign n7371 = ~n7370;
  assign n7410 = n7317 & n7421;
  assign n7396 = n7433 & n7434;
  assign n7411 = ~n7317;
  assign n7412 = n7445 ^ n7446;
  assign n7449 = n7445 & n7446;
  assign n7447 = ~n7445;
  assign n7233 = n7246 & n7247;
  assign n7223 = ~n7259;
  assign n7234 = ~n7246;
  assign n7260 = ~n7285;
  assign n7249 = ~n7286;
  assign n7276 = ~n7262;
  assign n7263 = ~n7298;
  assign n7302 = ~n7300;
  assign n7299 = n7266 & n7301;
  assign n7304 = n7340 ^ n7341;
  assign n7358 = n7371 & n221;
  assign n7354 = ~n7372;
  assign n7282 = ~n7383;
  assign n7356 = n7396 ^ n7397;
  assign n7319 = ~n7410;
  assign n7400 = n7411 & n7289;
  assign n3557 = n7412 ^ n4985;
  assign n7398 = ~n7396;
  assign n7435 = n7447 & n7448;
  assign n7375 = ~n7449;
  assign n7225 = n7223 & n7190;
  assign n7174 = ~n7233;
  assign n7228 = n7234 & n7235;
  assign n7213 = n7248 ^ n7249;
  assign n7187 = n7260 & n7261;
  assign n7236 = n7262 ^ n7263;
  assign n7264 = n7276 & n7277;
  assign n3318 = n7299 ^ n7300;
  assign n7287 = n7301 & n7302;
  assign n7278 = n7303 ^ n7304;
  assign n7305 = ~n7304;
  assign n7343 = n7354 & n7341;
  assign n7176 = n7356 ^ n7357;
  assign n7314 = ~n7358;
  assign n7355 = n7282 & n7243;
  assign n7385 = n7398 & n7399;
  assign n7291 = ~n7400;
  assign n3569 = ~n3557;
  assign n7413 = n7375 & n4985;
  assign n7387 = ~n7435;
  assign n5291 = n7212 ^ n7213;
  assign n7188 = ~n7225;
  assign n7198 = ~n7228;
  assign n7159 = n7213 & n7212;
  assign n7229 = n7236 & n417;
  assign n7224 = ~n7187;
  assign n7226 = ~n7236;
  assign n7237 = ~n7264;
  assign n7239 = n3318 & n6120;
  assign n7267 = n7278 & n4613;
  assign n3321 = ~n3318;
  assign n7265 = ~n7287;
  assign n7268 = ~n7278;
  assign n7240 = n7305 & n7306;
  assign n7325 = n7176 & n7342;
  assign n7313 = ~n7343;
  assign n7326 = ~n7176;
  assign n7280 = ~n7355;
  assign n7327 = n3569 & n5738;
  assign n7359 = ~n7385;
  assign n7401 = n7387 & n4983;
  assign n7386 = ~n7413;
  assign n7160 = n7187 ^ n7188;
  assign n7171 = n7198 & n7174;
  assign n6334 = ~n5291;
  assign n7162 = ~n7159;
  assign n7211 = n7223 & n7224;
  assign n7214 = n7226 & n7227;
  assign n7140 = ~n7229;
  assign n7172 = n7237 & n7238;
  assign n7215 = n7239 ^ n4649;
  assign n7182 = n7265 & n7266;
  assign n7194 = ~n7267;
  assign n7250 = n7268 & n4589;
  assign n7279 = n7313 & n7314;
  assign n7207 = ~n7325;
  assign n7315 = n7326 & n219;
  assign n7220 = n7327 ^ n4983;
  assign n7316 = n7359 & n7360;
  assign n7373 = n7386 & n7387;
  assign n7374 = ~n7401;
  assign n5230 = n7159 ^ n7160;
  assign n7089 = n7171 ^ n7172;
  assign n7161 = ~n7160;
  assign n7189 = ~n7211;
  assign n7166 = ~n7214;
  assign n7200 = n7215 & n7216;
  assign n7199 = ~n7172;
  assign n7201 = ~n7215;
  assign n7230 = ~n7182;
  assign n7231 = ~n7250;
  assign n7241 = n7279 ^ n7280;
  assign n7281 = ~n7279;
  assign n7293 = n7220 & n7307;
  assign n7178 = ~n7315;
  assign n7288 = n7316 ^ n7317;
  assign n7292 = ~n7220;
  assign n7318 = ~n7316;
  assign n7344 = ~n7373;
  assign n7361 = n7374 & n7375;
  assign n6219 = ~n5230;
  assign n7135 = n7161 & n7162;
  assign n7097 = ~n7089;
  assign n7164 = n7189 & n7190;
  assign n7163 = n7166 & n7140;
  assign n7191 = n7198 & n7199;
  assign n7124 = ~n7200;
  assign n7192 = n7201 & n7202;
  assign n7217 = n7230 & n7231;
  assign n7218 = n7231 & n7194;
  assign n7144 = n7240 ^ n7241;
  assign n7151 = n7241 & n7240;
  assign n7270 = n7281 & n7282;
  assign n7269 = n7288 ^ n7289;
  assign n7283 = n7292 & n7255;
  assign n7222 = ~n7293;
  assign n7308 = n7318 & n7319;
  assign n7328 = n7344 & n7345;
  assign n7329 = ~n7361;
  assign n7138 = ~n7135;
  assign n7136 = n7163 ^ n7164;
  assign n7165 = ~n7164;
  assign n7173 = ~n7191;
  assign n7149 = ~n7192;
  assign n7193 = ~n7217;
  assign n7183 = ~n7218;
  assign n7204 = n7144 & n4582;
  assign n7203 = ~n7144;
  assign n7253 = n7269 & n218;
  assign n7242 = ~n7270;
  assign n7251 = ~n7269;
  assign n7257 = ~n7283;
  assign n7290 = ~n7308;
  assign n7295 = ~n7328;
  assign n7320 = n7329 & n7330;
  assign n5193 = n7135 ^ n7136;
  assign n7137 = ~n7136;
  assign n7157 = n7165 & n7166;
  assign n7141 = n7173 & n7174;
  assign n7167 = n7124 & n7149;
  assign n3278 = n7182 ^ n7183;
  assign n7168 = n7193 & n7194;
  assign n7195 = n7203 & n4550;
  assign n7147 = ~n7204;
  assign n7205 = n7242 & n7243;
  assign n7244 = n7251 & n7252;
  assign n7132 = ~n7253;
  assign n7254 = n7290 & n7291;
  assign n7294 = ~n7320;
  assign n6194 = ~n5193;
  assign n7061 = n7137 & n7138;
  assign n7139 = ~n7157;
  assign n7150 = ~n7141;
  assign n7142 = ~n7167;
  assign n7145 = n7168 ^ n4550;
  assign n3286 = ~n3278;
  assign n7169 = ~n7168;
  assign n7170 = ~n7195;
  assign n7175 = n219 ^ n7205;
  assign n7206 = ~n7205;
  assign n7156 = ~n7244;
  assign n7219 = n7254 ^ n7255;
  assign n7256 = ~n7254;
  assign n3484 = n7294 & n7295;
  assign n7064 = ~n7061;
  assign n7114 = n7139 & n7140;
  assign n7030 = n7141 ^ n7142;
  assign n3223 = n7144 ^ n7145;
  assign n7143 = n7149 & n7150;
  assign n7133 = n3286 & n6076;
  assign n7158 = n7169 & n7170;
  assign n7152 = n7175 ^ n7176;
  assign n7197 = n7206 & n7207;
  assign n7208 = n7156 & n7132;
  assign n7196 = n7219 ^ n7220;
  assign n7245 = n7256 & n7257;
  assign n5864 = n7258 ^ n3484;
  assign n7232 = n3484 & n7271;
  assign n5016 = ~n3484;
  assign n7088 = n416 ^ n7114;
  assign n7118 = n7114 & n7122;
  assign n7119 = n7030 & n431;
  assign n7115 = ~n7114;
  assign n7116 = ~n7030;
  assign n3258 = ~n3223;
  assign n7072 = n7133 ^ n4589;
  assign n7123 = ~n7143;
  assign n7134 = n7151 ^ n7152;
  assign n7146 = ~n7158;
  assign n7127 = n7152 & n7151;
  assign n7186 = n7196 & n217;
  assign n7177 = ~n7197;
  assign n7154 = ~n7208;
  assign n7184 = ~n7196;
  assign n7210 = n7232 ^ n4926;
  assign n7221 = ~n7245;
  assign n5875 = ~n5864;
  assign n7062 = n7088 ^ n7089;
  assign n7109 = n7115 & n416;
  assign n7110 = n7116 & n7117;
  assign n7096 = ~n7118;
  assign n7032 = ~n7119;
  assign n7112 = n7072 & n7120;
  assign n7091 = n3258 & n5894;
  assign n7098 = n7123 & n7124;
  assign n7111 = ~n7072;
  assign n7125 = n7134 & n4536;
  assign n7068 = n7146 & n7147;
  assign n7126 = ~n7134;
  assign n7130 = ~n7127;
  assign n7153 = n7177 & n7178;
  assign n7179 = n7184 & n7185;
  assign n7085 = ~n7186;
  assign n7181 = n7209 ^ n7210;
  assign n7180 = n7221 & n7222;
  assign n6080 = n7061 ^ n7062;
  assign n7063 = ~n7062;
  assign n7075 = n7091 ^ n4550;
  assign n7090 = n7096 & n7097;
  assign n7071 = n7098 ^ n7099;
  assign n7074 = ~n7109;
  assign n7050 = ~n7110;
  assign n7100 = n7111 & n7099;
  assign n7058 = ~n7112;
  assign n7086 = ~n7098;
  assign n7079 = ~n7125;
  assign n7121 = n7126 & n4509;
  assign n7101 = ~n7068;
  assign n7128 = n7153 ^ n7154;
  assign n7155 = ~n7153;
  assign n7108 = ~n7179;
  assign n7037 = n7180 ^ n7181;
  assign n5153 = ~n6080;
  assign n7010 = n7063 & n7064;
  assign n6992 = n7071 ^ n7072;
  assign n7065 = n7075 & n7076;
  assign n7066 = ~n7075;
  assign n7073 = ~n7090;
  assign n7087 = ~n7100;
  assign n7102 = ~n7121;
  assign n7113 = n7127 ^ n7128;
  assign n7129 = ~n7128;
  assign n7148 = n7155 & n7156;
  assign n7105 = n7108 & n7085;
  assign n7048 = n6992 & n430;
  assign n7046 = ~n6992;
  assign n7025 = ~n7065;
  assign n7059 = n7066 & n7067;
  assign n7049 = n7073 & n7074;
  assign n7077 = n7086 & n7087;
  assign n7092 = n7101 & n7102;
  assign n7093 = n7102 & n7079;
  assign n7103 = n7113 & n4495;
  assign n7104 = ~n7113;
  assign n7080 = n7129 & n7130;
  assign n7131 = ~n7148;
  assign n7040 = n7046 & n7047;
  assign n6994 = ~n7048;
  assign n7029 = n431 ^ n7049;
  assign n7038 = ~n7059;
  assign n7051 = ~n7049;
  assign n7057 = ~n7077;
  assign n7078 = ~n7092;
  assign n7069 = ~n7093;
  assign n7052 = ~n7103;
  assign n7094 = n7104 & n4466;
  assign n7083 = ~n7080;
  assign n7106 = n7131 & n7132;
  assign n7011 = n7029 ^ n7030;
  assign n7013 = ~n7040;
  assign n7026 = n7025 & n7038;
  assign n7041 = n7050 & n7051;
  assign n7027 = n7057 & n7058;
  assign n3171 = n7068 ^ n7069;
  assign n7042 = n7078 & n7079;
  assign n7035 = ~n7094;
  assign n7081 = n7105 ^ n7106;
  assign n7107 = ~n7106;
  assign n5117 = n7010 ^ n7011;
  assign n6972 = n7011 & n7010;
  assign n6955 = n7026 ^ n7027;
  assign n7031 = ~n7041;
  assign n7039 = ~n7027;
  assign n3218 = ~n3171;
  assign n7053 = ~n7042;
  assign n7070 = n7035 & n7052;
  assign n7060 = n7080 ^ n7081;
  assign n7082 = ~n7081;
  assign n7095 = n7107 & n7108;
  assign n6003 = ~n5117;
  assign n6975 = ~n6972;
  assign n7003 = n6955 & n7015;
  assign n7004 = ~n6955;
  assign n7012 = n7031 & n7032;
  assign n7033 = n7038 & n7039;
  assign n7028 = n3218 & n5879;
  assign n7044 = n7052 & n7053;
  assign n7054 = n7060 & n4469;
  assign n7043 = ~n7070;
  assign n7055 = ~n7060;
  assign n7022 = n7082 & n7083;
  assign n7084 = ~n7095;
  assign n6977 = ~n7003;
  assign n7000 = n7004 & n429;
  assign n6991 = n430 ^ n7012;
  assign n7014 = ~n7012;
  assign n7016 = n7028 ^ n4509;
  assign n7024 = ~n7033;
  assign n3152 = n7042 ^ n7043;
  assign n7034 = ~n7044;
  assign n6997 = ~n7054;
  assign n7045 = n7055 & n4424;
  assign n7056 = n7084 & n7085;
  assign n6973 = n6991 ^ n6992;
  assign n6957 = ~n7000;
  assign n7002 = n7013 & n7014;
  assign n7005 = n7016 & n7017;
  assign n6965 = n7024 & n7025;
  assign n7006 = ~n7016;
  assign n7019 = n7034 & n7035;
  assign n3160 = ~n3152;
  assign n7021 = ~n7045;
  assign n7036 = n216 ^ n7056;
  assign n5073 = n6972 ^ n6973;
  assign n6974 = ~n6973;
  assign n6993 = ~n7002;
  assign n6970 = ~n7005;
  assign n7001 = n7006 & n7007;
  assign n6986 = ~n6965;
  assign n7008 = n3160 & n5829;
  assign n7020 = ~n7019;
  assign n7018 = n7021 & n6997;
  assign n7023 = n7036 ^ n7037;
  assign n5906 = ~n5073;
  assign n5794 = n6974 & n6975;
  assign n6976 = n6993 & n6994;
  assign n6987 = ~n7001;
  assign n6935 = n7008 ^ n4495;
  assign n3094 = n7018 ^ n7019;
  assign n7009 = n7020 & n7021;
  assign n6960 = n7022 ^ n7023;
  assign n6954 = n429 ^ n6976;
  assign n6978 = ~n6976;
  assign n6983 = n6986 & n6987;
  assign n6984 = n6987 & n6970;
  assign n6989 = n6935 & n6995;
  assign n6982 = n3094 & n5675;
  assign n6988 = ~n6935;
  assign n6999 = n6960 & n4416;
  assign n3096 = ~n3094;
  assign n6996 = ~n7009;
  assign n6998 = ~n6960;
  assign n5755 = n6954 ^ n6955;
  assign n6967 = n6977 & n6978;
  assign n6900 = n6982 ^ n4424;
  assign n6969 = ~n6983;
  assign n6966 = ~n6984;
  assign n6985 = n6988 & n6951;
  assign n6938 = ~n6989;
  assign n6979 = n6996 & n6997;
  assign n6990 = n6998 & n4379;
  assign n6962 = ~n6999;
  assign n6891 = n5755 & n5794;
  assign n6949 = n6965 ^ n6966;
  assign n6956 = ~n6967;
  assign n6964 = n6900 & n6968;
  assign n6950 = n6969 & n6970;
  assign n6963 = ~n6900;
  assign n6959 = n6979 ^ n4416;
  assign n6952 = ~n6985;
  assign n6980 = ~n6979;
  assign n6981 = ~n6990;
  assign n6947 = n6949 & n428;
  assign n6936 = n6950 ^ n6951;
  assign n6917 = n6956 & n6957;
  assign n3106 = n6959 ^ n6960;
  assign n6945 = ~n6949;
  assign n6958 = n6963 & n6925;
  assign n6902 = ~n6964;
  assign n6953 = ~n6950;
  assign n6971 = n6980 & n6981;
  assign n6928 = n6935 ^ n6936;
  assign n6940 = n6945 & n6946;
  assign n6911 = ~n6947;
  assign n6934 = n3106 & n5651;
  assign n6932 = ~n6917;
  assign n6948 = n6952 & n6953;
  assign n3100 = ~n3106;
  assign n6927 = ~n6958;
  assign n6961 = ~n6971;
  assign n6923 = n6928 & n427;
  assign n6919 = ~n6928;
  assign n6921 = n6934 ^ n4379;
  assign n6933 = ~n6940;
  assign n6937 = ~n6948;
  assign n6941 = n6961 & n6962;
  assign n6912 = n6919 & n6920;
  assign n6913 = n6921 & n6922;
  assign n6873 = ~n6923;
  assign n6914 = ~n6921;
  assign n6929 = n6932 & n6933;
  assign n6916 = n6933 & n6911;
  assign n6924 = n6937 & n6938;
  assign n3078 = n6941 ^ n6942;
  assign n6943 = ~n6941;
  assign n6894 = ~n6912;
  assign n6860 = ~n6913;
  assign n6904 = n6914 & n6915;
  assign n6892 = n6916 ^ n6917;
  assign n6899 = n6924 ^ n6925;
  assign n6910 = ~n6929;
  assign n6926 = ~n6924;
  assign n3085 = ~n3078;
  assign n6939 = n6943 & n6944;
  assign n3752 = n6891 ^ n6892;
  assign n6896 = n6894 & n6873;
  assign n6883 = n6899 ^ n6900;
  assign n6880 = ~n6904;
  assign n6893 = ~n6892;
  assign n6870 = n6910 & n6911;
  assign n6918 = n6926 & n6927;
  assign n6905 = n3085 & n5634;
  assign n6930 = ~n6939;
  assign n4971 = n3752 ^ n6803;
  assign n3754 = ~n3752;
  assign n6879 = n6883 & n426;
  assign n6850 = n6893 & n6891;
  assign n6885 = n6860 & n6880;
  assign n6871 = ~n6896;
  assign n6877 = ~n6883;
  assign n6895 = ~n6870;
  assign n6897 = n6905 ^ n4337;
  assign n6901 = ~n6918;
  assign n6907 = n6930 & n6931;
  assign n2728 = n4971 ^ n4953;
  assign n6776 = n3754 & n3807;
  assign n6851 = n6870 ^ n6871;
  assign n6874 = n6877 & n6878;
  assign n6833 = ~n6879;
  assign n6853 = ~n6850;
  assign n6865 = ~n6885;
  assign n6884 = n6894 & n6895;
  assign n6886 = n6897 & n6898;
  assign n6864 = n6901 & n6902;
  assign n6887 = ~n6897;
  assign n2955 = n6906 ^ n6907;
  assign n6908 = ~n6907;
  assign n4970 = ~n2728;
  assign n6835 = n6850 ^ n6851;
  assign n6854 = n6864 ^ n6865;
  assign n6852 = ~n6851;
  assign n6855 = ~n6874;
  assign n6872 = ~n6884;
  assign n6819 = ~n6886;
  assign n6882 = n6887 & n6888;
  assign n6881 = ~n6864;
  assign n6876 = n2955 & n5547;
  assign n3013 = ~n2955;
  assign n6903 = n6908 & n6909;
  assign n6821 = n4970 & n6829;
  assign n6822 = n4970 & n4953;
  assign n6830 = n6835 & n3768;
  assign n6831 = ~n6835;
  assign n6810 = n6852 & n6853;
  assign n6845 = n6854 & n425;
  assign n6836 = n6855 & n6833;
  assign n6843 = ~n6854;
  assign n6837 = n6872 & n6873;
  assign n6765 = n6876 ^ n4298;
  assign n6875 = n6880 & n6881;
  assign n6842 = ~n6882;
  assign n6889 = ~n6903;
  assign n6774 = ~n6821;
  assign n6802 = ~n6822;
  assign n6805 = ~n6830;
  assign n6823 = n6831 & n3710;
  assign n6811 = n6836 ^ n6837;
  assign n6813 = ~n6810;
  assign n6838 = n6843 & n6844;
  assign n6779 = ~n6845;
  assign n6858 = n6765 & n6861;
  assign n6856 = ~n6837;
  assign n6862 = n6819 & n6842;
  assign n6857 = ~n6765;
  assign n6859 = ~n6875;
  assign n6866 = n6889 & n6890;
  assign n6793 = n6802 & n6803;
  assign n6804 = n6805 & n6776;
  assign n6794 = n6810 ^ n6811;
  assign n6783 = ~n6823;
  assign n6812 = ~n6811;
  assign n6807 = ~n6838;
  assign n6846 = n6855 & n6856;
  assign n6847 = n6857 & n6789;
  assign n6767 = ~n6858;
  assign n6839 = n6859 & n6860;
  assign n6840 = ~n6862;
  assign n2992 = n6866 ^ n6867;
  assign n6868 = ~n6866;
  assign n6773 = ~n6793;
  assign n6784 = n6794 & n3674;
  assign n6782 = ~n6804;
  assign n6775 = n6783 & n6805;
  assign n6785 = ~n6794;
  assign n6762 = n6812 & n6813;
  assign n6816 = n6807 & n6779;
  assign n6824 = n6839 ^ n6840;
  assign n6832 = ~n6846;
  assign n6791 = ~n6847;
  assign n6841 = ~n6839;
  assign n3001 = ~n2992;
  assign n6863 = n6868 & n6869;
  assign n6750 = n6773 & n6774;
  assign n2695 = n6775 ^ n6776;
  assign n6722 = n6782 & n6783;
  assign n6737 = ~n6784;
  assign n6777 = n6785 & n3672;
  assign n6787 = ~n6816;
  assign n6817 = n6824 & n424;
  assign n6786 = n6832 & n6833;
  assign n6814 = ~n6824;
  assign n6834 = n6841 & n6842;
  assign n6825 = n3001 & n5484;
  assign n6848 = ~n6863;
  assign n6734 = n6750 ^ n6751;
  assign n6720 = n6750 ^ n6752;
  assign n2697 = ~n2695;
  assign n6760 = ~n6722;
  assign n6761 = ~n6777;
  assign n6763 = n6786 ^ n6787;
  assign n6808 = n6814 & n6815;
  assign n6728 = ~n6817;
  assign n6806 = ~n6786;
  assign n6743 = n6825 ^ n4235;
  assign n6818 = ~n6834;
  assign n6826 = n6848 & n6849;
  assign n4771 = n135 ^ n6720;
  assign n6692 = n6734 & n6735;
  assign n6560 = n6720 & n135;
  assign n6721 = n2697 & n4934;
  assign n6753 = n6760 & n6761;
  assign n6754 = n6761 & n6737;
  assign n6746 = n6762 ^ n6763;
  assign n6725 = n6763 & n6762;
  assign n6795 = n6806 & n6807;
  assign n6758 = ~n6808;
  assign n6797 = n6743 & n6809;
  assign n6788 = n6818 & n6819;
  assign n6796 = ~n6743;
  assign n6798 = n6826 ^ n4249;
  assign n6827 = ~n6826;
  assign n6703 = n6692 & n6665;
  assign n6414 = ~n4771;
  assign n6701 = ~n6692;
  assign n6672 = n6721 ^ n3768;
  assign n6739 = n6746 & n3574;
  assign n6736 = ~n6753;
  assign n6723 = ~n6754;
  assign n6738 = ~n6746;
  assign n6780 = n6758 & n6728;
  assign n6764 = n6788 ^ n6789;
  assign n6778 = ~n6795;
  assign n6792 = n6796 & n6707;
  assign n6745 = ~n6797;
  assign n2873 = n6798 ^ n6799;
  assign n6790 = ~n6788;
  assign n6820 = n6827 & n6828;
  assign n6664 = n6692 ^ n6672;
  assign n6693 = n6701 & n6702;
  assign n6644 = ~n6703;
  assign n2536 = n6722 ^ n6723;
  assign n6674 = n6736 & n6737;
  assign n6724 = n6738 & n3584;
  assign n6676 = ~n6739;
  assign n6681 = n6764 ^ n6765;
  assign n6755 = n6778 & n6779;
  assign n6756 = ~n6780;
  assign n6759 = n2873 & n5508;
  assign n6781 = n6790 & n6791;
  assign n6711 = ~n6792;
  assign n2932 = ~n2873;
  assign n6800 = ~n6820;
  assign n6642 = n6664 ^ n6665;
  assign n6671 = ~n6693;
  assign n2529 = ~n2536;
  assign n6704 = ~n6674;
  assign n6705 = ~n6724;
  assign n6726 = n6755 ^ n6756;
  assign n6740 = n6759 ^ n4198;
  assign n6757 = ~n6755;
  assign n6766 = ~n6781;
  assign n6770 = n6800 & n6801;
  assign n6634 = n6642 & n134;
  assign n6632 = ~n6642;
  assign n6666 = n6671 & n6672;
  assign n6667 = n2529 & n4881;
  assign n6694 = n6704 & n6705;
  assign n6673 = n6705 & n6676;
  assign n6606 = n6725 ^ n6726;
  assign n6622 = n6726 & n6725;
  assign n6729 = n6740 & n6741;
  assign n6730 = ~n6740;
  assign n6747 = n6757 & n6758;
  assign n6742 = n6766 & n6767;
  assign n2829 = n6769 ^ n6770;
  assign n6771 = ~n6770;
  assign n6619 = n6632 & n6633;
  assign n6562 = ~n6634;
  assign n6643 = ~n6666;
  assign n6645 = n6667 ^ n3672;
  assign n2410 = n6673 ^ n6674;
  assign n6675 = ~n6694;
  assign n6695 = n6606 & n3510;
  assign n6696 = ~n6606;
  assign n6653 = ~n6729;
  assign n6715 = n6730 & n6731;
  assign n6706 = n6742 ^ n6743;
  assign n6727 = ~n6747;
  assign n6744 = ~n6742;
  assign n6733 = n2829 & n5426;
  assign n2879 = ~n2829;
  assign n6768 = n6771 & n6772;
  assign n6597 = ~n6619;
  assign n6548 = n6643 & n6644;
  assign n6637 = n6645 & n6646;
  assign n6620 = n2410 & n4834;
  assign n6635 = ~n6645;
  assign n2472 = ~n2410;
  assign n6647 = n6675 & n6676;
  assign n6608 = ~n6695;
  assign n6684 = n6696 & n3522;
  assign n6685 = n6706 ^ n6707;
  assign n6682 = ~n6715;
  assign n6708 = n6727 & n6728;
  assign n6712 = n6733 ^ n4156;
  assign n6732 = n6744 & n6745;
  assign n6748 = ~n6768;
  assign n6584 = n6597 & n6560;
  assign n6559 = n6597 & n6562;
  assign n6600 = n6620 ^ n3584;
  assign n6598 = ~n6548;
  assign n6621 = n6635 & n6636;
  assign n6564 = ~n6637;
  assign n6605 = n6647 ^ n3522;
  assign n6648 = ~n6647;
  assign n6649 = ~n6684;
  assign n6679 = n6685 & n438;
  assign n6677 = ~n6685;
  assign n6688 = n6653 & n6682;
  assign n6697 = n6708 & n6709;
  assign n6698 = n6712 & n6713;
  assign n6686 = ~n6708;
  assign n6699 = ~n6712;
  assign n6710 = ~n6732;
  assign n6716 = n6748 & n6749;
  assign n4721 = n6559 ^ n6560;
  assign n6561 = ~n6584;
  assign n6586 = n6600 & n6601;
  assign n2365 = n6605 ^ n6606;
  assign n6587 = ~n6600;
  assign n6599 = ~n6621;
  assign n6638 = n6648 & n6649;
  assign n6668 = n6677 & n6678;
  assign n6575 = ~n6679;
  assign n6655 = n6686 ^ n6681;
  assign n6657 = ~n6688;
  assign n6687 = n6686 & n439;
  assign n6680 = ~n6697;
  assign n6581 = ~n6698;
  assign n6689 = n6699 & n6700;
  assign n6656 = n6710 & n6711;
  assign n2850 = n6716 ^ n6717;
  assign n6718 = ~n6716;
  assign n4748 = ~n4721;
  assign n6534 = n6561 & n6562;
  assign n6492 = ~n6586;
  assign n6569 = n6587 & n6588;
  assign n6585 = n6598 & n6599;
  assign n6589 = n6564 & n6599;
  assign n2355 = ~n2365;
  assign n6607 = ~n6638;
  assign n6623 = n439 ^ n6655;
  assign n6639 = n6656 ^ n6657;
  assign n6612 = ~n6668;
  assign n6669 = n6680 & n6681;
  assign n6651 = ~n6687;
  assign n6617 = ~n6689;
  assign n6683 = ~n6656;
  assign n2860 = ~n2850;
  assign n6714 = n6718 & n6719;
  assign n6526 = n6534 & n6535;
  assign n6515 = ~n6534;
  assign n6528 = ~n6569;
  assign n6536 = n2355 & n4783;
  assign n6563 = ~n6585;
  assign n6549 = ~n6589;
  assign n6602 = n6607 & n6608;
  assign n6565 = n6622 ^ n6623;
  assign n6570 = n6623 & n6622;
  assign n6626 = n6639 & n437;
  assign n6609 = n6612 & n6575;
  assign n6624 = ~n6639;
  assign n6650 = ~n6669;
  assign n6658 = n6617 & n6581;
  assign n6670 = n6682 & n6683;
  assign n6659 = n2860 & n5412;
  assign n6690 = ~n6714;
  assign n6516 = n6515 & n133;
  assign n6497 = ~n6526;
  assign n6451 = n6536 ^ n3510;
  assign n6537 = n6528 & n6492;
  assign n6498 = n6548 ^ n6549;
  assign n6501 = n6563 & n6564;
  assign n6591 = n6565 & n3450;
  assign n6550 = ~n6602;
  assign n6590 = ~n6565;
  assign n6613 = n6624 & n6625;
  assign n6506 = ~n6626;
  assign n6610 = n6650 & n6651;
  assign n6615 = ~n6658;
  assign n6640 = n6659 ^ n4111;
  assign n6652 = ~n6670;
  assign n6660 = n6690 & n6691;
  assign n6490 = n6497 & n6498;
  assign n6482 = n6515 ^ n6498;
  assign n6465 = ~n6516;
  assign n6499 = n6451 & n6517;
  assign n6500 = ~n6451;
  assign n6502 = ~n6537;
  assign n6527 = ~n6501;
  assign n6529 = n6550 ^ n6565;
  assign n6573 = n6590 & n3463;
  assign n6520 = ~n6591;
  assign n6571 = n6609 ^ n6610;
  assign n6542 = ~n6613;
  assign n6611 = ~n6610;
  assign n6627 = n6640 & n6641;
  assign n6614 = n6652 & n6653;
  assign n6628 = ~n6640;
  assign n2709 = n6660 ^ n6661;
  assign n6662 = ~n6660;
  assign n6439 = n133 ^ n6482;
  assign n6464 = ~n6490;
  assign n6452 = ~n6499;
  assign n6493 = n6500 & n6407;
  assign n6483 = n6501 ^ n6502;
  assign n6518 = n6527 & n6528;
  assign n2295 = n3450 ^ n6529;
  assign n6441 = n6570 ^ n6571;
  assign n6551 = ~n6573;
  assign n6578 = n6542 & n6506;
  assign n6572 = ~n6571;
  assign n6603 = n6611 & n6612;
  assign n6592 = n6614 ^ n6615;
  assign n6511 = ~n6627;
  assign n6618 = n6628 & n6629;
  assign n6616 = ~n6614;
  assign n2807 = ~n2709;
  assign n6654 = n6662 & n6663;
  assign n4699 = n6439 ^ n4721;
  assign n6338 = n6439 & n4721;
  assign n6374 = n6464 & n6465;
  assign n6468 = n6483 & n132;
  assign n6409 = ~n6493;
  assign n6466 = ~n6483;
  assign n6491 = ~n6518;
  assign n2188 = ~n2295;
  assign n6538 = n6550 & n6551;
  assign n6457 = ~n6441;
  assign n6503 = n6572 & n6570;
  assign n6540 = ~n6578;
  assign n6579 = n6592 & n436;
  assign n6574 = ~n6603;
  assign n6576 = ~n6592;
  assign n6604 = n6616 & n6617;
  assign n6546 = ~n6618;
  assign n6593 = n2807 & n5350;
  assign n6630 = ~n6654;
  assign n6237 = ~n4699;
  assign n6421 = ~n6374;
  assign n6454 = n6466 & n6467;
  assign n6387 = ~n6468;
  assign n6450 = n6491 & n6492;
  assign n6455 = n2188 & n4750;
  assign n6519 = ~n6538;
  assign n6539 = n6574 & n6575;
  assign n6566 = n6576 & n6577;
  assign n6430 = ~n6579;
  assign n6582 = n6546 & n6511;
  assign n6567 = n6593 ^ n4070;
  assign n6580 = ~n6604;
  assign n6594 = n6630 & n6631;
  assign n6406 = n6450 ^ n6451;
  assign n6422 = ~n6454;
  assign n6423 = n6455 ^ n3463;
  assign n6453 = ~n6450;
  assign n6484 = n6519 & n6520;
  assign n6504 = n6539 ^ n6540;
  assign n6541 = ~n6539;
  assign n6475 = ~n6566;
  assign n6554 = n6567 & n6568;
  assign n6543 = n6580 & n6581;
  assign n6544 = ~n6582;
  assign n6552 = ~n6567;
  assign n6555 = n6594 ^ n4106;
  assign n6595 = ~n6594;
  assign n6388 = n6406 ^ n6407;
  assign n6405 = n6421 & n6422;
  assign n6410 = n6422 & n6387;
  assign n6411 = n6423 & n6424;
  assign n6412 = ~n6423;
  assign n6440 = n6452 & n6453;
  assign n6442 = n6484 ^ n3410;
  assign n6486 = n6484 & n3410;
  assign n6485 = ~n6484;
  assign n6348 = n6503 ^ n6504;
  assign n6425 = n6504 & n6503;
  assign n6530 = n6541 & n6542;
  assign n6531 = n6475 & n6430;
  assign n6354 = n6543 ^ n6544;
  assign n6547 = n6552 & n6553;
  assign n6435 = ~n6554;
  assign n2676 = n6555 ^ n6556;
  assign n6545 = ~n6543;
  assign n6583 = n6595 & n6596;
  assign n6373 = n6388 & n131;
  assign n6371 = ~n6388;
  assign n6386 = ~n6405;
  assign n6375 = ~n6410;
  assign n6346 = ~n6411;
  assign n6398 = n6412 & n6413;
  assign n6408 = ~n6440;
  assign n2207 = n6441 ^ n6442;
  assign n6469 = n6485 & n3401;
  assign n6456 = ~n6486;
  assign n6471 = n6348 & n3369;
  assign n6470 = ~n6348;
  assign n6428 = ~n6425;
  assign n6509 = n6354 & n435;
  assign n6505 = ~n6530;
  assign n6473 = ~n6531;
  assign n6507 = ~n6354;
  assign n6521 = n2676 & n6533;
  assign n6495 = n2676 & n5300;
  assign n6532 = n6545 & n6546;
  assign n6480 = ~n6547;
  assign n2777 = ~n2676;
  assign n6557 = ~n6583;
  assign n6363 = n6371 & n6372;
  assign n6301 = ~n6373;
  assign n6339 = n6374 ^ n6375;
  assign n6299 = n6386 & n6387;
  assign n6377 = ~n6398;
  assign n6329 = n6408 & n6409;
  assign n6376 = n2207 & n4714;
  assign n6399 = n2207 & n6414;
  assign n2108 = ~n2207;
  assign n6443 = n6456 & n6457;
  assign n6416 = ~n6469;
  assign n6458 = n6470 & n3353;
  assign n6350 = ~n6471;
  assign n6394 = n6495 ^ n4015;
  assign n6472 = n6505 & n6506;
  assign n6494 = n6507 & n6508;
  assign n6358 = ~n6509;
  assign n6512 = n6480 & n6435;
  assign n5404 = ~n6521;
  assign n6513 = n2777 & n5380;
  assign n6510 = ~n6532;
  assign n6523 = n6557 & n6558;
  assign n4667 = n6338 ^ n6339;
  assign n6257 = n6339 & n6338;
  assign n6341 = ~n6363;
  assign n6340 = ~n6299;
  assign n6289 = n6376 ^ n3410;
  assign n6365 = n6377 & n6346;
  assign n6378 = ~n6329;
  assign n6389 = n2108 & n4771;
  assign n4786 = ~n6399;
  assign n6415 = ~n6443;
  assign n6381 = ~n6458;
  assign n6426 = n6472 ^ n6473;
  assign n6461 = n6394 & n6476;
  assign n6460 = ~n6394;
  assign n6474 = ~n6472;
  assign n6392 = ~n6494;
  assign n6477 = n6510 & n6511;
  assign n6478 = ~n6512;
  assign n5383 = ~n6513;
  assign n2740 = n6522 ^ n6523;
  assign n6524 = ~n6523;
  assign n6151 = ~n4667;
  assign n6327 = n6340 & n6341;
  assign n6298 = n6341 & n6301;
  assign n6342 = n6289 & n6250;
  assign n6343 = ~n6289;
  assign n6330 = ~n6365;
  assign n6364 = n6377 & n6378;
  assign n4774 = ~n6389;
  assign n6379 = n6415 & n6416;
  assign n6305 = n6425 ^ n6426;
  assign n6427 = ~n6426;
  assign n6445 = n6460 & n6356;
  assign n6396 = ~n6461;
  assign n6459 = n6474 & n6475;
  assign n6444 = n6477 ^ n6478;
  assign n6479 = ~n6477;
  assign n6487 = n2740 & n6496;
  assign n6463 = n2740 & n5295;
  assign n2724 = ~n2740;
  assign n6514 = n6524 & n6525;
  assign n6258 = n6298 ^ n6299;
  assign n6300 = ~n6327;
  assign n6303 = n6329 ^ n6330;
  assign n6261 = ~n6342;
  assign n6328 = n6343 & n6344;
  assign n6345 = ~n6364;
  assign n6347 = n6379 ^ n3369;
  assign n6380 = ~n6379;
  assign n6272 = ~n6305;
  assign n6311 = n6427 & n6428;
  assign n6433 = n6444 & n434;
  assign n6360 = ~n6445;
  assign n6429 = ~n6459;
  assign n6431 = ~n6444;
  assign n6436 = n6463 ^ n4044;
  assign n6462 = n6479 & n6480;
  assign n6481 = n2724 & n5341;
  assign n5368 = ~n6487;
  assign n6488 = ~n6514;
  assign n4653 = n6257 ^ n6258;
  assign n6259 = ~n6258;
  assign n6199 = n6300 & n6301;
  assign n6287 = n6303 & n130;
  assign n6285 = ~n6303;
  assign n6302 = ~n6328;
  assign n6331 = n6345 & n6346;
  assign n2130 = n6347 ^ n6348;
  assign n6366 = n6380 & n6381;
  assign n6314 = ~n6311;
  assign n6390 = n6429 & n6430;
  assign n6417 = n6431 & n6432;
  assign n6278 = ~n6433;
  assign n6420 = n6436 & n6437;
  assign n6418 = ~n6436;
  assign n6434 = ~n6462;
  assign n5344 = ~n6481;
  assign n6447 = n6488 & n6489;
  assign n6065 = ~n4653;
  assign n6161 = n6259 & n6257;
  assign n6247 = ~n6199;
  assign n6270 = n6285 & n6286;
  assign n6212 = ~n6287;
  assign n6269 = n2130 & n4673;
  assign n6288 = ~n6331;
  assign n2151 = ~n2130;
  assign n6349 = ~n6366;
  assign n6353 = n435 ^ n6390;
  assign n6391 = ~n6390;
  assign n6321 = ~n6417;
  assign n6400 = n6418 & n6419;
  assign n6282 = ~n6420;
  assign n6393 = n6434 & n6435;
  assign n2556 = n6446 ^ n6447;
  assign n6448 = ~n6447;
  assign n6196 = n6269 ^ n3353;
  assign n6248 = ~n6270;
  assign n6249 = n6288 ^ n6289;
  assign n6284 = n6288 & n6302;
  assign n6304 = n6349 & n6350;
  assign n6312 = n6353 ^ n6354;
  assign n6382 = n6391 & n6392;
  assign n6383 = n6321 & n6278;
  assign n6355 = n6393 ^ n6394;
  assign n6325 = ~n6400;
  assign n6395 = ~n6393;
  assign n6401 = n2556 & n5327;
  assign n6385 = n2556 & n5213;
  assign n2664 = ~n2556;
  assign n6438 = n6448 & n6449;
  assign n6233 = n6247 & n6248;
  assign n6225 = n6249 ^ n6250;
  assign n6236 = n6248 & n6212;
  assign n6260 = ~n6284;
  assign n6262 = n6304 ^ n6305;
  assign n6307 = n6304 & n3318;
  assign n6290 = n6311 ^ n6312;
  assign n6306 = ~n6304;
  assign n6313 = ~n6312;
  assign n6332 = n6355 ^ n6356;
  assign n6357 = ~n6382;
  assign n6319 = ~n6383;
  assign n6322 = n6325 & n6282;
  assign n6243 = n6385 ^ n3946;
  assign n6384 = n6395 & n6396;
  assign n5329 = ~n6401;
  assign n6397 = n2664 & n6402;
  assign n6403 = ~n6438;
  assign n6215 = n6225 & n129;
  assign n6211 = ~n6233;
  assign n6213 = ~n6225;
  assign n6200 = ~n6236;
  assign n6234 = n6260 & n6261;
  assign n2039 = n3318 ^ n6262;
  assign n6273 = n6290 & n3278;
  assign n6291 = n6306 & n3321;
  assign n6271 = ~n6307;
  assign n6274 = ~n6290;
  assign n6275 = n6313 & n6314;
  assign n6317 = n6332 & n433;
  assign n6315 = ~n6332;
  assign n6318 = n6357 & n6358;
  assign n6351 = n6243 & n6361;
  assign n6352 = ~n6243;
  assign n6359 = ~n6384;
  assign n5309 = ~n6397;
  assign n6367 = n6403 & n6404;
  assign n6162 = n6199 ^ n6200;
  assign n6139 = n6211 & n6212;
  assign n6197 = n6213 & n6214;
  assign n6141 = ~n6215;
  assign n6226 = n6234 & n6235;
  assign n6198 = n2039 & n4626;
  assign n6227 = n2039 & n6237;
  assign n6216 = ~n6234;
  assign n2045 = ~n2039;
  assign n6263 = n6271 & n6272;
  assign n6167 = ~n6273;
  assign n6264 = n6274 & n3286;
  assign n6239 = ~n6291;
  assign n6308 = n6315 & n6316;
  assign n6206 = ~n6317;
  assign n6276 = n6318 ^ n6319;
  assign n6320 = ~n6318;
  assign n6208 = ~n6351;
  assign n6333 = n6352 & n6204;
  assign n6323 = n6359 & n6360;
  assign n2608 = n6367 ^ n6368;
  assign n6369 = ~n6367;
  assign n4595 = n6161 ^ n6162;
  assign n6099 = n6162 & n6161;
  assign n6183 = ~n6139;
  assign n6182 = ~n6197;
  assign n6082 = n6198 ^ n3318;
  assign n6180 = n6216 ^ n6196;
  assign n6217 = n6216 & n6181;
  assign n6195 = ~n6226;
  assign n4718 = ~n6227;
  assign n6218 = n2045 & n4699;
  assign n6238 = ~n6263;
  assign n6202 = ~n6264;
  assign n6087 = n6275 ^ n6276;
  assign n6191 = n6276 & n6275;
  assign n6241 = ~n6308;
  assign n6309 = n6320 & n6321;
  assign n6126 = n6322 ^ n6323;
  assign n6245 = ~n6333;
  assign n6324 = ~n6323;
  assign n6335 = n2608 & n5291;
  assign n2486 = ~n2608;
  assign n6362 = n6369 & n6370;
  assign n5961 = ~n4595;
  assign n6150 = n6180 ^ n6181;
  assign n6165 = n6182 & n6183;
  assign n6138 = n6182 & n6141;
  assign n6187 = n6195 & n6196;
  assign n6164 = ~n6217;
  assign n4701 = ~n6218;
  assign n6188 = n6238 & n6239;
  assign n6228 = n6202 & n6167;
  assign n6265 = n6241 & n6206;
  assign n6279 = n6126 & n6292;
  assign n6277 = ~n6309;
  assign n6280 = ~n6126;
  assign n6310 = n6324 & n6325;
  assign n6326 = n2486 & n6334;
  assign n5272 = ~n6335;
  assign n6293 = n2486 & n5150;
  assign n6336 = ~n6362;
  assign n6100 = n6138 ^ n6139;
  assign n6137 = n6150 & n128;
  assign n6135 = ~n6150;
  assign n6140 = ~n6165;
  assign n6163 = ~n6187;
  assign n6201 = ~n6188;
  assign n6189 = ~n6228;
  assign n6230 = ~n6265;
  assign n6229 = n6277 & n6278;
  assign n6173 = ~n6279;
  assign n6266 = n6280 & n432;
  assign n6267 = n6293 ^ n3913;
  assign n6281 = ~n6310;
  assign n5293 = ~n6326;
  assign n6294 = n6336 & n6337;
  assign n4576 = n6099 ^ n6100;
  assign n6103 = ~n6100;
  assign n6116 = n6135 & n6136;
  assign n6062 = ~n6137;
  assign n6047 = n6140 & n6141;
  assign n6117 = n6163 & n6164;
  assign n1979 = n6188 ^ n6189;
  assign n6190 = n6201 & n6202;
  assign n6192 = n6229 ^ n6230;
  assign n6240 = ~n6229;
  assign n6128 = ~n6266;
  assign n6253 = n6267 & n6268;
  assign n6242 = n6281 & n6282;
  assign n6251 = ~n6267;
  assign n6254 = n6294 ^ n6295;
  assign n6296 = ~n6294;
  assign n5914 = ~n4576;
  assign n6005 = n6103 & n6099;
  assign n6101 = ~n6116;
  assign n6081 = n6117 ^ n6118;
  assign n6102 = ~n6047;
  assign n6121 = n6117 & n6118;
  assign n6119 = ~n6117;
  assign n6152 = n1979 & n4667;
  assign n1976 = ~n1979;
  assign n6166 = ~n6190;
  assign n5986 = n6191 ^ n6192;
  assign n6089 = n6192 & n6191;
  assign n6231 = n6240 & n6241;
  assign n6203 = n6242 ^ n6243;
  assign n6246 = n6251 & n6252;
  assign n6132 = ~n6253;
  assign n2401 = n3901 ^ n6254;
  assign n6244 = ~n6242;
  assign n6283 = n6296 & n6297;
  assign n5980 = n6081 ^ n6082;
  assign n6010 = ~n6005;
  assign n6083 = n6101 & n6102;
  assign n6084 = n6101 & n6062;
  assign n6110 = n6119 & n6120;
  assign n6104 = ~n6121;
  assign n6111 = n1976 & n4613;
  assign n6142 = n1976 & n6151;
  assign n4669 = ~n6152;
  assign n6122 = n6166 & n6167;
  assign n6154 = n5986 & n3171;
  assign n6153 = ~n5986;
  assign n6092 = n6203 ^ n6204;
  assign n6205 = ~n6231;
  assign n6220 = n2401 & n5230;
  assign n6193 = n2401 & n5185;
  assign n6232 = n6244 & n6245;
  assign n6178 = ~n6246;
  assign n2403 = ~n2401;
  assign n6255 = ~n6283;
  assign n6046 = n5980 & n143;
  assign n6044 = ~n5980;
  assign n6061 = ~n6083;
  assign n6048 = ~n6084;
  assign n6085 = n6104 & n6082;
  assign n6064 = ~n6110;
  assign n6031 = n6111 ^ n3278;
  assign n6086 = n6122 ^ n3258;
  assign n6124 = n6122 & n3258;
  assign n4688 = ~n6142;
  assign n6123 = ~n6122;
  assign n6143 = n6153 & n3218;
  assign n5989 = ~n6154;
  assign n6170 = n6092 & n447;
  assign n6168 = ~n6092;
  assign n6096 = n6193 ^ n3901;
  assign n6171 = n6205 & n6206;
  assign n6175 = n6178 & n6132;
  assign n6209 = n2403 & n6219;
  assign n5257 = ~n6220;
  assign n6207 = ~n6232;
  assign n6222 = n6255 & n6256;
  assign n6040 = n6044 & n6045;
  assign n5964 = ~n6046;
  assign n6006 = n6047 ^ n6048;
  assign n6029 = n6061 & n6062;
  assign n6063 = ~n6085;
  assign n6077 = n6031 & n5982;
  assign n1927 = n6086 ^ n6087;
  assign n6075 = ~n6031;
  assign n6112 = n6123 & n3223;
  assign n6105 = ~n6124;
  assign n6036 = ~n6143;
  assign n6155 = n6168 & n6169;
  assign n6056 = ~n6170;
  assign n6125 = n432 ^ n6171;
  assign n6158 = n6096 & n6174;
  assign n6157 = ~n6096;
  assign n6172 = ~n6171;
  assign n6176 = n6207 & n6208;
  assign n5233 = ~n6209;
  assign n2285 = n6221 ^ n6222;
  assign n6223 = ~n6222;
  assign n4516 = n6005 ^ n6006;
  assign n5979 = n143 ^ n6029;
  assign n6007 = ~n6040;
  assign n6009 = ~n6006;
  assign n6008 = ~n6029;
  assign n6030 = n6063 & n6064;
  assign n6049 = n1927 & n6065;
  assign n6066 = n6075 & n6076;
  assign n6033 = ~n6077;
  assign n1917 = ~n1927;
  assign n6088 = n6105 & n6087;
  assign n6068 = ~n6112;
  assign n6090 = n6125 ^ n6126;
  assign n6094 = ~n6155;
  assign n6145 = n6157 & n6054;
  assign n6098 = ~n6158;
  assign n6156 = n6172 & n6173;
  assign n5970 = n6175 ^ n6176;
  assign n6177 = ~n6176;
  assign n6184 = n2285 & n6194;
  assign n6160 = n2285 & n5145;
  assign n2426 = ~n2285;
  assign n6210 = n6223 & n6224;
  assign n5939 = n5979 ^ n5980;
  assign n5787 = ~n4516;
  assign n5995 = n6007 & n6008;
  assign n5938 = n6009 & n6010;
  assign n5981 = n6030 ^ n6031;
  assign n6032 = ~n6030;
  assign n6012 = n1917 & n4582;
  assign n6041 = n1917 & n4653;
  assign n4633 = ~n6049;
  assign n5984 = ~n6066;
  assign n6067 = ~n6088;
  assign n6069 = n6089 ^ n6090;
  assign n6014 = n6090 & n6089;
  assign n6129 = n5970 & n6144;
  assign n6058 = ~n6145;
  assign n6127 = ~n6156;
  assign n6130 = ~n5970;
  assign n6026 = n6160 ^ n3852;
  assign n6159 = n6177 & n6178;
  assign n6179 = n2426 & n5193;
  assign n5219 = ~n6184;
  assign n6185 = ~n6210;
  assign n4472 = n5938 ^ n5939;
  assign n5940 = ~n5939;
  assign n5877 = n5981 ^ n5982;
  assign n5963 = ~n5995;
  assign n5941 = ~n5938;
  assign n5945 = n6012 ^ n3223;
  assign n6011 = n6032 & n6033;
  assign n4655 = ~n6041;
  assign n6034 = n6067 & n6068;
  assign n6051 = n6069 & n3152;
  assign n6050 = ~n6069;
  assign n6091 = n6127 & n6128;
  assign n6022 = ~n6129;
  assign n6113 = n6130 & n446;
  assign n6114 = n6026 & n6133;
  assign n6115 = ~n6026;
  assign n6131 = ~n6159;
  assign n5195 = ~n6179;
  assign n6146 = n6185 & n6186;
  assign n5760 = ~n4472;
  assign n5833 = n5940 & n5941;
  assign n5942 = n5877 & n5959;
  assign n5920 = n5963 & n5964;
  assign n5943 = ~n5877;
  assign n5966 = n5945 & n5985;
  assign n5965 = ~n5945;
  assign n5983 = ~n6011;
  assign n5987 = n6034 ^ n3171;
  assign n6035 = ~n6034;
  assign n6042 = n6050 & n3160;
  assign n5899 = ~n6051;
  assign n6052 = n6091 ^ n6092;
  assign n6093 = ~n6091;
  assign n5974 = ~n6113;
  assign n6028 = ~n6114;
  assign n6106 = n6115 & n5972;
  assign n6095 = n6131 & n6132;
  assign n6107 = n6146 ^ n6147;
  assign n6148 = ~n6146;
  assign n5836 = ~n5833;
  assign n5876 = n142 ^ n5920;
  assign n5911 = ~n5942;
  assign n5921 = n5943 & n142;
  assign n5912 = ~n5920;
  assign n5960 = n5965 & n5894;
  assign n5946 = ~n5966;
  assign n5944 = n5983 & n5984;
  assign n1840 = n5986 ^ n5987;
  assign n6013 = n6035 & n6036;
  assign n5952 = ~n6042;
  assign n6015 = n447 ^ n6052;
  assign n6078 = n6093 & n6094;
  assign n6053 = n6095 ^ n6096;
  assign n5976 = ~n6106;
  assign n2220 = n3775 ^ n6107;
  assign n6097 = ~n6095;
  assign n6134 = n6148 & n6149;
  assign n5834 = n5876 ^ n5877;
  assign n5892 = n5911 & n5912;
  assign n5867 = ~n5921;
  assign n5893 = n5944 ^ n5945;
  assign n5896 = ~n5960;
  assign n5913 = n1840 & n4536;
  assign n5948 = n1840 & n5961;
  assign n5947 = ~n5944;
  assign n1867 = ~n1840;
  assign n5988 = ~n6013;
  assign n5996 = n5952 & n5899;
  assign n5818 = n6014 ^ n6015;
  assign n6016 = ~n6015;
  assign n5884 = n6053 ^ n6054;
  assign n6055 = ~n6078;
  assign n6070 = n2220 & n6080;
  assign n6043 = n2220 & n5102;
  assign n6079 = n6097 & n6098;
  assign n2388 = ~n2220;
  assign n6108 = ~n6134;
  assign n4430 = n5833 ^ n5834;
  assign n5835 = ~n5834;
  assign n5866 = ~n5892;
  assign n5868 = n5893 ^ n5894;
  assign n5878 = n5913 ^ n3218;
  assign n5922 = n5946 & n5947;
  assign n5923 = n1867 & n4595;
  assign n4619 = ~n5948;
  assign n5949 = n5988 & n5989;
  assign n5968 = n5818 & n3094;
  assign n5950 = ~n5996;
  assign n5967 = ~n5818;
  assign n5925 = n6016 & n6014;
  assign n6019 = n5884 & n445;
  assign n6017 = ~n5884;
  assign n6023 = n6043 ^ n3775;
  assign n6020 = n6055 & n6056;
  assign n6059 = n2388 & n5153;
  assign n5178 = ~n6070;
  assign n6057 = ~n6079;
  assign n6071 = n6108 & n6109;
  assign n5669 = ~n4430;
  assign n5730 = n5835 & n5836;
  assign n5782 = n5866 & n5867;
  assign n5853 = n5868 & n141;
  assign n5851 = ~n5868;
  assign n5871 = n5878 & n5879;
  assign n5869 = ~n5878;
  assign n5895 = ~n5922;
  assign n4598 = ~n5923;
  assign n1825 = n5949 ^ n5950;
  assign n5951 = ~n5949;
  assign n5962 = n5967 & n3096;
  assign n5858 = ~n5968;
  assign n5928 = ~n5925;
  assign n5997 = n6017 & n6018;
  assign n5886 = ~n6019;
  assign n5969 = n446 ^ n6020;
  assign n5999 = n6023 & n6024;
  assign n6000 = ~n6023;
  assign n6021 = ~n6020;
  assign n6025 = n6057 & n6058;
  assign n5156 = ~n6059;
  assign n6037 = n6071 ^ n6072;
  assign n6073 = ~n6071;
  assign n5812 = ~n5782;
  assign n5837 = n5851 & n5852;
  assign n5784 = ~n5853;
  assign n5854 = n5869 & n5870;
  assign n5796 = ~n5871;
  assign n5785 = n5895 & n5896;
  assign n5897 = n1825 & n5914;
  assign n1812 = ~n1825;
  assign n5924 = n5951 & n5952;
  assign n5821 = ~n5962;
  assign n5926 = n5969 ^ n5970;
  assign n5934 = ~n5997;
  assign n5888 = ~n5999;
  assign n5990 = n6000 & n6001;
  assign n5998 = n6021 & n6022;
  assign n5971 = n6025 ^ n6026;
  assign n2262 = n3639 ^ n6037;
  assign n6027 = ~n6025;
  assign n6060 = n6073 & n6074;
  assign n5813 = ~n5837;
  assign n5827 = ~n5854;
  assign n5828 = ~n5785;
  assign n5855 = n1812 & n4466;
  assign n4560 = ~n5897;
  assign n5880 = n1812 & n4576;
  assign n5898 = ~n5924;
  assign n5900 = n5925 ^ n5926;
  assign n5927 = ~n5926;
  assign n5953 = n5971 ^ n5972;
  assign n5936 = ~n5990;
  assign n5973 = ~n5998;
  assign n5991 = n2262 & n6003;
  assign n6002 = n6027 & n6028;
  assign n2104 = ~n2262;
  assign n6038 = ~n6060;
  assign n5799 = n5812 & n5813;
  assign n5781 = n5813 & n5784;
  assign n5814 = n5827 & n5828;
  assign n5815 = n5827 & n5796;
  assign n5723 = n5855 ^ n3160;
  assign n4578 = ~n5880;
  assign n5856 = n5898 & n5899;
  assign n5882 = n5900 & n3106;
  assign n5881 = ~n5900;
  assign n5839 = n5927 & n5928;
  assign n5931 = n5953 & n444;
  assign n5929 = ~n5953;
  assign n5954 = n5936 & n5888;
  assign n5932 = n5973 & n5974;
  assign n5120 = ~n5991;
  assign n5977 = n2104 & n5117;
  assign n5955 = n2104 & n5050;
  assign n5975 = ~n6002;
  assign n5992 = n6038 & n6039;
  assign n5743 = n5781 ^ n5782;
  assign n5783 = ~n5799;
  assign n5795 = ~n5814;
  assign n5786 = ~n5815;
  assign n5817 = n5723 & n5829;
  assign n5816 = ~n5723;
  assign n5819 = n5856 ^ n3094;
  assign n5857 = ~n5856;
  assign n5872 = n5881 & n3100;
  assign n5792 = ~n5882;
  assign n5915 = n5929 & n5930;
  assign n5807 = ~n5931;
  assign n5883 = n445 ^ n5932;
  assign n5902 = ~n5954;
  assign n5805 = n5955 ^ n3639;
  assign n5933 = ~n5932;
  assign n5901 = n5975 & n5976;
  assign n5140 = ~n5977;
  assign n5956 = n5992 ^ n3569;
  assign n5994 = n5992 & n6004;
  assign n5993 = ~n5992;
  assign n5620 = n5730 ^ n5743;
  assign n5683 = n5743 & n5730;
  assign n5731 = ~n5743;
  assign n5744 = n5783 & n5784;
  assign n5745 = n5785 ^ n5786;
  assign n5756 = n5795 & n5796;
  assign n5800 = n5816 & n5757;
  assign n5726 = ~n5817;
  assign n1752 = n5818 ^ n5819;
  assign n5838 = n5857 & n5858;
  assign n5752 = ~n5872;
  assign n5840 = n5883 ^ n5884;
  assign n5873 = n5901 ^ n5902;
  assign n5844 = ~n5915;
  assign n5903 = n5805 & n5847;
  assign n5916 = n5933 & n5934;
  assign n5904 = ~n5805;
  assign n2182 = n5956 ^ n5957;
  assign n5935 = ~n5901;
  assign n5978 = n5993 & n5957;
  assign n5909 = ~n5994;
  assign n5632 = n5730 ^ n5731;
  assign n5716 = n5744 ^ n5745;
  assign n5748 = n5745 & n140;
  assign n5724 = n5756 ^ n5757;
  assign n5718 = ~n5744;
  assign n5746 = ~n5745;
  assign n5758 = ~n5756;
  assign n5761 = n1752 & n4469;
  assign n5788 = n1752 & n4516;
  assign n5759 = ~n5800;
  assign n1786 = ~n1752;
  assign n5820 = ~n5838;
  assign n5789 = n5792 & n5752;
  assign n5822 = n5839 ^ n5840;
  assign n5802 = n5840 & n5839;
  assign n5861 = n5873 & n443;
  assign n5841 = n5844 & n5807;
  assign n5859 = ~n5873;
  assign n5849 = ~n5903;
  assign n5889 = n5904 & n5905;
  assign n5885 = ~n5916;
  assign n5907 = n2182 & n5073;
  assign n5917 = n5935 & n5936;
  assign n2194 = ~n2182;
  assign n5958 = n5909 & n3557;
  assign n5919 = ~n5978;
  assign n5684 = n140 ^ n5716;
  assign n5667 = n5723 ^ n5724;
  assign n5732 = n5746 & n5747;
  assign n5687 = ~n5748;
  assign n5749 = n5758 & n5759;
  assign n5697 = n5761 ^ n3096;
  assign n5767 = n1786 & n5787;
  assign n4542 = ~n5788;
  assign n5790 = n5820 & n5821;
  assign n5801 = n5822 & n3085;
  assign n5689 = ~n5822;
  assign n5845 = n5859 & n5860;
  assign n5740 = ~n5861;
  assign n5842 = n5885 & n5886;
  assign n5810 = ~n5889;
  assign n5890 = n2194 & n5906;
  assign n5076 = ~n5907;
  assign n5862 = n2194 & n4985;
  assign n5887 = ~n5917;
  assign n5918 = ~n5958;
  assign n5937 = n5919 & n3569;
  assign n4365 = n5683 ^ n5684;
  assign n5613 = n5684 & n5683;
  assign n5695 = n5667 & n139;
  assign n5693 = ~n5667;
  assign n5717 = ~n5732;
  assign n5728 = n5697 & n5733;
  assign n5725 = ~n5749;
  assign n5727 = ~n5697;
  assign n4519 = ~n5767;
  assign n1687 = n5789 ^ n5790;
  assign n5791 = ~n5790;
  assign n5722 = ~n5801;
  assign n5797 = n5689 & n3078;
  assign n5803 = n5841 ^ n5842;
  assign n5776 = ~n5845;
  assign n5778 = n5862 ^ n3557;
  assign n5843 = ~n5842;
  assign n5846 = n5887 & n5888;
  assign n5078 = ~n5890;
  assign n5910 = n5918 & n5919;
  assign n5908 = ~n5937;
  assign n5582 = ~n4365;
  assign n5685 = n5693 & n5694;
  assign n5643 = ~n5695;
  assign n5703 = n5717 & n5718;
  assign n5696 = n5725 & n5726;
  assign n5719 = n5727 & n5675;
  assign n5698 = ~n5728;
  assign n5750 = n1687 & n5760;
  assign n5729 = n1687 & n4416;
  assign n1743 = ~n1687;
  assign n5768 = n5791 & n5792;
  assign n5692 = ~n5797;
  assign n5671 = n5802 ^ n5803;
  assign n5735 = n5803 & n5802;
  assign n5808 = n5776 & n5740;
  assign n5823 = n5778 & n5831;
  assign n5830 = n5843 & n5844;
  assign n5804 = n5846 ^ n5847;
  assign n5824 = ~n5778;
  assign n5848 = ~n5846;
  assign n5891 = n5908 & n5909;
  assign n5874 = ~n5910;
  assign n5664 = ~n5685;
  assign n5674 = n5696 ^ n5697;
  assign n5686 = ~n5703;
  assign n5699 = ~n5696;
  assign n5677 = ~n5719;
  assign n5628 = n5729 ^ n3106;
  assign n5734 = n1743 & n4472;
  assign n4499 = ~n5750;
  assign n5751 = ~n5768;
  assign n5769 = n5671 & n2955;
  assign n5770 = ~n5671;
  assign n5753 = ~n5735;
  assign n5711 = n5804 ^ n5805;
  assign n5774 = ~n5808;
  assign n5780 = ~n5823;
  assign n5811 = n5824 & n5738;
  assign n5806 = ~n5830;
  assign n5832 = n5848 & n5849;
  assign n5865 = n5874 & n5875;
  assign n5863 = ~n5891;
  assign n5600 = n5674 ^ n5675;
  assign n5666 = n5686 & n5687;
  assign n5688 = n5698 & n5699;
  assign n4475 = ~n5734;
  assign n5720 = n5751 & n5752;
  assign n5673 = ~n5769;
  assign n5762 = n5770 & n3013;
  assign n5771 = n5711 & n5793;
  assign n5772 = ~n5711;
  assign n5773 = n5806 & n5807;
  assign n5742 = ~n5811;
  assign n5809 = ~n5832;
  assign n5850 = n5863 & n5864;
  assign n5826 = ~n5865;
  assign n5641 = n5666 ^ n5667;
  assign n5665 = ~n5666;
  assign n5676 = ~n5688;
  assign n5690 = n5720 ^ n3078;
  assign n5721 = ~n5720;
  assign n5647 = ~n5762;
  assign n5713 = ~n5771;
  assign n5763 = n5772 & n442;
  assign n5736 = n5773 ^ n5774;
  assign n5775 = ~n5773;
  assign n5777 = n5809 & n5810;
  assign n5825 = ~n5850;
  assign n5614 = n139 ^ n5641;
  assign n5655 = n5664 & n5665;
  assign n5648 = n5676 & n5677;
  assign n1667 = n5689 ^ n5690;
  assign n5704 = n5721 & n5722;
  assign n5622 = n5735 ^ n5736;
  assign n5658 = n5736 & n5753;
  assign n5682 = ~n5763;
  assign n5764 = n5775 & n5776;
  assign n5737 = n5777 ^ n5778;
  assign n5779 = ~n5777;
  assign n1998 = n5825 & n5826;
  assign n4302 = n5613 ^ n5614;
  assign n5570 = n5614 & n5613;
  assign n5627 = n5648 ^ n5649;
  assign n5642 = ~n5655;
  assign n5652 = n5648 & n5649;
  assign n5650 = ~n5648;
  assign n5668 = n1667 & n4430;
  assign n5653 = n1667 & n4370;
  assign n1722 = ~n1667;
  assign n5691 = ~n5704;
  assign n5706 = n5622 & n3001;
  assign n5705 = ~n5622;
  assign n5661 = n5737 ^ n5738;
  assign n5739 = ~n5764;
  assign n5765 = n5779 & n5780;
  assign n5754 = n5794 ^ n1998;
  assign n5766 = n1998 & n5798;
  assign n3653 = ~n1998;
  assign n5530 = ~n4302;
  assign n5558 = n5627 ^ n5628;
  assign n5615 = n5642 & n5643;
  assign n5644 = n5650 & n5651;
  assign n5635 = ~n5652;
  assign n5561 = n5653 ^ n3085;
  assign n4455 = ~n5668;
  assign n5656 = n1722 & n5669;
  assign n5670 = n5691 & n5692;
  assign n5700 = n5705 & n2992;
  assign n5624 = ~n5706;
  assign n5709 = n5661 & n441;
  assign n5707 = ~n5661;
  assign n5710 = n5739 & n5740;
  assign n5053 = n5754 ^ n5755;
  assign n5741 = ~n5765;
  assign n5680 = n5766 ^ n3484;
  assign n5603 = n5558 & n137;
  assign n5592 = n5615 ^ n5600;
  assign n5601 = ~n5558;
  assign n5617 = n5615 & n5626;
  assign n5630 = n5561 & n5634;
  assign n5629 = n5635 & n5628;
  assign n5616 = ~n5615;
  assign n5606 = ~n5644;
  assign n5631 = ~n5561;
  assign n4432 = ~n5656;
  assign n5645 = n5670 ^ n5671;
  assign n5672 = ~n5670;
  assign n5598 = ~n5700;
  assign n5701 = n5707 & n5708;
  assign n5640 = ~n5709;
  assign n5678 = n5710 ^ n5711;
  assign n5712 = ~n5710;
  assign n5714 = n5741 & n5742;
  assign n5057 = ~n5053;
  assign n5571 = n138 ^ n5592;
  assign n5594 = n5601 & n5602;
  assign n5538 = ~n5603;
  assign n5604 = n5616 & n138;
  assign n5599 = ~n5617;
  assign n5605 = ~n5629;
  assign n5564 = ~n5630;
  assign n5618 = n5631 & n5586;
  assign n1591 = n5645 ^ n3013;
  assign n5657 = n5672 & n5673;
  assign n5659 = n442 ^ n5678;
  assign n5663 = ~n5701;
  assign n5702 = n5712 & n5713;
  assign n5679 = n5714 ^ n5715;
  assign n5490 = n5570 ^ n5571;
  assign n5515 = n5571 & n5570;
  assign n5560 = ~n5594;
  assign n5593 = n5599 & n5600;
  assign n5581 = ~n5604;
  assign n5585 = n5605 & n5606;
  assign n5588 = ~n5618;
  assign n5619 = n1591 & n5632;
  assign n1684 = ~n1591;
  assign n5646 = ~n5657;
  assign n5577 = n5658 ^ n5659;
  assign n5609 = n5659 & n5658;
  assign n5612 = n5679 ^ n5680;
  assign n5681 = ~n5702;
  assign n4264 = ~n5490;
  assign n5562 = n5585 ^ n5586;
  assign n5580 = ~n5593;
  assign n5587 = ~n5585;
  assign n4386 = ~n5619;
  assign n5607 = n1684 & n5620;
  assign n5595 = n1684 & n4359;
  assign n5621 = n5646 & n5647;
  assign n5636 = n5577 & n2932;
  assign n5637 = ~n5577;
  assign n5625 = ~n5609;
  assign n5660 = n5681 & n5682;
  assign n5518 = n5561 ^ n5562;
  assign n5557 = n5580 & n5581;
  assign n5583 = n5587 & n5588;
  assign n5523 = n5595 ^ n2955;
  assign n4412 = ~n5607;
  assign n5596 = n5621 ^ n5622;
  assign n5623 = ~n5621;
  assign n5553 = ~n5636;
  assign n5633 = n5637 & n2873;
  assign n5638 = n5660 ^ n5661;
  assign n5662 = ~n5660;
  assign n5545 = n5518 & n136;
  assign n5536 = n5557 ^ n5558;
  assign n5543 = ~n5518;
  assign n5559 = ~n5557;
  assign n5563 = ~n5583;
  assign n5575 = n5523 & n5547;
  assign n5573 = ~n5523;
  assign n4409 = n4412 & n4386;
  assign n1528 = n2992 ^ n5596;
  assign n5608 = n5623 & n5624;
  assign n5579 = ~n5633;
  assign n5610 = n441 ^ n5638;
  assign n5654 = n5662 & n5663;
  assign n5516 = n137 ^ n5536;
  assign n5539 = n5543 & n5544;
  assign n5497 = ~n5545;
  assign n5554 = n5559 & n5560;
  assign n5546 = n5563 & n5564;
  assign n5566 = n5573 & n5574;
  assign n5525 = ~n5575;
  assign n5572 = n1528 & n5582;
  assign n1608 = ~n1528;
  assign n5597 = ~n5608;
  assign n5511 = n5609 ^ n5610;
  assign n5568 = n5610 & n5625;
  assign n5639 = ~n5654;
  assign n4223 = n5515 ^ n5516;
  assign n5476 = n5516 & n5515;
  assign n5519 = ~n5539;
  assign n5522 = n5546 ^ n5547;
  assign n5537 = ~n5554;
  assign n5548 = ~n5546;
  assign n5549 = ~n5566;
  assign n4343 = ~n5572;
  assign n5565 = n1608 & n4365;
  assign n5555 = n1608 & n4235;
  assign n5576 = n5597 & n5598;
  assign n5589 = n5511 & n2879;
  assign n5590 = ~n5511;
  assign n5611 = n5639 & n5640;
  assign n5457 = ~n4223;
  assign n5479 = ~n5476;
  assign n5456 = n5522 ^ n5523;
  assign n5517 = n5537 & n5538;
  assign n5540 = n5548 & n5549;
  assign n5505 = n5555 ^ n2992;
  assign n4367 = ~n5565;
  assign n5556 = n5576 ^ n5577;
  assign n5578 = ~n5576;
  assign n5514 = ~n5589;
  assign n5584 = n5590 & n2829;
  assign n5591 = n5611 ^ n5612;
  assign n5502 = n5456 & n5509;
  assign n5495 = n5517 ^ n5518;
  assign n5503 = ~n5456;
  assign n5520 = ~n5517;
  assign n5524 = ~n5540;
  assign n5531 = n5505 & n5541;
  assign n5532 = ~n5505;
  assign n1499 = n5556 ^ n2932;
  assign n5567 = n5578 & n5579;
  assign n5535 = ~n5584;
  assign n5569 = n440 ^ n5591;
  assign n5477 = n136 ^ n5495;
  assign n5481 = ~n5502;
  assign n5498 = n5503 & n151;
  assign n5510 = n5519 & n5520;
  assign n5504 = n5524 & n5525;
  assign n5507 = ~n5531;
  assign n5527 = n5532 & n5484;
  assign n5529 = n1499 & n4302;
  assign n5521 = n1499 & n4249;
  assign n1551 = ~n1499;
  assign n5552 = ~n5567;
  assign n5473 = n5568 ^ n5569;
  assign n4180 = n5476 ^ n5477;
  assign n5478 = ~n5477;
  assign n5459 = ~n5498;
  assign n5483 = n5504 ^ n5505;
  assign n5496 = ~n5510;
  assign n5506 = ~n5504;
  assign n5444 = n5521 ^ n2873;
  assign n5487 = ~n5527;
  assign n4325 = ~n5529;
  assign n5526 = n1551 & n5530;
  assign n5533 = n5552 & n5553;
  assign n5550 = n5473 & n2850;
  assign n5551 = ~n5473;
  assign n5401 = ~n4180;
  assign n5433 = n5478 & n5479;
  assign n5438 = n5483 ^ n5484;
  assign n5480 = n5496 & n5497;
  assign n5499 = n5506 & n5507;
  assign n5500 = n5444 & n5508;
  assign n5501 = ~n5444;
  assign n4305 = ~n5526;
  assign n5512 = n5533 ^ n2829;
  assign n5534 = ~n5533;
  assign n5475 = ~n5550;
  assign n5542 = n5551 & n2860;
  assign n5436 = ~n5433;
  assign n5465 = n5438 & n150;
  assign n5455 = n151 ^ n5480;
  assign n5463 = ~n5438;
  assign n5482 = ~n5480;
  assign n5486 = ~n5499;
  assign n5446 = ~n5500;
  assign n5491 = n5501 & n5467;
  assign n1523 = n5511 ^ n5512;
  assign n5528 = n5534 & n5535;
  assign n5494 = ~n5542;
  assign n5434 = n5455 ^ n5456;
  assign n5460 = n5463 & n5464;
  assign n5417 = ~n5465;
  assign n5470 = n5481 & n5482;
  assign n5466 = n5486 & n5487;
  assign n5469 = ~n5491;
  assign n5489 = n1523 & n4264;
  assign n1513 = ~n1523;
  assign n5513 = ~n5528;
  assign n5364 = n5433 ^ n5434;
  assign n5435 = ~n5434;
  assign n5440 = ~n5460;
  assign n5443 = n5466 ^ n5467;
  assign n5458 = ~n5470;
  assign n5468 = ~n5466;
  assign n4266 = ~n5489;
  assign n5485 = n1513 & n5490;
  assign n5471 = n1513 & n4202;
  assign n5492 = n5513 & n5514;
  assign n5369 = ~n5364;
  assign n5395 = n5435 & n5436;
  assign n5398 = n5443 ^ n5444;
  assign n5437 = n5458 & n5459;
  assign n5461 = n5468 & n5469;
  assign n5406 = n5471 ^ n2829;
  assign n4286 = ~n5485;
  assign n5472 = n5492 ^ n2860;
  assign n5493 = ~n5492;
  assign n5424 = n5398 & n149;
  assign n5415 = n5437 ^ n5438;
  assign n5422 = ~n5398;
  assign n5439 = ~n5437;
  assign n5445 = ~n5461;
  assign n5452 = n5406 & n5426;
  assign n5450 = ~n5406;
  assign n1471 = n5472 ^ n5473;
  assign n5488 = n5493 & n5494;
  assign n5396 = n150 ^ n5415;
  assign n5418 = n5422 & n5423;
  assign n5376 = ~n5424;
  assign n5429 = n5439 & n5440;
  assign n5425 = n5445 & n5446;
  assign n5447 = n5450 & n5451;
  assign n5408 = ~n5452;
  assign n5449 = n1471 & n5457;
  assign n1456 = ~n1471;
  assign n5474 = ~n5488;
  assign n5325 = n5395 ^ n5396;
  assign n5356 = n5396 & n5395;
  assign n5400 = ~n5418;
  assign n5405 = n5425 ^ n5426;
  assign n5416 = ~n5429;
  assign n5427 = ~n5425;
  assign n5428 = ~n5447;
  assign n4225 = ~n5449;
  assign n5442 = n1456 & n4223;
  assign n5430 = n1456 & n4171;
  assign n5462 = n5474 & n5475;
  assign n5330 = ~n5325;
  assign n5359 = ~n5356;
  assign n5361 = n5405 ^ n5406;
  assign n5397 = n5416 & n5417;
  assign n5419 = n5427 & n5428;
  assign n5371 = n5430 ^ n2850;
  assign n4245 = ~n5442;
  assign n5454 = n5462 & n2807;
  assign n5453 = ~n5462;
  assign n5384 = n5361 & n5391;
  assign n5374 = n5397 ^ n5398;
  assign n5385 = ~n5361;
  assign n5399 = ~n5397;
  assign n5407 = ~n5419;
  assign n5410 = n5371 & n5388;
  assign n5411 = ~n5371;
  assign n5448 = n5453 & n2709;
  assign n5432 = ~n5454;
  assign n5357 = n149 ^ n5374;
  assign n5363 = ~n5384;
  assign n5377 = n5385 & n148;
  assign n5392 = n5399 & n5400;
  assign n5387 = n5407 & n5408;
  assign n5390 = ~n5410;
  assign n5409 = n5411 & n5412;
  assign n5431 = n5432 & n5441;
  assign n5421 = ~n5448;
  assign n4024 = n5356 ^ n5357;
  assign n5358 = ~n5357;
  assign n5337 = ~n5377;
  assign n5370 = n5387 ^ n5388;
  assign n5375 = ~n5392;
  assign n5389 = ~n5387;
  assign n5373 = ~n5409;
  assign n5420 = ~n5431;
  assign n5414 = n5421 & n5432;
  assign n5318 = n5358 & n5359;
  assign n5321 = n5370 ^ n5371;
  assign n5360 = n5375 & n5376;
  assign n5378 = n5389 & n5390;
  assign n1362 = n5413 ^ n5414;
  assign n5402 = n5420 & n5421;
  assign n5345 = n5321 & n5352;
  assign n5335 = n5360 ^ n5361;
  assign n5346 = ~n5321;
  assign n5362 = ~n5360;
  assign n5372 = ~n5378;
  assign n5393 = n1362 & n5401;
  assign n5381 = n1362 & n4121;
  assign n5379 = n5402 ^ n2676;
  assign n1327 = ~n1362;
  assign n5403 = ~n5402;
  assign n5319 = n148 ^ n5335;
  assign n5323 = ~n5345;
  assign n5338 = n5346 & n147;
  assign n5353 = n5362 & n5363;
  assign n5347 = n5372 & n5373;
  assign n1349 = n5379 ^ n5380;
  assign n5331 = n5381 ^ n2807;
  assign n5386 = n1327 & n4180;
  assign n4209 = ~n5393;
  assign n5394 = n5403 & n5404;
  assign n3998 = n5318 ^ n5319;
  assign n5279 = n5319 & n5318;
  assign n5304 = ~n5338;
  assign n5332 = n5347 ^ n5348;
  assign n5336 = ~n5353;
  assign n5351 = n5347 & n5348;
  assign n5349 = ~n5347;
  assign n5365 = n1349 & n5369;
  assign n1270 = ~n1349;
  assign n4183 = ~n5386;
  assign n5382 = ~n5394;
  assign n5259 = ~n3998;
  assign n5282 = ~n5279;
  assign n5284 = n5331 ^ n5332;
  assign n5320 = n5336 & n5337;
  assign n5339 = n5349 & n5350;
  assign n5334 = ~n5351;
  assign n5354 = n1270 & n5364;
  assign n4136 = ~n5365;
  assign n5340 = n1270 & n4015;
  assign n5366 = n5382 & n5383;
  assign n5312 = n5284 & n146;
  assign n5302 = n5320 ^ n5321;
  assign n5310 = ~n5284;
  assign n5322 = ~n5320;
  assign n5333 = n5334 & n5331;
  assign n5316 = ~n5339;
  assign n5274 = n5340 ^ n2676;
  assign n4167 = ~n5354;
  assign n5342 = n5366 ^ n2740;
  assign n5367 = ~n5366;
  assign n5280 = n147 ^ n5302;
  assign n5305 = n5310 & n5311;
  assign n5266 = ~n5312;
  assign n5313 = n5322 & n5323;
  assign n5315 = ~n5333;
  assign n4164 = n4167 & n4136;
  assign n1205 = n5341 ^ n5342;
  assign n5355 = n5367 & n5368;
  assign n3951 = n5279 ^ n5280;
  assign n5281 = ~n5280;
  assign n5286 = ~n5305;
  assign n5303 = ~n5313;
  assign n5297 = n5315 & n5316;
  assign n5324 = n1205 & n5330;
  assign n1254 = ~n1205;
  assign n5343 = ~n5355;
  assign n5210 = ~n3951;
  assign n5243 = n5281 & n5282;
  assign n5273 = n5297 ^ n5298;
  assign n5283 = n5303 & n5304;
  assign n5301 = n5297 & n5298;
  assign n5299 = ~n5297;
  assign n4087 = ~n5324;
  assign n5314 = n1254 & n5325;
  assign n5306 = n1254 & n4055;
  assign n5326 = n5343 & n5344;
  assign n5246 = ~n5243;
  assign n5238 = n5273 ^ n5274;
  assign n5264 = n5283 ^ n5284;
  assign n5285 = ~n5283;
  assign n5294 = n5299 & n5300;
  assign n5287 = ~n5301;
  assign n5227 = n5306 ^ n2740;
  assign n4119 = ~n5314;
  assign n5307 = n5326 ^ n5327;
  assign n5328 = ~n5326;
  assign n5244 = n146 ^ n5264;
  assign n5262 = n5238 & n145;
  assign n5260 = ~n5238;
  assign n5275 = n5285 & n5286;
  assign n5276 = n5287 & n5274;
  assign n5268 = ~n5294;
  assign n5289 = n5227 & n5295;
  assign n5288 = ~n5227;
  assign n5296 = n4119 & n4087;
  assign n1228 = n5307 ^ n2664;
  assign n5317 = n5328 & n5329;
  assign n3915 = n5243 ^ n5244;
  assign n5245 = ~n5244;
  assign n5258 = n5260 & n5261;
  assign n5224 = ~n5262;
  assign n5265 = ~n5275;
  assign n5267 = ~n5276;
  assign n5277 = n5288 & n5249;
  assign n5229 = ~n5289;
  assign n4117 = ~n5296;
  assign n1223 = ~n1228;
  assign n5308 = ~n5317;
  assign n5180 = ~n3915;
  assign n5197 = n5245 & n5246;
  assign n5236 = ~n5258;
  assign n5263 = n5265 & n5266;
  assign n5248 = n5267 & n5268;
  assign n5251 = ~n5277;
  assign n5269 = n1223 & n3971;
  assign n5290 = n5308 & n5309;
  assign n5200 = ~n5197;
  assign n5226 = n5248 ^ n5249;
  assign n5237 = ~n5263;
  assign n5250 = ~n5248;
  assign n5189 = n5269 ^ n2556;
  assign n5270 = n5290 ^ n5291;
  assign n5292 = ~n5290;
  assign n5202 = n5226 ^ n5227;
  assign n5234 = n5236 & n5237;
  assign n5222 = n5237 ^ n5238;
  assign n5240 = n5250 & n5251;
  assign n5254 = n5189 & n5213;
  assign n5252 = ~n5189;
  assign n1088 = n2608 ^ n5270;
  assign n5278 = n5292 & n5293;
  assign n5209 = n5202 & n144;
  assign n5198 = n145 ^ n5222;
  assign n5207 = ~n5202;
  assign n5223 = ~n5234;
  assign n5228 = ~n5240;
  assign n5241 = n5252 & n5253;
  assign n5191 = ~n5254;
  assign n5247 = n1088 & n5259;
  assign n5235 = n1088 & n3872;
  assign n1140 = ~n1088;
  assign n5271 = ~n5278;
  assign n3892 = n5197 ^ n5198;
  assign n5203 = n5207 & n5208;
  assign n5167 = ~n5209;
  assign n5199 = ~n5198;
  assign n5201 = n5223 & n5224;
  assign n5212 = n5228 & n5229;
  assign n5172 = n5235 ^ n2608;
  assign n5215 = ~n5241;
  assign n5239 = n1140 & n3998;
  assign n4021 = ~n5247;
  assign n5255 = n5271 & n5272;
  assign n5141 = ~n3892;
  assign n5158 = n5199 & n5200;
  assign n5183 = n5201 ^ n5202;
  assign n5186 = ~n5203;
  assign n5188 = n5212 ^ n5213;
  assign n5187 = ~n5201;
  assign n5214 = ~n5212;
  assign n5220 = n5172 & n5225;
  assign n5221 = ~n5172;
  assign n4001 = ~n5239;
  assign n5231 = n5255 ^ n2401;
  assign n5256 = ~n5255;
  assign n5159 = n144 ^ n5183;
  assign n5184 = n5186 & n5187;
  assign n5126 = n5188 ^ n5189;
  assign n5161 = ~n5158;
  assign n5205 = n5214 & n5215;
  assign n5174 = ~n5220;
  assign n5216 = n5221 & n5150;
  assign n1029 = n5230 ^ n5231;
  assign n5242 = n5256 & n5257;
  assign n5101 = n5158 ^ n5159;
  assign n5160 = ~n5159;
  assign n5168 = n5126 & n5179;
  assign n5166 = ~n5184;
  assign n5169 = ~n5126;
  assign n5190 = ~n5205;
  assign n5152 = ~n5216;
  assign n5211 = n1029 & n3951;
  assign n5196 = n1029 & n3901;
  assign n1074 = ~n1029;
  assign n5232 = ~n5242;
  assign n5091 = ~n5101;
  assign n5104 = n5160 & n5161;
  assign n5146 = n5166 & n5167;
  assign n5148 = ~n5168;
  assign n5162 = n5169 & n159;
  assign n5171 = n5190 & n5191;
  assign n5113 = n5196 ^ n2401;
  assign n5204 = n1074 & n5210;
  assign n3981 = ~n5211;
  assign n5217 = n5232 & n5233;
  assign n5125 = n159 ^ n5146;
  assign n5107 = ~n5104;
  assign n5147 = ~n5146;
  assign n5128 = ~n5162;
  assign n5149 = n5171 ^ n5172;
  assign n5173 = ~n5171;
  assign n5182 = n5113 & n5185;
  assign n5181 = ~n5113;
  assign n3953 = ~n5204;
  assign n5192 = n5217 ^ n2426;
  assign n5218 = ~n5217;
  assign n5105 = n5125 ^ n5126;
  assign n5144 = n5147 & n5148;
  assign n5109 = n5149 ^ n5150;
  assign n5164 = n5173 & n5174;
  assign n5175 = n5181 & n5134;
  assign n5115 = ~n5182;
  assign n974 = n5192 ^ n5193;
  assign n5206 = n5218 & n5219;
  assign n5038 = n5104 ^ n5105;
  assign n5106 = ~n5105;
  assign n5131 = n5109 & n158;
  assign n5127 = ~n5144;
  assign n5129 = ~n5109;
  assign n5151 = ~n5164;
  assign n5136 = ~n5175;
  assign n5170 = n974 & n5180;
  assign n5157 = n974 & n3852;
  assign n1020 = ~n974;
  assign n5194 = ~n5206;
  assign n5055 = ~n5038;
  assign n5061 = n5106 & n5107;
  assign n5108 = n5127 & n5128;
  assign n5121 = n5129 & n5130;
  assign n5086 = ~n5131;
  assign n5133 = n5151 & n5152;
  assign n5068 = n5157 ^ n2285;
  assign n3939 = ~n5170;
  assign n5163 = n1020 & n3915;
  assign n5176 = n5194 & n5195;
  assign n5084 = n5108 ^ n5109;
  assign n5110 = ~n5108;
  assign n5111 = ~n5121;
  assign n5112 = n5133 ^ n5134;
  assign n5135 = ~n5133;
  assign n5143 = n5068 & n5145;
  assign n5142 = ~n5068;
  assign n3918 = ~n5163;
  assign n5154 = n5176 ^ n2220;
  assign n5177 = ~n5176;
  assign n5062 = n158 ^ n5084;
  assign n5103 = n5110 & n5111;
  assign n5064 = n5112 ^ n5113;
  assign n5123 = n5135 & n5136;
  assign n5137 = n5142 & n5093;
  assign n5070 = ~n5143;
  assign n957 = n5153 ^ n5154;
  assign n5165 = n5177 & n5178;
  assign n3701 = n5061 ^ n5062;
  assign n5019 = n5062 & n5061;
  assign n5089 = n5064 & n157;
  assign n5085 = ~n5103;
  assign n5087 = ~n5064;
  assign n5114 = ~n5123;
  assign n5095 = ~n5137;
  assign n5132 = n957 & n5141;
  assign n905 = ~n957;
  assign n5155 = ~n5165;
  assign n5063 = n5085 & n5086;
  assign n5079 = n5087 & n5088;
  assign n5041 = ~n5089;
  assign n5092 = n5114 & n5115;
  assign n5122 = n905 & n3892;
  assign n3869 = ~n5132;
  assign n5116 = n905 & n3665;
  assign n5138 = n5155 & n5156;
  assign n5037 = n5063 ^ n5064;
  assign n5065 = ~n5063;
  assign n5066 = ~n5079;
  assign n5067 = n5092 ^ n5093;
  assign n5094 = ~n5092;
  assign n5026 = n5116 ^ n2220;
  assign n3894 = ~n5122;
  assign n5118 = n5138 ^ n2262;
  assign n5139 = ~n5138;
  assign n5020 = n157 ^ n5037;
  assign n5058 = n5065 & n5066;
  assign n5022 = n5067 ^ n5068;
  assign n5081 = n5094 & n5095;
  assign n5097 = n5026 & n5102;
  assign n5096 = ~n5026;
  assign n844 = n5117 ^ n5118;
  assign n5124 = n5139 & n5140;
  assign n3828 = n5019 ^ n5020;
  assign n4991 = n5020 & n5019;
  assign n5044 = n5022 & n156;
  assign n5040 = ~n5058;
  assign n5042 = ~n5022;
  assign n5069 = ~n5081;
  assign n5082 = n5096 & n5046;
  assign n5028 = ~n5097;
  assign n5090 = n844 & n5101;
  assign n927 = ~n844;
  assign n5119 = ~n5124;
  assign n3826 = ~n3828;
  assign n4994 = ~n4991;
  assign n5021 = n5040 & n5041;
  assign n5033 = n5042 & n5043;
  assign n5008 = ~n5044;
  assign n5045 = n5069 & n5070;
  assign n5048 = ~n5082;
  assign n3805 = ~n5090;
  assign n5080 = n927 & n5091;
  assign n5071 = n927 & n3639;
  assign n5098 = n5119 & n5120;
  assign n2773 = n3826 ^ n2728;
  assign n3861 = n3826 & n2728;
  assign n5006 = n5021 ^ n5022;
  assign n5023 = ~n5021;
  assign n5024 = ~n5033;
  assign n5025 = n5045 ^ n5046;
  assign n5047 = ~n5045;
  assign n5000 = n5071 ^ n2262;
  assign n3844 = ~n5080;
  assign n5072 = n5098 ^ n2194;
  assign n5100 = n5098 & n5076;
  assign n5099 = ~n5098;
  assign n4990 = n3861 & n2695;
  assign n78252 = ~n2773;
  assign n3845 = ~n3861;
  assign n4992 = n156 ^ n5006;
  assign n5018 = n5023 & n5024;
  assign n4996 = n5025 ^ n5026;
  assign n5034 = n5047 & n5048;
  assign n5051 = n5000 & n5013;
  assign n5049 = ~n5000;
  assign n5059 = n3844 & n3805;
  assign n785 = n5072 ^ n5073;
  assign n5083 = n5099 & n5078;
  assign n5077 = ~n5100;
  assign n4969 = n78252 & n3807;
  assign n4988 = n3845 & n2697;
  assign n4956 = ~n4990;
  assign n4975 = n4991 ^ n4992;
  assign n4993 = ~n4992;
  assign n5011 = n4996 & n155;
  assign n5007 = ~n5018;
  assign n5009 = ~n4996;
  assign n5027 = ~n5034;
  assign n5035 = n5049 & n5050;
  assign n5015 = ~n5051;
  assign n5039 = n785 & n5055;
  assign n3842 = ~n5059;
  assign n817 = ~n785;
  assign n5074 = n5077 & n5078;
  assign n5075 = ~n5083;
  assign n4952 = n4969 ^ n4970;
  assign n4949 = n4969 ^ n4971;
  assign n4954 = n4975 ^ n3845;
  assign n4976 = ~n4988;
  assign n4957 = n4993 & n4994;
  assign n4995 = n5007 & n5008;
  assign n5004 = n5009 & n5010;
  assign n4979 = ~n5011;
  assign n5012 = n5027 & n5028;
  assign n5002 = ~n5035;
  assign n5032 = n817 & n5038;
  assign n3729 = ~n5039;
  assign n5029 = n817 & n3557;
  assign n5056 = ~n5074;
  assign n5060 = n5075 & n5076;
  assign n3328 = n359 ^ n4949;
  assign n4933 = n4952 & n4953;
  assign n3779 = n2695 ^ n4954;
  assign n4950 = ~n4949;
  assign n4972 = n4976 & n4975;
  assign n4966 = ~n4957;
  assign n4977 = n4995 ^ n4996;
  assign n4997 = ~n4995;
  assign n4998 = ~n5004;
  assign n4999 = n5012 ^ n5013;
  assign n5014 = ~n5012;
  assign n4964 = n5029 ^ n2182;
  assign n3766 = ~n5032;
  assign n5054 = n5056 & n5057;
  assign n5052 = ~n5060;
  assign n4904 = n4933 ^ n4934;
  assign n4921 = n3779 & n3710;
  assign n4937 = n4933 & n4934;
  assign n4615 = ~n3328;
  assign n4935 = ~n4933;
  assign n4890 = n4950 & n359;
  assign n2638 = ~n3779;
  assign n4955 = ~n4972;
  assign n4958 = n155 ^ n4977;
  assign n4989 = n4997 & n4998;
  assign n4960 = n4999 ^ n5000;
  assign n5005 = n5014 & n5015;
  assign n4968 = ~n4964;
  assign n5017 = n3766 & n3729;
  assign n5036 = n5052 & n5053;
  assign n5031 = ~n5054;
  assign n4903 = n4921 ^ n2697;
  assign n78251 = n2638 ^ n2773;
  assign n4929 = n4935 & n4936;
  assign n3910 = n2638 & n2773;
  assign n4899 = ~n4937;
  assign n4930 = n4890 & n358;
  assign n4927 = ~n4890;
  assign n4938 = n4955 & n4956;
  assign n4924 = n4957 ^ n4958;
  assign n4914 = n4958 & n4966;
  assign n4980 = n4960 & n4987;
  assign n4978 = ~n4989;
  assign n4981 = ~n4960;
  assign n5001 = ~n5005;
  assign n3764 = ~n5017;
  assign n5030 = ~n5036;
  assign n4891 = n4903 ^ n4904;
  assign n4922 = n4927 & n4928;
  assign n4910 = ~n4929;
  assign n4877 = ~n4930;
  assign n4912 = n4938 ^ n4924;
  assign n4940 = n4938 & n2529;
  assign n4939 = ~n4938;
  assign n4959 = n4978 & n4979;
  assign n4962 = ~n4980;
  assign n4973 = n4981 & n154;
  assign n4982 = n5001 & n5002;
  assign n726 = n5030 & n5031;
  assign n4871 = n4890 ^ n4891;
  assign n4905 = n4910 & n4903;
  assign n3693 = n2536 ^ n4912;
  assign n4897 = ~n4922;
  assign n4931 = n4939 & n2536;
  assign n4923 = ~n4940;
  assign n4941 = n4959 ^ n4960;
  assign n4961 = ~n4959;
  assign n4943 = ~n4973;
  assign n4963 = n4982 ^ n4983;
  assign n4986 = n4982 & n4983;
  assign n4984 = ~n4982;
  assign n5003 = n726 & n5016;
  assign n2184 = ~n726;
  assign n4857 = n358 ^ n4871;
  assign n4892 = n4891 & n4897;
  assign n4898 = ~n4905;
  assign n4893 = n3693 & n3674;
  assign n2598 = ~n3693;
  assign n4913 = n4923 & n4924;
  assign n4907 = ~n4931;
  assign n4915 = n154 ^ n4941;
  assign n4951 = n4961 & n4962;
  assign n4918 = n4963 ^ n4964;
  assign n4974 = n4984 & n4985;
  assign n4967 = ~n4986;
  assign n4908 = n5003 ^ n1998;
  assign n3265 = n4857 ^ n3328;
  assign n4815 = n4857 & n4615;
  assign n4876 = ~n4892;
  assign n4861 = n4893 ^ n2536;
  assign n4878 = n4898 & n4899;
  assign n78250 = n3910 ^ n2598;
  assign n4859 = n2598 & n3910;
  assign n4906 = ~n4913;
  assign n4873 = n4914 ^ n4915;
  assign n4916 = ~n4915;
  assign n4944 = n4918 & n4946;
  assign n4942 = ~n4951;
  assign n4945 = ~n4918;
  assign n4965 = n4967 & n4968;
  assign n4948 = ~n4974;
  assign n4583 = ~n3265;
  assign n4818 = ~n4815;
  assign n4845 = n4876 & n4877;
  assign n4860 = n4878 ^ n4879;
  assign n4882 = n4878 & n4879;
  assign n4869 = ~n4861;
  assign n4880 = ~n4878;
  assign n4894 = n4906 & n4907;
  assign n4885 = n4916 & n4914;
  assign n4917 = n4942 & n4943;
  assign n4920 = ~n4944;
  assign n4932 = n4945 & n153;
  assign n4947 = ~n4965;
  assign n4846 = n4860 ^ n4861;
  assign n4863 = n4845 & n4867;
  assign n4862 = ~n4845;
  assign n4872 = n4880 & n4881;
  assign n4868 = ~n4882;
  assign n4874 = n4894 ^ n2410;
  assign n4896 = n4894 & n2410;
  assign n4895 = ~n4894;
  assign n4900 = n4917 ^ n4918;
  assign n4919 = ~n4917;
  assign n4902 = ~n4932;
  assign n4925 = n4947 & n4948;
  assign n4831 = n4845 ^ n4846;
  assign n4847 = ~n4846;
  assign n4858 = n4862 & n357;
  assign n4848 = ~n4863;
  assign n4864 = n4868 & n4869;
  assign n4854 = ~n4872;
  assign n2531 = n4873 ^ n4874;
  assign n4884 = n4895 & n2472;
  assign n4883 = ~n4896;
  assign n4886 = n153 ^ n4900;
  assign n4911 = n4919 & n4920;
  assign n4909 = n4925 ^ n4926;
  assign n4816 = n357 ^ n4831;
  assign n4842 = n4847 & n4848;
  assign n4833 = ~n4858;
  assign n78249 = n4859 ^ n2531;
  assign n4853 = ~n4864;
  assign n4823 = n2531 & n4859;
  assign n3713 = ~n2531;
  assign n4875 = n4883 & n4873;
  assign n4866 = ~n4884;
  assign n4836 = n4885 ^ n4886;
  assign n4887 = ~n4886;
  assign n4889 = n4908 ^ n4909;
  assign n4901 = ~n4911;
  assign n4538 = n4815 ^ n4816;
  assign n4817 = ~n4816;
  assign n4832 = ~n4842;
  assign n4849 = n4853 & n4854;
  assign n4843 = n3713 & n3574;
  assign n4865 = ~n4875;
  assign n4855 = n4887 & n4885;
  assign n4888 = n4901 & n4902;
  assign n4546 = ~n4538;
  assign n4775 = n4817 & n4818;
  assign n4802 = n4832 & n4833;
  assign n4822 = n4843 ^ n2410;
  assign n4814 = ~n4849;
  assign n4850 = n4865 & n4866;
  assign n4870 = n4888 ^ n4889;
  assign n4778 = ~n4775;
  assign n4820 = n4802 & n4824;
  assign n4819 = ~n4802;
  assign n4821 = n4814 ^ n4834;
  assign n4828 = n4822 & n4834;
  assign n4829 = ~n4822;
  assign n4835 = n4850 ^ n2355;
  assign n4852 = n4850 & n2355;
  assign n4851 = ~n4850;
  assign n4856 = n152 ^ n4870;
  assign n4812 = n4819 & n356;
  assign n4807 = ~n4820;
  assign n4803 = n4821 ^ n4822;
  assign n4801 = ~n4828;
  assign n4825 = n4829 & n4830;
  assign n2433 = n4835 ^ n4836;
  assign n4844 = n4851 & n2365;
  assign n4839 = ~n4852;
  assign n4796 = n4855 ^ n4856;
  assign n4789 = n4802 ^ n4803;
  assign n4804 = n4803 & n4807;
  assign n4793 = ~n4812;
  assign n78248 = n4823 ^ n2433;
  assign n4787 = n2433 & n4823;
  assign n4813 = ~n4825;
  assign n3662 = ~n2433;
  assign n4837 = n4839 & n4836;
  assign n4827 = ~n4844;
  assign n4841 = n4796 & n2188;
  assign n4840 = ~n4796;
  assign n4776 = n356 ^ n4789;
  assign n4792 = ~n4804;
  assign n4808 = n4813 & n4814;
  assign n4805 = n3662 & n3510;
  assign n4826 = ~n4837;
  assign n4838 = n4840 & n2295;
  assign n4811 = ~n4841;
  assign n3209 = n4775 ^ n4776;
  assign n4777 = ~n4776;
  assign n4753 = n4792 & n4793;
  assign n4767 = n4805 ^ n2365;
  assign n4800 = ~n4808;
  assign n4809 = n4826 & n4827;
  assign n4799 = ~n4838;
  assign n4504 = ~n3209;
  assign n4723 = n4777 & n4778;
  assign n4745 = ~n4753;
  assign n4791 = n4767 & n4794;
  assign n4795 = n4800 & n4801;
  assign n4790 = ~n4767;
  assign n4797 = n4809 ^ n2295;
  assign n4810 = ~n4809;
  assign n4726 = ~n4723;
  assign n4788 = n4790 & n4783;
  assign n4781 = ~n4791;
  assign n4782 = ~n4795;
  assign n2383 = n4796 ^ n4797;
  assign n4806 = n4810 & n4811;
  assign n4779 = n4781 & n4782;
  assign n4766 = n4782 ^ n4783;
  assign n78247 = n4787 ^ n2383;
  assign n4761 = n2383 & n4787;
  assign n4769 = ~n4788;
  assign n3565 = ~n2383;
  assign n4798 = ~n4806;
  assign n4754 = n4766 ^ n4767;
  assign n4768 = ~n4779;
  assign n4770 = n3565 & n3450;
  assign n4784 = n4798 & n4799;
  assign n4738 = n4753 ^ n4754;
  assign n4755 = n4754 & n4762;
  assign n4756 = ~n4754;
  assign n4765 = n4768 & n4769;
  assign n4736 = n4770 ^ n2295;
  assign n4772 = n4784 ^ n2207;
  assign n4785 = ~n4784;
  assign n4724 = n355 ^ n4738;
  assign n4744 = ~n4755;
  assign n4749 = n4756 & n355;
  assign n4757 = n4736 & n4763;
  assign n4747 = ~n4765;
  assign n4758 = ~n4736;
  assign n2281 = n4771 ^ n4772;
  assign n4780 = n4785 & n4786;
  assign n4451 = n4723 ^ n4724;
  assign n4725 = ~n4724;
  assign n4739 = n4744 & n4745;
  assign n4730 = ~n4749;
  assign n4735 = n4747 ^ n4750;
  assign n4746 = ~n4757;
  assign n4751 = n4758 & n4750;
  assign n78246 = n4761 ^ n2281;
  assign n4704 = n2281 & n4761;
  assign n3537 = ~n2281;
  assign n4773 = ~n4780;
  assign n3155 = ~n4451;
  assign n4675 = n4725 & n4726;
  assign n4707 = n4735 ^ n4736;
  assign n4729 = ~n4739;
  assign n4740 = n4746 & n4747;
  assign n4732 = ~n4751;
  assign n4741 = n3537 & n3401;
  assign n4764 = n4773 & n4774;
  assign n4719 = n4707 & n4727;
  assign n4728 = n4729 & n4730;
  assign n4720 = ~n4707;
  assign n4731 = ~n4740;
  assign n4696 = n4741 ^ n2207;
  assign n4760 = n4764 & n2130;
  assign n4759 = ~n4764;
  assign n4705 = ~n4719;
  assign n4710 = n4720 & n354;
  assign n4706 = ~n4728;
  assign n4711 = n4731 & n4732;
  assign n4752 = n4759 & n2151;
  assign n4743 = ~n4760;
  assign n4702 = n4705 & n4706;
  assign n4692 = n4706 ^ n4707;
  assign n4694 = ~n4710;
  assign n4695 = n4711 ^ n4712;
  assign n4715 = n4711 & n4712;
  assign n4713 = ~n4711;
  assign n4742 = n4743 & n4748;
  assign n4734 = ~n4752;
  assign n4676 = n354 ^ n4692;
  assign n4678 = n4695 ^ n4696;
  assign n4693 = ~n4702;
  assign n4708 = n4713 & n4714;
  assign n4703 = ~n4715;
  assign n4733 = ~n4742;
  assign n4737 = n4734 & n4743;
  assign n4408 = n4675 ^ n4676;
  assign n4637 = n4676 & n4675;
  assign n4684 = n4678 & n353;
  assign n4677 = n4693 & n4694;
  assign n4682 = ~n4678;
  assign n4697 = n4703 & n4696;
  assign n4690 = ~n4708;
  assign n4716 = n4733 & n4734;
  assign n4722 = ~n4737;
  assign n4417 = ~n4408;
  assign n4640 = ~n4637;
  assign n4659 = n4677 ^ n4678;
  assign n4679 = n4682 & n4683;
  assign n4647 = ~n4684;
  assign n4663 = ~n4677;
  assign n4689 = ~n4697;
  assign n4698 = n4716 ^ n2039;
  assign n2212 = n4721 ^ n4722;
  assign n4717 = ~n4716;
  assign n4638 = n353 ^ n4659;
  assign n4662 = ~n4679;
  assign n4670 = n4689 & n4690;
  assign n2112 = n4698 ^ n4699;
  assign n78245 = n4704 ^ n2212;
  assign n4681 = n2212 & n4704;
  assign n4709 = n4717 & n4718;
  assign n3473 = ~n2212;
  assign n3066 = n4637 ^ n4638;
  assign n4639 = ~n4638;
  assign n4660 = n4662 & n4663;
  assign n4657 = n4670 ^ n4671;
  assign n4674 = n4670 & n4671;
  assign n4672 = ~n4670;
  assign n3417 = ~n2112;
  assign n4685 = ~n4681;
  assign n4691 = n3473 & n3369;
  assign n4700 = ~n4709;
  assign n4390 = ~n3066;
  assign n4584 = n4639 & n4640;
  assign n4646 = ~n4660;
  assign n4664 = n4672 & n4673;
  assign n4661 = ~n4674;
  assign n78260 = n4681 ^ n3417;
  assign n4651 = n3417 & n4685;
  assign n4665 = n3417 & n3321;
  assign n4656 = n4691 ^ n2130;
  assign n4686 = n4700 & n4701;
  assign n4641 = n4646 & n4647;
  assign n4624 = n4656 ^ n4657;
  assign n4658 = n4661 & n4656;
  assign n4643 = ~n4664;
  assign n4603 = n4665 ^ n2039;
  assign n4666 = n4686 ^ n1976;
  assign n4687 = ~n4686;
  assign n4636 = n4624 & n352;
  assign n4621 = ~n4641;
  assign n4634 = ~n4624;
  assign n4642 = ~n4658;
  assign n4650 = n4603 & n4626;
  assign n4648 = ~n4603;
  assign n2042 = n4666 ^ n4667;
  assign n4680 = n4687 & n4688;
  assign n4601 = n4621 ^ n4624;
  assign n4629 = n4634 & n4635;
  assign n4600 = ~n4636;
  assign n4625 = n4642 & n4643;
  assign n4644 = n4648 & n4649;
  assign n4605 = ~n4650;
  assign n78259 = n4651 ^ n2042;
  assign n3374 = ~n2042;
  assign n4668 = ~n4680;
  assign n4585 = n352 ^ n4601;
  assign n4602 = n4625 ^ n4626;
  assign n4620 = ~n4629;
  assign n4627 = ~n4625;
  assign n4628 = ~n4644;
  assign n4609 = n3374 & n4651;
  assign n4630 = n3374 & n3278;
  assign n4652 = n4668 & n4669;
  assign n4329 = n4584 ^ n4585;
  assign n4528 = n4585 & n4584;
  assign n4571 = n4602 ^ n4603;
  assign n4611 = n4620 & n4621;
  assign n4622 = n4627 & n4628;
  assign n4563 = n4630 ^ n1979;
  assign n4623 = ~n4609;
  assign n4631 = n4652 ^ n4653;
  assign n4654 = ~n4652;
  assign n4321 = ~n4329;
  assign n4586 = n4571 & n4592;
  assign n4587 = ~n4571;
  assign n4599 = ~n4611;
  assign n4604 = ~n4622;
  assign n4614 = n4563 & n4589;
  assign n4612 = ~n4563;
  assign n1981 = n1927 ^ n4631;
  assign n4645 = n4654 & n4655;
  assign n4569 = ~n4586;
  assign n4580 = n4587 & n367;
  assign n4593 = n4599 & n4600;
  assign n4588 = n4604 & n4605;
  assign n4606 = n4612 & n4613;
  assign n4591 = ~n4614;
  assign n4579 = n1981 & n4623;
  assign n4616 = n1981 & n3328;
  assign n4610 = ~n1981;
  assign n4632 = ~n4645;
  assign n4555 = ~n4580;
  assign n4562 = n4588 ^ n4589;
  assign n4570 = ~n4593;
  assign n4590 = ~n4588;
  assign n4565 = ~n4606;
  assign n78258 = n4609 ^ n4610;
  assign n4594 = n4610 & n3223;
  assign n4607 = n4610 & n4615;
  assign n3308 = ~n4616;
  assign n4617 = n4632 & n4633;
  assign n4532 = n4562 ^ n4563;
  assign n4561 = n4569 & n4570;
  assign n4553 = n4570 ^ n4571;
  assign n4581 = n4590 & n4591;
  assign n4521 = n4594 ^ n1917;
  assign n3330 = ~n4607;
  assign n4596 = n4617 ^ n1840;
  assign n4618 = ~n4617;
  assign n4529 = n367 ^ n4553;
  assign n4547 = n4532 & n4556;
  assign n4548 = ~n4532;
  assign n4554 = ~n4561;
  assign n4564 = ~n4581;
  assign n4572 = n4521 & n4582;
  assign n4573 = ~n4521;
  assign n1912 = n4595 ^ n4596;
  assign n4608 = n4618 & n4619;
  assign n2981 = n4528 ^ n4529;
  assign n4530 = ~n4529;
  assign n4534 = ~n4547;
  assign n4544 = n4548 & n366;
  assign n4531 = n4554 & n4555;
  assign n4549 = n4564 & n4565;
  assign n4524 = ~n4572;
  assign n4566 = n4573 & n4550;
  assign n78257 = n4579 ^ n1912;
  assign n4543 = n1912 & n4579;
  assign n4574 = n1912 & n4583;
  assign n3288 = ~n1912;
  assign n4597 = ~n4608;
  assign n4283 = ~n2981;
  assign n4487 = n4530 & n4528;
  assign n4512 = n4531 ^ n4532;
  assign n4514 = ~n4544;
  assign n4533 = ~n4531;
  assign n4522 = n4549 ^ n4550;
  assign n4551 = ~n4549;
  assign n4552 = ~n4566;
  assign n4557 = n3288 & n3171;
  assign n4567 = n3288 & n3265;
  assign n3267 = ~n4574;
  assign n4575 = n4597 & n4598;
  assign n4488 = n366 ^ n4512;
  assign n4490 = ~n4487;
  assign n4492 = n4521 ^ n4522;
  assign n4520 = n4533 & n4534;
  assign n4545 = n4551 & n4552;
  assign n4480 = n4557 ^ n1867;
  assign n3290 = ~n4567;
  assign n4558 = n4575 ^ n4576;
  assign n4577 = ~n4575;
  assign n2940 = n4487 ^ n4488;
  assign n4489 = ~n4488;
  assign n4507 = n4492 & n365;
  assign n4505 = ~n4492;
  assign n4513 = ~n4520;
  assign n4523 = ~n4545;
  assign n4537 = n4480 & n4509;
  assign n4535 = ~n4480;
  assign n1853 = n4558 ^ n1825;
  assign n4568 = n4577 & n4578;
  assign n4252 = ~n2940;
  assign n4446 = n4489 & n4490;
  assign n4501 = n4505 & n4506;
  assign n4462 = ~n4507;
  assign n4491 = n4513 & n4514;
  assign n4508 = n4523 & n4524;
  assign n4525 = n4535 & n4536;
  assign n4511 = ~n4537;
  assign n78256 = n4543 ^ n1853;
  assign n4500 = n1853 & n4543;
  assign n4539 = n1853 & n4546;
  assign n3217 = ~n1853;
  assign n4559 = ~n4568;
  assign n4449 = ~n4446;
  assign n4470 = n4491 ^ n4492;
  assign n4479 = ~n4501;
  assign n4478 = ~n4491;
  assign n4481 = n4508 ^ n4509;
  assign n4510 = ~n4508;
  assign n4483 = ~n4525;
  assign n4503 = ~n4500;
  assign n4515 = n3217 & n3152;
  assign n4526 = n3217 & n4538;
  assign n3232 = ~n4539;
  assign n4540 = n4559 & n4560;
  assign n4447 = n365 ^ n4470;
  assign n4476 = n4478 & n4479;
  assign n4435 = n4480 ^ n4481;
  assign n4502 = n4510 & n4511;
  assign n4439 = n4515 ^ n1812;
  assign n3251 = ~n4526;
  assign n4517 = n4540 ^ n1752;
  assign n4541 = ~n4540;
  assign n2923 = n4446 ^ n4447;
  assign n4448 = ~n4447;
  assign n4463 = n4435 & n4471;
  assign n4461 = ~n4476;
  assign n4464 = ~n4435;
  assign n4482 = ~n4502;
  assign n4493 = n4439 & n4466;
  assign n4494 = ~n4439;
  assign n3248 = n3251 & n3232;
  assign n3162 = n4516 ^ n4517;
  assign n4527 = n4541 & n4542;
  assign n4206 = ~n2923;
  assign n4391 = n4448 & n4449;
  assign n4434 = n4461 & n4462;
  assign n4437 = ~n4463;
  assign n4456 = n4464 & n364;
  assign n4465 = n4482 & n4483;
  assign n4441 = ~n4493;
  assign n4484 = n4494 & n4495;
  assign n78255 = n4500 ^ n3162;
  assign n4444 = n3162 & n4503;
  assign n4477 = n3162 & n3096;
  assign n4496 = n3162 & n4504;
  assign n1826 = ~n3162;
  assign n4518 = ~n4527;
  assign n4418 = n4434 ^ n4435;
  assign n4436 = ~n4434;
  assign n4420 = ~n4456;
  assign n4438 = n4465 ^ n4466;
  assign n4467 = ~n4465;
  assign n4398 = n4477 ^ n1752;
  assign n4468 = ~n4484;
  assign n4460 = ~n4444;
  assign n3211 = ~n4496;
  assign n4485 = n1826 & n3209;
  assign n4497 = n4518 & n4519;
  assign n4392 = n364 ^ n4418;
  assign n4433 = n4436 & n4437;
  assign n4394 = n4438 ^ n4439;
  assign n4457 = n4467 & n4468;
  assign n4458 = n4398 & n4469;
  assign n4459 = ~n4398;
  assign n3195 = ~n4485;
  assign n4473 = n4497 ^ n1687;
  assign n4498 = ~n4497;
  assign n2861 = n4391 ^ n4392;
  assign n4347 = n4392 & n4391;
  assign n4421 = n4394 & n4427;
  assign n4419 = ~n4433;
  assign n4422 = ~n4394;
  assign n4440 = ~n4457;
  assign n4400 = ~n4458;
  assign n4450 = n4459 & n4424;
  assign n1785 = n4472 ^ n4473;
  assign n4486 = n4498 & n4499;
  assign n4163 = ~n2861;
  assign n4350 = ~n4347;
  assign n4393 = n4419 & n4420;
  assign n4396 = ~n4421;
  assign n4414 = n4422 & n363;
  assign n4423 = n4440 & n4441;
  assign n4426 = ~n4450;
  assign n4413 = n1785 & n4460;
  assign n4452 = n1785 & n3155;
  assign n4445 = ~n1785;
  assign n4474 = ~n4486;
  assign n4372 = n4393 ^ n4394;
  assign n4395 = ~n4393;
  assign n4374 = ~n4414;
  assign n4397 = n4423 ^ n4424;
  assign n4425 = ~n4423;
  assign n78254 = n4444 ^ n4445;
  assign n4428 = n4445 & n3100;
  assign n4442 = n4445 & n4451;
  assign n3158 = ~n4452;
  assign n4453 = n4474 & n4475;
  assign n4348 = n363 ^ n4372;
  assign n4388 = n4395 & n4396;
  assign n4352 = n4397 ^ n4398;
  assign n4415 = n4425 & n4426;
  assign n4356 = n4428 ^ n1687;
  assign n3179 = ~n4442;
  assign n4429 = n4453 ^ n1722;
  assign n4454 = ~n4453;
  assign n4143 = n4347 ^ n4348;
  assign n4349 = ~n4348;
  assign n4377 = n4352 & n362;
  assign n4373 = ~n4388;
  assign n4375 = ~n4352;
  assign n4399 = ~n4415;
  assign n4405 = n4356 & n4416;
  assign n4404 = ~n4356;
  assign n1756 = n4429 ^ n4430;
  assign n4443 = n4454 & n4455;
  assign n4134 = ~n4143;
  assign n4307 = n4349 & n4350;
  assign n4351 = n4373 & n4374;
  assign n4368 = n4375 & n4376;
  assign n4332 = ~n4377;
  assign n4378 = n4399 & n4400;
  assign n4401 = n4404 & n4379;
  assign n4358 = ~n4405;
  assign n78253 = n4413 ^ n1756;
  assign n4387 = n1756 & n4413;
  assign n4407 = n1756 & n4417;
  assign n4406 = ~n1756;
  assign n4431 = ~n4443;
  assign n4330 = n4351 ^ n4352;
  assign n4353 = ~n4351;
  assign n4354 = ~n4368;
  assign n4355 = n4378 ^ n4379;
  assign n4380 = ~n4378;
  assign n4381 = ~n4401;
  assign n4389 = ~n4387;
  assign n4383 = n4406 & n3078;
  assign n3115 = ~n4407;
  assign n4402 = n4406 & n4408;
  assign n4410 = n4431 & n4432;
  assign n4308 = n362 ^ n4330;
  assign n4344 = n4353 & n4354;
  assign n4310 = n4355 ^ n4356;
  assign n4369 = n4380 & n4381;
  assign n4314 = n4383 ^ n1667;
  assign n3138 = ~n4402;
  assign n3023 = n4409 ^ n4410;
  assign n4411 = ~n4410;
  assign n4085 = n4307 ^ n4308;
  assign n4267 = n4308 & n4307;
  assign n4335 = n4310 & n361;
  assign n4331 = ~n4344;
  assign n4333 = ~n4310;
  assign n4357 = ~n4369;
  assign n4363 = n4314 & n4370;
  assign n4362 = ~n4314;
  assign n3135 = n3138 & n3115;
  assign n78268 = n4387 ^ n3023;
  assign n4319 = n3023 & n4389;
  assign n4371 = n3023 & n3013;
  assign n4384 = n3023 & n4390;
  assign n1723 = ~n3023;
  assign n4403 = n4411 & n4412;
  assign n4094 = ~n4085;
  assign n4309 = n4331 & n4332;
  assign n4326 = n4333 & n4334;
  assign n4293 = ~n4335;
  assign n4336 = n4357 & n4358;
  assign n4360 = n4362 & n4337;
  assign n4316 = ~n4363;
  assign n4276 = n4371 ^ n1684;
  assign n4328 = ~n4319;
  assign n4382 = n1723 & n3066;
  assign n3091 = ~n4384;
  assign n4385 = ~n4403;
  assign n4291 = n4309 ^ n4310;
  assign n4311 = ~n4309;
  assign n4312 = ~n4326;
  assign n4313 = n4336 ^ n4337;
  assign n4338 = ~n4336;
  assign n4345 = n4276 & n4359;
  assign n4339 = ~n4360;
  assign n4346 = ~n4276;
  assign n3069 = ~n4382;
  assign n4364 = n4385 & n4386;
  assign n4271 = n361 ^ n4291;
  assign n4306 = n4311 & n4312;
  assign n4273 = n4313 ^ n4314;
  assign n4327 = n4338 & n4339;
  assign n4279 = ~n4345;
  assign n4340 = n4346 & n4298;
  assign n4341 = n4364 ^ n4365;
  assign n4366 = ~n4364;
  assign n4007 = n4267 ^ n4271;
  assign n4229 = n4271 & n4267;
  assign n4268 = ~n4271;
  assign n4296 = n4273 & n360;
  assign n4292 = ~n4306;
  assign n4294 = ~n4273;
  assign n4315 = ~n4327;
  assign n4300 = ~n4340;
  assign n1659 = n4341 ^ n1528;
  assign n4361 = n4366 & n4367;
  assign n4002 = n4267 ^ n4268;
  assign n4272 = n4292 & n4293;
  assign n4288 = n4294 & n4295;
  assign n4255 = ~n4296;
  assign n4297 = n4315 & n4316;
  assign n4287 = n1659 & n4328;
  assign n4322 = n1659 & n4329;
  assign n4320 = ~n1659;
  assign n4342 = ~n4361;
  assign n4253 = n4272 ^ n4273;
  assign n4274 = ~n4272;
  assign n4275 = ~n4288;
  assign n4277 = n4297 ^ n4298;
  assign n4299 = ~n4297;
  assign n78267 = n4319 ^ n4320;
  assign n4290 = ~n4287;
  assign n4301 = n4320 & n2992;
  assign n4317 = n4320 & n4321;
  assign n3028 = ~n4322;
  assign n4323 = n4342 & n4343;
  assign n4230 = n360 ^ n4253;
  assign n4269 = n4274 & n4275;
  assign n4213 = n4276 ^ n4277;
  assign n4289 = n4299 & n4300;
  assign n4240 = n4301 ^ n1608;
  assign n3053 = ~n4317;
  assign n4303 = n4323 ^ n1499;
  assign n4324 = ~n4323;
  assign n3977 = n4229 ^ n4230;
  assign n4185 = n4230 & n4229;
  assign n4258 = n4213 & n375;
  assign n4254 = ~n4269;
  assign n4256 = ~n4213;
  assign n4278 = ~n4289;
  assign n3050 = n3053 & n3028;
  assign n3006 = n4302 ^ n4303;
  assign n4318 = n4324 & n4325;
  assign n3984 = ~n3977;
  assign n4188 = ~n4185;
  assign n4231 = n4254 & n4255;
  assign n4246 = n4256 & n4257;
  assign n4215 = ~n4258;
  assign n4259 = n4278 & n4279;
  assign n78266 = n4287 ^ n3006;
  assign n4227 = n3006 & n4290;
  assign n4270 = n3006 & n2932;
  assign n4282 = n3006 & n2981;
  assign n1610 = ~n3006;
  assign n4304 = ~n4318;
  assign n4212 = n375 ^ n4231;
  assign n4232 = ~n4231;
  assign n4233 = ~n4246;
  assign n4234 = n4259 ^ n4240;
  assign n4261 = n4259 & n4262;
  assign n4260 = ~n4259;
  assign n4175 = n4270 ^ n1551;
  assign n4251 = ~n4227;
  assign n3008 = ~n4282;
  assign n4280 = n1610 & n4283;
  assign n4284 = n4304 & n4305;
  assign n4186 = n4212 ^ n4213;
  assign n4226 = n4232 & n4233;
  assign n4190 = n4234 ^ n4235;
  assign n4247 = n4260 & n4235;
  assign n4250 = n4175 & n4198;
  assign n4239 = ~n4261;
  assign n4248 = ~n4175;
  assign n2984 = ~n4280;
  assign n4263 = n4284 ^ n1513;
  assign n4285 = ~n4284;
  assign n2600 = n4185 ^ n4186;
  assign n4187 = ~n4186;
  assign n4216 = n4190 & n4218;
  assign n4214 = ~n4226;
  assign n4217 = ~n4190;
  assign n4236 = n4239 & n4240;
  assign n4220 = ~n4247;
  assign n4241 = n4248 & n4249;
  assign n4200 = ~n4250;
  assign n1583 = n4263 ^ n4264;
  assign n4281 = n4285 & n4286;
  assign n3935 = ~n2600;
  assign n4151 = n4187 & n4188;
  assign n4189 = n4214 & n4215;
  assign n4192 = ~n4216;
  assign n4211 = n4217 & n374;
  assign n4219 = ~n4236;
  assign n4178 = ~n4241;
  assign n4210 = n1583 & n4251;
  assign n4242 = n1583 & n4252;
  assign n4228 = ~n1583;
  assign n4265 = ~n4281;
  assign n4145 = ~n4151;
  assign n4172 = n4189 ^ n4190;
  assign n4191 = ~n4189;
  assign n4174 = ~n4211;
  assign n4197 = n4219 & n4220;
  assign n78265 = n4227 ^ n4228;
  assign n4221 = n4228 & n2879;
  assign n4237 = n4228 & n2940;
  assign n2943 = ~n4242;
  assign n4243 = n4265 & n4266;
  assign n4152 = n374 ^ n4172;
  assign n4184 = n4191 & n4192;
  assign n4176 = n4197 ^ n4198;
  assign n4199 = ~n4197;
  assign n4129 = n4221 ^ n1523;
  assign n2968 = ~n4237;
  assign n4222 = n4243 ^ n1471;
  assign n4244 = ~n4243;
  assign n3890 = n4151 ^ n4152;
  assign n4144 = ~n4152;
  assign n4141 = n4175 ^ n4176;
  assign n4173 = ~n4184;
  assign n4193 = n4199 & n4200;
  assign n4203 = n4129 & n4156;
  assign n4201 = ~n4129;
  assign n1515 = n4222 ^ n4223;
  assign n4238 = n4244 & n4245;
  assign n2572 = ~n3890;
  assign n4095 = n4144 & n4145;
  assign n4153 = n4141 & n4169;
  assign n4170 = n4173 & n4174;
  assign n4154 = ~n4141;
  assign n4177 = ~n4193;
  assign n4194 = n4201 & n4202;
  assign n4158 = ~n4203;
  assign n78264 = n4210 ^ n1515;
  assign n4168 = n1515 & n4210;
  assign n4205 = n1515 & n2923;
  assign n4204 = ~n1515;
  assign n4224 = ~n4238;
  assign n4098 = ~n4095;
  assign n4139 = ~n4153;
  assign n4146 = n4154 & n373;
  assign n4140 = ~n4170;
  assign n4155 = n4177 & n4178;
  assign n4131 = ~n4194;
  assign n4179 = n4204 & n2850;
  assign n2904 = ~n4205;
  assign n4195 = n4204 & n4206;
  assign n4207 = n4224 & n4225;
  assign n4127 = n4139 & n4140;
  assign n4123 = n4140 ^ n4141;
  assign n4125 = ~n4146;
  assign n4128 = n4155 ^ n4156;
  assign n4157 = ~n4155;
  assign n4089 = n4179 ^ n1456;
  assign n2925 = ~n4195;
  assign n4181 = n4207 ^ n1362;
  assign n4208 = ~n4207;
  assign n4096 = n373 ^ n4123;
  assign n4124 = ~n4127;
  assign n4100 = n4128 ^ n4129;
  assign n4147 = n4157 & n4158;
  assign n4160 = n4089 & n4171;
  assign n4159 = ~n4089;
  assign n1415 = n4180 ^ n4181;
  assign n4196 = n4208 & n4209;
  assign n3853 = n4095 ^ n4096;
  assign n4097 = ~n4096;
  assign n4108 = n4100 & n4120;
  assign n4099 = n4124 & n4125;
  assign n4109 = ~n4100;
  assign n4130 = ~n4147;
  assign n4148 = n4159 & n4111;
  assign n4082 = ~n4160;
  assign n78263 = n4168 ^ n1415;
  assign n4137 = n1415 & n4168;
  assign n4162 = n1415 & n2861;
  assign n4161 = ~n1415;
  assign n4182 = ~n4196;
  assign n3840 = ~n3853;
  assign n4056 = n4097 & n4098;
  assign n4074 = n4099 ^ n4100;
  assign n4101 = ~n4108;
  assign n4103 = n4109 & n372;
  assign n4102 = ~n4099;
  assign n4110 = n4130 & n4131;
  assign n4113 = ~n4148;
  assign n4142 = ~n4137;
  assign n4132 = n4161 & n2709;
  assign n2864 = ~n4162;
  assign n4149 = n4161 & n4163;
  assign n4165 = n4182 & n4183;
  assign n4057 = n372 ^ n4074;
  assign n4059 = ~n4056;
  assign n4088 = n4101 & n4102;
  assign n4076 = ~n4103;
  assign n4090 = n4110 ^ n4111;
  assign n4112 = ~n4110;
  assign n4051 = n4132 ^ n1362;
  assign n2886 = ~n4149;
  assign n4138 = n4164 ^ n4165;
  assign n4166 = ~n4165;
  assign n3803 = n4056 ^ n4057;
  assign n4058 = ~n4057;
  assign n4075 = ~n4088;
  assign n4077 = n4089 ^ n4090;
  assign n4104 = n4112 & n4113;
  assign n4114 = n4051 & n4121;
  assign n4115 = ~n4051;
  assign n78262 = n4137 ^ n4138;
  assign n4079 = n4138 & n4142;
  assign n4122 = n4138 & n2777;
  assign n4133 = n4138 & n4143;
  assign n1395 = ~n4138;
  assign n4150 = n4166 & n4167;
  assign n2417 = ~n3803;
  assign n4009 = n4058 & n4059;
  assign n4028 = n4075 & n4076;
  assign n4068 = n4077 & n371;
  assign n4066 = ~n4077;
  assign n4081 = ~n4104;
  assign n4053 = ~n4114;
  assign n4105 = n4115 & n4070;
  assign n4035 = n4122 ^ n1349;
  assign n4093 = ~n4079;
  assign n2842 = ~n4133;
  assign n4126 = n1395 & n4134;
  assign n4135 = ~n4150;
  assign n4048 = ~n4028;
  assign n4061 = n4066 & n4067;
  assign n4030 = ~n4068;
  assign n4069 = n4081 & n4082;
  assign n4072 = ~n4105;
  assign n4092 = n4035 & n4106;
  assign n4091 = ~n4035;
  assign n2814 = ~n4126;
  assign n4116 = n4135 & n4136;
  assign n4049 = ~n4061;
  assign n4050 = n4069 ^ n4070;
  assign n4071 = ~n4069;
  assign n4083 = n4091 & n4015;
  assign n4037 = ~n4092;
  assign n2839 = n2842 & n2814;
  assign n1320 = n4116 ^ n4117;
  assign n4118 = ~n4116;
  assign n4042 = n4048 & n4049;
  assign n4027 = n4049 & n4030;
  assign n3986 = n4050 ^ n4051;
  assign n4062 = n4071 & n4072;
  assign n4017 = ~n4083;
  assign n4004 = n1320 & n4093;
  assign n4084 = n1320 & n4094;
  assign n4080 = ~n1320;
  assign n4107 = n4118 & n4119;
  assign n4010 = n4027 ^ n4028;
  assign n4033 = n3986 & n370;
  assign n4029 = ~n4042;
  assign n4031 = ~n3986;
  assign n4052 = ~n4062;
  assign n78261 = n4079 ^ n4080;
  assign n4018 = ~n4004;
  assign n4063 = n4080 & n2724;
  assign n2771 = ~n4084;
  assign n4078 = n4080 & n4085;
  assign n4086 = ~n4107;
  assign n2332 = n4009 ^ n4010;
  assign n3954 = n4010 & n4009;
  assign n4011 = n4029 & n4030;
  assign n4025 = n4031 & n4032;
  assign n3988 = ~n4033;
  assign n4034 = n4052 & n4053;
  assign n4054 = n4063 ^ n1254;
  assign n2795 = ~n4078;
  assign n4073 = n4086 & n4087;
  assign n3738 = ~n2332;
  assign n3985 = n370 ^ n4011;
  assign n4012 = ~n4011;
  assign n4013 = ~n4025;
  assign n4014 = n4034 ^ n4035;
  assign n4036 = ~n4034;
  assign n4045 = n4054 & n4055;
  assign n4043 = ~n4054;
  assign n2792 = n2795 & n2771;
  assign n4065 = n4073 & n1223;
  assign n4064 = ~n4073;
  assign n3959 = n3985 ^ n3986;
  assign n4006 = n4012 & n4013;
  assign n3961 = n4014 ^ n4015;
  assign n4026 = n4036 & n4037;
  assign n4040 = n4043 & n4044;
  assign n3968 = ~n4045;
  assign n4060 = n4064 & n1228;
  assign n4047 = ~n4065;
  assign n3654 = n3954 ^ n3959;
  assign n3922 = n3959 & n3954;
  assign n3955 = ~n3959;
  assign n3991 = n3961 & n369;
  assign n3987 = ~n4006;
  assign n3989 = ~n3961;
  assign n4016 = ~n4026;
  assign n3995 = ~n4040;
  assign n4046 = n4047 & n4024;
  assign n4039 = ~n4060;
  assign n3641 = n3954 ^ n3955;
  assign n3925 = ~n3922;
  assign n3960 = n3987 & n3988;
  assign n3982 = n3989 & n3990;
  assign n3944 = ~n3991;
  assign n3992 = n4016 & n4017;
  assign n4022 = n3995 & n3968;
  assign n4038 = ~n4046;
  assign n4041 = n4039 & n4047;
  assign n3942 = n3960 ^ n3961;
  assign n3962 = ~n3960;
  assign n3963 = ~n3982;
  assign n3994 = ~n3992;
  assign n3993 = ~n4022;
  assign n4019 = n4038 & n4039;
  assign n4023 = ~n4041;
  assign n3923 = n369 ^ n3942;
  assign n3956 = n3962 & n3963;
  assign n3975 = n3992 ^ n3993;
  assign n3983 = n3994 & n3995;
  assign n3999 = n4019 ^ n1088;
  assign n4005 = n4023 ^ n4024;
  assign n4020 = ~n4019;
  assign n3903 = n3922 ^ n3923;
  assign n3924 = ~n3923;
  assign n3943 = ~n3956;
  assign n3966 = n3975 & n368;
  assign n3964 = ~n3975;
  assign n3967 = ~n3983;
  assign n1183 = n3998 ^ n3999;
  assign n78276 = n4004 ^ n4005;
  assign n3996 = n4005 & n2664;
  assign n4003 = n4005 & n4007;
  assign n3974 = n4005 & n4018;
  assign n4008 = n4020 & n4021;
  assign n1293 = ~n4005;
  assign n2749 = n3903 ^ n3828;
  assign n3846 = n3903 & n2773;
  assign n3904 = n3903 & n3910;
  assign n3895 = n3924 & n3925;
  assign n3919 = n3943 & n3944;
  assign n3957 = n3964 & n3965;
  assign n3906 = ~n3966;
  assign n3945 = n3967 & n3968;
  assign n78275 = n3974 ^ n1183;
  assign n3978 = n1183 & n3984;
  assign n3976 = ~n1183;
  assign n3929 = n3996 ^ n1228;
  assign n3997 = n1293 & n4002;
  assign n2746 = ~n4003;
  assign n4000 = ~n4008;
  assign n2748 = n2749 ^ n2728;
  assign n3883 = ~n3846;
  assign n3831 = ~n3904;
  assign n3926 = ~n3919;
  assign n3928 = n3945 ^ n3946;
  assign n3927 = ~n3957;
  assign n3947 = ~n3945;
  assign n3934 = n3976 & n3974;
  assign n3969 = n3929 & n3946;
  assign n3949 = n3976 & n2608;
  assign n3972 = n3976 & n3977;
  assign n2657 = ~n3978;
  assign n3970 = ~n3929;
  assign n2719 = ~n3997;
  assign n3979 = n4000 & n4001;
  assign n3825 = n2748 & n2728;
  assign n3854 = n2748 & n3861;
  assign n78348 = ~n2748;
  assign n3875 = n3883 & n3779;
  assign n3921 = n3926 & n3927;
  assign n3857 = n3928 ^ n3929;
  assign n3940 = n3927 & n3906;
  assign n3885 = n3949 ^ n1088;
  assign n3948 = ~n3969;
  assign n3958 = n3970 & n3971;
  assign n2689 = ~n3972;
  assign n3950 = n3979 ^ n1074;
  assign n2743 = n2746 & n2719;
  assign n3980 = ~n3979;
  assign n3806 = n3825 ^ n78252;
  assign n3829 = n3825 & n3845;
  assign n3827 = ~n3825;
  assign n3793 = ~n3854;
  assign n3862 = ~n3875;
  assign n3907 = n3857 & n3911;
  assign n3905 = ~n3921;
  assign n3908 = ~n3857;
  assign n3920 = ~n3940;
  assign n3941 = n3947 & n3948;
  assign n2686 = n2689 & n2657;
  assign n1125 = n3950 ^ n3951;
  assign n3931 = ~n3958;
  assign n3973 = n3980 & n3981;
  assign n3739 = n3806 & n3807;
  assign n3810 = n3793 & n3826;
  assign n3811 = n3827 & n3828;
  assign n3791 = ~n3829;
  assign n3876 = n3905 & n3906;
  assign n3878 = ~n3907;
  assign n3897 = n3908 & n383;
  assign n3896 = n3919 ^ n3920;
  assign n78274 = n3934 ^ n1125;
  assign n3930 = ~n3941;
  assign n3936 = n1125 & n2600;
  assign n2543 = ~n1125;
  assign n3952 = ~n3973;
  assign n3769 = n3739 & n3710;
  assign n3767 = ~n3739;
  assign n3790 = ~n3810;
  assign n3792 = ~n3811;
  assign n3856 = n383 ^ n3876;
  assign n3863 = n3895 ^ n3896;
  assign n3877 = ~n3876;
  assign n3859 = ~n3897;
  assign n3812 = n3896 & n3895;
  assign n3912 = n3930 & n3931;
  assign n3873 = n2543 & n3934;
  assign n3914 = n2543 & n2403;
  assign n3932 = n2543 & n3935;
  assign n2603 = ~n3936;
  assign n3937 = n3952 & n3953;
  assign n3750 = n3767 & n3768;
  assign n3703 = ~n3769;
  assign n3780 = n3790 & n3791;
  assign n3781 = n3792 & n3793;
  assign n3813 = n3856 ^ n3857;
  assign n3855 = n3862 & n3863;
  assign n3847 = n3863 ^ n3779;
  assign n3870 = n3877 & n3878;
  assign n3815 = ~n3812;
  assign n3909 = n3912 & n3913;
  assign n3900 = n3914 ^ n1029;
  assign n3898 = ~n3912;
  assign n3902 = ~n3873;
  assign n2632 = ~n3932;
  assign n3916 = n3937 ^ n974;
  assign n3938 = ~n3937;
  assign n3730 = ~n3750;
  assign n3753 = ~n3780;
  assign n3751 = ~n3781;
  assign n3783 = n3812 ^ n3813;
  assign n78347 = n3846 ^ n3847;
  assign n3814 = ~n3813;
  assign n3830 = ~n3855;
  assign n3858 = ~n3870;
  assign n3871 = n3898 ^ n3885;
  assign n3888 = n3900 & n3901;
  assign n3899 = n3898 & n3872;
  assign n3884 = ~n3909;
  assign n3886 = ~n3900;
  assign n1076 = n3915 ^ n3916;
  assign n3933 = n3938 & n3939;
  assign n3740 = n3751 & n3752;
  assign n3741 = n3753 & n3754;
  assign n3770 = ~n3783;
  assign n3778 = n78347 & n2695;
  assign n3743 = n3814 & n3815;
  assign n2730 = ~n78347;
  assign n3782 = n3830 & n3831;
  assign n3816 = n3858 & n3859;
  assign n3817 = n3871 ^ n3872;
  assign n3879 = n3884 & n3885;
  assign n3880 = n3886 & n3887;
  assign n3799 = ~n3888;
  assign n3865 = ~n3899;
  assign n3824 = n1076 & n3902;
  assign n3889 = n1076 & n2572;
  assign n3874 = ~n1076;
  assign n3917 = ~n3933;
  assign n3718 = ~n3740;
  assign n3719 = ~n3741;
  assign n3731 = n3778 ^ n3779;
  assign n3742 = n3782 ^ n3783;
  assign n3795 = n3782 & n3693;
  assign n3746 = ~n3743;
  assign n3794 = ~n3782;
  assign n3785 = n3816 ^ n3817;
  assign n3808 = ~n3816;
  assign n3850 = n3817 & n382;
  assign n3848 = ~n3817;
  assign n78273 = n3873 ^ n3874;
  assign n3864 = ~n3879;
  assign n3834 = ~n3880;
  assign n3866 = n3874 & n2426;
  assign n2534 = ~n3889;
  assign n3881 = n3874 & n3890;
  assign n3891 = n3917 & n3918;
  assign n3691 = n3718 & n3719;
  assign n3717 = n3730 & n3731;
  assign n3709 = n3739 ^ n3731;
  assign n2565 = n3742 ^ n3693;
  assign n3744 = n382 ^ n3785;
  assign n3784 = n3794 & n2598;
  assign n3771 = ~n3795;
  assign n3832 = n3848 & n3849;
  assign n3773 = ~n3850;
  assign n3818 = n3864 & n3865;
  assign n3860 = n3834 & n3799;
  assign n3851 = n3866 ^ n974;
  assign n2574 = ~n3881;
  assign n3867 = n3891 ^ n3892;
  assign n3893 = ~n3891;
  assign n3112 = n71 ^ n3691;
  assign n3690 = n3709 ^ n3710;
  assign n3694 = ~n3691;
  assign n3702 = ~n3717;
  assign n3692 = n2565 & n2536;
  assign n3616 = n2565 & n78347;
  assign n2682 = ~n2565;
  assign n3720 = n3743 ^ n3744;
  assign n3755 = n3770 & n3771;
  assign n3745 = ~n3744;
  assign n3733 = ~n3784;
  assign n3809 = ~n3832;
  assign n3835 = n3851 & n3852;
  assign n3833 = ~n3818;
  assign n3819 = ~n3860;
  assign n3836 = ~n3851;
  assign n1010 = n957 ^ n3867;
  assign n3882 = n3893 & n3894;
  assign n3124 = ~n3112;
  assign n3686 = n3690 & n70;
  assign n3644 = n3692 ^ n3693;
  assign n3606 = n3694 & n71;
  assign n78346 = n2682 ^ n78347;
  assign n3684 = ~n3690;
  assign n3671 = n3702 & n3703;
  assign n3622 = ~n3616;
  assign n3711 = n3720 & n2531;
  assign n3712 = ~n3720;
  assign n3677 = n3745 & n3746;
  assign n3732 = ~n3755;
  assign n3796 = n3808 & n3809;
  assign n3797 = n3818 ^ n3819;
  assign n78272 = n3824 ^ n1010;
  assign n3820 = n3833 & n3834;
  assign n3725 = ~n3835;
  assign n3821 = n3836 & n3837;
  assign n3776 = n1010 & n3824;
  assign n3839 = n1010 & n3853;
  assign n3838 = ~n1010;
  assign n3868 = ~n3882;
  assign n3643 = n3671 ^ n3672;
  assign n3670 = n3684 & n3685;
  assign n3619 = ~n3686;
  assign n3675 = n3671 & n3672;
  assign n3673 = ~n3671;
  assign n3660 = ~n3711;
  assign n3704 = n3712 & n3713;
  assign n3658 = n3732 & n3733;
  assign n3680 = ~n3677;
  assign n3772 = ~n3796;
  assign n3788 = n3797 & n381;
  assign n3786 = ~n3797;
  assign n3798 = ~n3820;
  assign n3759 = ~n3821;
  assign n3801 = ~n3776;
  assign n3800 = n3838 & n2388;
  assign n2458 = ~n3839;
  assign n3822 = n3838 & n3840;
  assign n3841 = n3868 & n3869;
  assign n3617 = n3643 ^ n3644;
  assign n3655 = ~n3670;
  assign n3663 = n3673 & n3674;
  assign n3656 = ~n3675;
  assign n3688 = ~n3704;
  assign n3687 = ~n3658;
  assign n3707 = n3772 & n3773;
  assign n3774 = n3786 & n3787;
  assign n3706 = ~n3788;
  assign n3757 = n3798 & n3799;
  assign n3756 = n3759 & n3725;
  assign n3696 = n3800 ^ n957;
  assign n2501 = ~n3822;
  assign n977 = n3841 ^ n3842;
  assign n3843 = ~n3841;
  assign n3605 = n3617 & n69;
  assign n3603 = ~n3617;
  assign n3645 = n3606 & n3655;
  assign n3646 = n3655 & n3619;
  assign n3647 = n3644 & n3656;
  assign n3621 = ~n3663;
  assign n3676 = n3687 & n3688;
  assign n3657 = n3688 & n3660;
  assign n3734 = ~n3707;
  assign n3650 = n3756 ^ n3757;
  assign n3735 = ~n3774;
  assign n3760 = n3696 & n3775;
  assign n3758 = ~n3757;
  assign n3761 = ~n3696;
  assign n2498 = n2501 & n2458;
  assign n3802 = n977 & n2417;
  assign n3777 = ~n977;
  assign n3823 = n3843 & n3844;
  assign n3594 = n3603 & n3604;
  assign n3550 = ~n3605;
  assign n3618 = ~n3645;
  assign n3607 = ~n3646;
  assign n3620 = ~n3647;
  assign n2503 = n3657 ^ n3658;
  assign n3659 = ~n3676;
  assign n3721 = n3734 & n3735;
  assign n3722 = n3650 & n3736;
  assign n3737 = n3735 & n3706;
  assign n3723 = ~n3650;
  assign n3747 = n3758 & n3759;
  assign n3698 = ~n3760;
  assign n3748 = n3761 & n3665;
  assign n78271 = n3776 ^ n3777;
  assign n3716 = n3777 & n3801;
  assign n3762 = n3777 & n2262;
  assign n2378 = ~n3802;
  assign n3789 = n3777 & n3803;
  assign n3804 = ~n3823;
  assign n3582 = ~n3594;
  assign n3580 = n3606 ^ n3607;
  assign n78345 = n3616 ^ n2503;
  assign n3540 = n3618 & n3619;
  assign n3589 = n3620 & n3621;
  assign n3595 = n2503 & n2472;
  assign n2616 = ~n2503;
  assign n3623 = n3659 & n3660;
  assign n3705 = ~n3721;
  assign n3683 = ~n3722;
  assign n3714 = n3723 & n380;
  assign n3708 = ~n3737;
  assign n3724 = ~n3747;
  assign n3668 = ~n3748;
  assign n3599 = n3762 ^ n927;
  assign n2419 = ~n3789;
  assign n3763 = n3804 & n3805;
  assign n3049 = n3580 ^ n3112;
  assign n3059 = n3580 ^ n3124;
  assign n3571 = n3582 & n3550;
  assign n3506 = n3580 & n3112;
  assign n3562 = n3589 ^ n3584;
  assign n3583 = n3595 ^ n2531;
  assign n3581 = ~n3540;
  assign n3552 = ~n3589;
  assign n3560 = n2616 & n3622;
  assign n3626 = ~n3623;
  assign n3681 = n3705 & n3706;
  assign n3678 = n3707 ^ n3708;
  assign n3652 = ~n3714;
  assign n3695 = n3724 & n3725;
  assign n877 = n3763 ^ n3764;
  assign n3765 = ~n3763;
  assign n3541 = ~n3571;
  assign n3570 = n3581 & n3582;
  assign n3519 = ~n3506;
  assign n3573 = n3583 & n3584;
  assign n3561 = ~n3583;
  assign n3572 = ~n3560;
  assign n3661 = n3677 ^ n3678;
  assign n3649 = n380 ^ n3681;
  assign n3682 = ~n3681;
  assign n3679 = ~n3678;
  assign n3664 = n3695 ^ n3696;
  assign n3697 = ~n3695;
  assign n78270 = n3716 ^ n877;
  assign n3727 = n877 & n3738;
  assign n3726 = ~n877;
  assign n3749 = n3765 & n3766;
  assign n3507 = n3540 ^ n3541;
  assign n3508 = n3561 ^ n3562;
  assign n3549 = ~n3570;
  assign n3551 = ~n3573;
  assign n3563 = n3561 & n3574;
  assign n3610 = n3649 ^ n3650;
  assign n3648 = n3661 & n3662;
  assign n3624 = ~n3661;
  assign n3613 = n3664 ^ n3665;
  assign n3609 = n3679 & n3680;
  assign n3666 = n3682 & n3683;
  assign n3689 = n3697 & n3698;
  assign n3630 = n3726 & n3716;
  assign n3699 = n3726 & n2182;
  assign n2290 = ~n3727;
  assign n3715 = n3726 & n2332;
  assign n3728 = ~n3749;
  assign n1691 = n3506 ^ n3507;
  assign n3458 = n3507 & n3519;
  assign n3532 = n3508 & n68;
  assign n3542 = n3549 & n3550;
  assign n3530 = ~n3508;
  assign n3544 = n3551 & n3552;
  assign n3524 = ~n3563;
  assign n3534 = n3609 ^ n3610;
  assign n3590 = n3623 ^ n3624;
  assign n3611 = ~n3610;
  assign n3625 = ~n3648;
  assign n3632 = n3624 & n2433;
  assign n3635 = n3613 & n379;
  assign n3633 = ~n3613;
  assign n3651 = ~n3666;
  assign n3667 = ~n3689;
  assign n3527 = n3699 ^ n817;
  assign n2303 = ~n3715;
  assign n3700 = n3728 & n3729;
  assign n3025 = ~n1691;
  assign n3461 = ~n3458;
  assign n3520 = n3530 & n3531;
  assign n3476 = ~n3532;
  assign n3500 = ~n3542;
  assign n3523 = ~n3544;
  assign n2392 = n2433 ^ n3590;
  assign n3554 = n3611 & n3609;
  assign n3608 = n3625 & n3626;
  assign n3592 = ~n3632;
  assign n3627 = n3633 & n3634;
  assign n3576 = ~n3635;
  assign n3612 = n3651 & n3652;
  assign n3636 = n3667 & n3668;
  assign n3669 = n3700 ^ n3701;
  assign n3485 = n3500 ^ n3508;
  assign n3499 = ~n3520;
  assign n3447 = n3523 & n3524;
  assign n78344 = n3560 ^ n2392;
  assign n3498 = n2392 & n3572;
  assign n3543 = n2392 & n2365;
  assign n2569 = ~n2392;
  assign n3591 = ~n3608;
  assign n3585 = n3612 ^ n3613;
  assign n3596 = ~n3627;
  assign n3597 = ~n3612;
  assign n3598 = n3636 ^ n3637;
  assign n3640 = n3636 & n3637;
  assign n3638 = ~n3636;
  assign n3631 = n3669 ^ n726;
  assign n3459 = n68 ^ n3485;
  assign n3494 = n3499 & n3500;
  assign n3495 = ~n3447;
  assign n3521 = n3543 ^ n2433;
  assign n3555 = n379 ^ n3585;
  assign n3564 = n3591 & n3592;
  assign n3593 = n3596 & n3597;
  assign n3586 = n3598 ^ n3599;
  assign n78269 = n3630 ^ n3631;
  assign n3628 = n3638 & n3639;
  assign n3614 = ~n3640;
  assign n3615 = n3631 & n3653;
  assign n3642 = n3631 & n3654;
  assign n832 = ~n3631;
  assign n1625 = n3458 ^ n3459;
  assign n3460 = ~n3459;
  assign n3475 = ~n3494;
  assign n3511 = n3521 & n3522;
  assign n3509 = ~n3521;
  assign n3536 = n3554 ^ n3555;
  assign n3533 = n3564 ^ n3565;
  assign n3491 = n3555 & n3554;
  assign n3567 = n3564 & n3565;
  assign n3566 = ~n3564;
  assign n3579 = n3586 & n378;
  assign n3575 = ~n3593;
  assign n3577 = ~n3586;
  assign n3600 = n3614 & n3599;
  assign n3456 = n3615 ^ n726;
  assign n3588 = ~n3628;
  assign n3629 = n832 & n3641;
  assign n3601 = ~n3642;
  assign n2964 = ~n1625;
  assign n3389 = n3460 & n3461;
  assign n3428 = n3475 & n3476;
  assign n3501 = n3509 & n3510;
  assign n3487 = ~n3511;
  assign n2340 = n3533 ^ n3534;
  assign n3526 = n3536 & n3537;
  assign n3525 = ~n3536;
  assign n3553 = n3566 & n2383;
  assign n3545 = ~n3567;
  assign n3516 = n3575 & n3576;
  assign n3568 = n3577 & n3578;
  assign n3518 = ~n3579;
  assign n3587 = ~n3600;
  assign n3602 = ~n3629;
  assign n3414 = ~n3428;
  assign n3486 = n3487 & n3495;
  assign n78343 = n3498 ^ n2340;
  assign n3471 = ~n3501;
  assign n2478 = ~n2340;
  assign n3514 = n3525 & n2281;
  assign n3489 = ~n3526;
  assign n3535 = n3545 & n3534;
  assign n3513 = ~n3553;
  assign n3547 = ~n3516;
  assign n3546 = ~n3568;
  assign n3556 = n3587 & n3588;
  assign n2266 = n3601 & n3602;
  assign n3470 = ~n3486;
  assign n3477 = n3471 & n3487;
  assign n3478 = n2478 & n2295;
  assign n3442 = n2478 & n3498;
  assign n3465 = ~n3514;
  assign n3512 = ~n3535;
  assign n3538 = n3546 & n3547;
  assign n3515 = n3546 & n3518;
  assign n3528 = n3556 ^ n3557;
  assign n3559 = n3556 & n3569;
  assign n3558 = ~n3556;
  assign n2248 = ~n2266;
  assign n3407 = n3470 & n3471;
  assign n3448 = ~n3477;
  assign n3462 = n3478 ^ n2383;
  assign n3490 = n3489 & n3465;
  assign n3466 = n3512 & n3513;
  assign n3492 = n3515 ^ n3516;
  assign n3482 = n3527 ^ n3528;
  assign n3517 = ~n3538;
  assign n3548 = n3558 & n3557;
  assign n3539 = ~n3559;
  assign n3429 = n3447 ^ n3448;
  assign n3443 = ~n3407;
  assign n3451 = n3462 & n3463;
  assign n3449 = ~n3462;
  assign n3467 = ~n3490;
  assign n3472 = n3491 ^ n3492;
  assign n3436 = n3492 & n3491;
  assign n3488 = ~n3466;
  assign n3496 = n3482 & n3502;
  assign n3503 = n3517 & n3518;
  assign n3497 = ~n3482;
  assign n3529 = n3539 & n3527;
  assign n3505 = ~n3548;
  assign n3412 = n3428 ^ n3429;
  assign n3432 = n3429 & n67;
  assign n3430 = ~n3429;
  assign n3446 = n3449 & n3450;
  assign n3434 = ~n3451;
  assign n2237 = n3466 ^ n3467;
  assign n3468 = n3472 & n3473;
  assign n3469 = ~n3472;
  assign n3479 = n3488 & n3489;
  assign n3439 = ~n3436;
  assign n3480 = ~n3496;
  assign n3493 = n3497 & n377;
  assign n3481 = ~n3503;
  assign n3504 = ~n3529;
  assign n3390 = n67 ^ n3412;
  assign n3426 = n3430 & n3431;
  assign n3392 = ~n3432;
  assign n78342 = n3442 ^ n2237;
  assign n3433 = n3434 & n3443;
  assign n3420 = ~n3446;
  assign n2384 = ~n2237;
  assign n3444 = ~n3468;
  assign n3452 = n3469 & n2212;
  assign n3464 = ~n3479;
  assign n3474 = n3480 & n3481;
  assign n3453 = n3481 ^ n3482;
  assign n3455 = ~n3493;
  assign n3483 = n3504 & n3505;
  assign n2920 = n3389 ^ n3390;
  assign n3331 = n3390 & n3389;
  assign n3413 = ~n3426;
  assign n3419 = ~n3433;
  assign n3427 = n3434 & n3420;
  assign n3421 = n2384 & n2108;
  assign n3399 = n2384 & n3442;
  assign n3423 = ~n3452;
  assign n3437 = n377 ^ n3453;
  assign n3425 = n3464 & n3465;
  assign n3454 = ~n3474;
  assign n3457 = n3483 ^ n3484;
  assign n2933 = ~n2920;
  assign n3406 = n3413 & n3414;
  assign n3359 = n3419 & n3420;
  assign n3409 = n3421 ^ n2281;
  assign n3408 = ~n3427;
  assign n3405 = ~n3399;
  assign n3404 = n3436 ^ n3437;
  assign n3424 = n3423 & n3444;
  assign n3438 = ~n3437;
  assign n3445 = ~n3425;
  assign n3440 = n3454 & n3455;
  assign n3441 = n3456 ^ n3457;
  assign n3391 = ~n3406;
  assign n3393 = n3407 ^ n3408;
  assign n3402 = n3409 & n3410;
  assign n3386 = ~n3359;
  assign n3400 = ~n3409;
  assign n3415 = n3404 & n2112;
  assign n2169 = n3424 ^ n3425;
  assign n3416 = ~n3404;
  assign n3395 = n3438 & n3439;
  assign n3418 = n3440 ^ n3441;
  assign n3435 = n3444 & n3445;
  assign n3348 = n3391 & n3392;
  assign n3385 = n3393 & n66;
  assign n78341 = n3399 ^ n2169;
  assign n3383 = ~n3393;
  assign n3394 = n3400 & n3401;
  assign n3382 = ~n3402;
  assign n3387 = n2169 & n2151;
  assign n3378 = ~n3415;
  assign n3411 = n3416 & n3417;
  assign n3396 = n376 ^ n3418;
  assign n2345 = ~n2169;
  assign n3422 = ~n3435;
  assign n3365 = ~n3348;
  assign n3379 = n3383 & n3384;
  assign n3350 = ~n3385;
  assign n3380 = n3382 & n3386;
  assign n3372 = n3387 ^ n2212;
  assign n3367 = ~n3394;
  assign n3339 = n3395 ^ n3396;
  assign n3358 = n2345 & n3405;
  assign n3398 = ~n3411;
  assign n3403 = n3422 & n3423;
  assign n3368 = n3372 & n3353;
  assign n3364 = ~n3379;
  assign n3366 = ~n3380;
  assign n3375 = n3382 & n3367;
  assign n3376 = n3339 & n2042;
  assign n3333 = ~n3372;
  assign n3373 = ~n3339;
  assign n3381 = n3403 ^ n3404;
  assign n3397 = ~n3403;
  assign n3362 = n3364 & n3365;
  assign n3347 = n3364 & n3350;
  assign n3352 = n3366 & n3367;
  assign n3354 = ~n3368;
  assign n3363 = n3333 & n3369;
  assign n3370 = n3373 & n3374;
  assign n3360 = ~n3375;
  assign n3345 = ~n3376;
  assign n2074 = n3381 ^ n2112;
  assign n3388 = n3397 & n3398;
  assign n3332 = n3347 ^ n3348;
  assign n3334 = n3352 ^ n3353;
  assign n3313 = n3359 ^ n3360;
  assign n3349 = ~n3362;
  assign n3355 = ~n3352;
  assign n3337 = ~n3363;
  assign n3351 = n2074 & n2045;
  assign n3361 = ~n3370;
  assign n2232 = ~n2074;
  assign n3377 = ~n3388;
  assign n2892 = n3331 ^ n3332;
  assign n3324 = n3333 ^ n3334;
  assign n3294 = n3332 & n3331;
  assign n3343 = n3313 & n65;
  assign n3335 = n3349 & n3350;
  assign n3299 = n3351 ^ n2112;
  assign n3346 = n3354 & n3355;
  assign n3341 = ~n3313;
  assign n78356 = n3358 ^ n2232;
  assign n3311 = n2232 & n3358;
  assign n3371 = n3377 & n3378;
  assign n3316 = n3324 & n64;
  assign n2883 = ~n2892;
  assign n3314 = ~n3324;
  assign n3297 = ~n3294;
  assign n3312 = n65 ^ n3335;
  assign n3338 = n3341 & n3342;
  assign n3303 = ~n3343;
  assign n3326 = ~n3335;
  assign n3305 = ~n3299;
  assign n3336 = ~n3346;
  assign n3357 = ~n3371;
  assign n3295 = n3312 ^ n3313;
  assign n3309 = n3314 & n3315;
  assign n3262 = ~n3316;
  assign n3317 = n3336 & n3337;
  assign n3325 = ~n3338;
  assign n3340 = n3357 ^ n2042;
  assign n3356 = n3357 & n3361;
  assign n1444 = n3294 ^ n3295;
  assign n3296 = ~n3295;
  assign n3281 = ~n3309;
  assign n3298 = n3317 ^ n3318;
  assign n3319 = n3325 & n3326;
  assign n3322 = n3317 & n3318;
  assign n3320 = ~n3317;
  assign n2174 = n3339 ^ n3340;
  assign n3344 = ~n3356;
  assign n2851 = ~n1444;
  assign n3252 = n3296 & n3297;
  assign n3292 = n3281 & n3262;
  assign n3241 = n3298 ^ n3299;
  assign n78355 = n3311 ^ n2174;
  assign n3302 = ~n3319;
  assign n3310 = n3320 & n3321;
  assign n3304 = ~n3322;
  assign n3291 = n2174 & n3311;
  assign n2005 = ~n2174;
  assign n3327 = n3344 & n3345;
  assign n3273 = n3241 & n3280;
  assign n3255 = ~n3252;
  assign n3269 = ~n3292;
  assign n3274 = ~n3241;
  assign n3268 = n3302 & n3303;
  assign n3300 = n3304 & n3305;
  assign n3284 = ~n3310;
  assign n3301 = n2005 & n1979;
  assign n3293 = ~n3291;
  assign n3306 = n3327 ^ n3328;
  assign n3329 = ~n3327;
  assign n3253 = n3268 ^ n3269;
  assign n3242 = ~n3273;
  assign n3270 = n3274 & n79;
  assign n3282 = ~n3268;
  assign n3283 = ~n3300;
  assign n3285 = n3301 ^ n2042;
  assign n1947 = n1981 ^ n3306;
  assign n3323 = n3329 & n3330;
  assign n2822 = n3252 ^ n3253;
  assign n3254 = ~n3253;
  assign n3228 = ~n3270;
  assign n3275 = n3281 & n3282;
  assign n3236 = n3283 & n3284;
  assign n3276 = n3285 & n3286;
  assign n78354 = n3291 ^ n1947;
  assign n3239 = n1947 & n3293;
  assign n3271 = n1947 & n1927;
  assign n3277 = ~n3285;
  assign n2080 = ~n1947;
  assign n3307 = ~n3323;
  assign n2811 = ~n2822;
  assign n3200 = n3254 & n3255;
  assign n3257 = n3271 ^ n1981;
  assign n3261 = ~n3275;
  assign n3263 = ~n3236;
  assign n3260 = ~n3276;
  assign n3272 = n3277 & n3278;
  assign n3247 = ~n3239;
  assign n3287 = n3307 & n3308;
  assign n3212 = ~n3200;
  assign n3256 = n3257 & n3258;
  assign n3240 = n3261 & n3262;
  assign n3196 = ~n3257;
  assign n3259 = n3263 & n3260;
  assign n3246 = ~n3272;
  assign n3264 = n3287 ^ n3288;
  assign n3289 = ~n3287;
  assign n3225 = n3240 ^ n3241;
  assign n3226 = ~n3256;
  assign n3244 = n3196 & n3223;
  assign n3243 = ~n3240;
  assign n3245 = ~n3259;
  assign n3235 = n3246 & n3260;
  assign n1889 = n3264 ^ n3265;
  assign n3279 = n3289 & n3290;
  assign n3201 = n79 ^ n3225;
  assign n3186 = n3235 ^ n3236;
  assign n78353 = n3239 ^ n1889;
  assign n3234 = n3242 & n3243;
  assign n3204 = ~n3244;
  assign n3237 = n3245 & n3246;
  assign n3233 = n1889 & n1867;
  assign n1958 = ~n1889;
  assign n3266 = ~n3279;
  assign n1331 = n3200 ^ n3201;
  assign n3166 = n3201 & n3212;
  assign n3220 = n3186 & n3229;
  assign n3188 = n3233 ^ n1912;
  assign n3221 = ~n3186;
  assign n3227 = ~n3234;
  assign n3222 = ~n3237;
  assign n3224 = n1958 & n3247;
  assign n3249 = n3266 & n3267;
  assign n2769 = ~n1331;
  assign n3169 = ~n3166;
  assign n3213 = n3188 & n3218;
  assign n3205 = ~n3220;
  assign n3215 = n3221 & n78;
  assign n3197 = n3222 ^ n3223;
  assign n3219 = n3222 & n3226;
  assign n3202 = n3227 & n3228;
  assign n3214 = ~n3188;
  assign n3230 = ~n3224;
  assign n1832 = n3248 ^ n3249;
  assign n3250 = ~n3249;
  assign n3150 = n3196 ^ n3197;
  assign n3185 = n78 ^ n3202;
  assign n3190 = ~n3213;
  assign n3207 = n3214 & n3171;
  assign n3192 = ~n3215;
  assign n3203 = ~n3219;
  assign n3206 = ~n3202;
  assign n78352 = n3224 ^ n1832;
  assign n3175 = n1832 & n3230;
  assign n3216 = n1832 & n1825;
  assign n1933 = ~n1832;
  assign n3238 = n3250 & n3251;
  assign n3167 = n3185 ^ n3186;
  assign n3183 = n3150 & n77;
  assign n3181 = ~n3150;
  assign n3187 = n3203 & n3204;
  assign n3198 = n3205 & n3206;
  assign n3174 = ~n3207;
  assign n3131 = n3216 ^ n3217;
  assign n3176 = ~n3175;
  assign n3231 = ~n3238;
  assign n2726 = n3166 ^ n3167;
  assign n3168 = ~n3167;
  assign n3180 = n3181 & n3182;
  assign n3144 = ~n3183;
  assign n3170 = n3187 ^ n3188;
  assign n3189 = ~n3187;
  assign n3191 = ~n3198;
  assign n3208 = n3231 & n3232;
  assign n2716 = ~n2726;
  assign n3127 = n3168 & n3169;
  assign n3120 = n3170 ^ n3171;
  assign n3163 = ~n3180;
  assign n3184 = n3189 & n3190;
  assign n3172 = n3191 & n3192;
  assign n3193 = n3208 ^ n3209;
  assign n3210 = ~n3208;
  assign n3148 = n3120 & n76;
  assign n3130 = ~n3127;
  assign n3146 = ~n3120;
  assign n3149 = n77 ^ n3172;
  assign n3173 = ~n3184;
  assign n3164 = ~n3172;
  assign n1804 = n3193 ^ n1826;
  assign n3199 = n3210 & n3211;
  assign n3142 = n3146 & n3147;
  assign n3103 = ~n3148;
  assign n3128 = n3149 ^ n3150;
  assign n3159 = n3163 & n3164;
  assign n3151 = n3173 & n3174;
  assign n78351 = n3175 ^ n1804;
  assign n3161 = n1804 & n1786;
  assign n1894 = ~n1804;
  assign n3194 = ~n3199;
  assign n1237 = n3127 ^ n3128;
  assign n3125 = ~n3142;
  assign n3129 = ~n3128;
  assign n3132 = n3151 ^ n3152;
  assign n3143 = ~n3159;
  assign n3154 = n3151 & n3160;
  assign n3073 = n3161 ^ n3162;
  assign n3153 = ~n3151;
  assign n3134 = n1894 & n3176;
  assign n3177 = n3194 & n3195;
  assign n2665 = ~n1237;
  assign n3070 = n3129 & n3130;
  assign n3080 = n3131 ^ n3132;
  assign n3139 = n3143 & n3144;
  assign n3145 = n3153 & n3152;
  assign n3140 = ~n3154;
  assign n3141 = ~n3134;
  assign n3156 = n3177 ^ n1785;
  assign n3178 = ~n3177;
  assign n3108 = n3080 & n3117;
  assign n3109 = ~n3080;
  assign n3119 = ~n3139;
  assign n3133 = n3140 & n3131;
  assign n3122 = ~n3145;
  assign n1858 = n3155 ^ n3156;
  assign n3165 = n3178 & n3179;
  assign n3082 = ~n3108;
  assign n3104 = n3109 & n75;
  assign n3092 = n3119 ^ n3120;
  assign n3118 = n3125 & n3119;
  assign n3121 = ~n3133;
  assign n78350 = n3134 ^ n1858;
  assign n3116 = n1858 & n3141;
  assign n3123 = n1858 & n1743;
  assign n1766 = ~n1858;
  assign n3157 = ~n3165;
  assign n3071 = n76 ^ n3092;
  assign n3062 = ~n3104;
  assign n3102 = ~n3118;
  assign n3093 = n3121 & n3122;
  assign n3105 = n3123 ^ n1785;
  assign n3111 = ~n3116;
  assign n3136 = n3157 & n3158;
  assign n1186 = n3070 ^ n3071;
  assign n3035 = n3071 & n3070;
  assign n3072 = n3093 ^ n3094;
  assign n3079 = n3102 & n3103;
  assign n3097 = n3093 & n3094;
  assign n3098 = n3105 & n3106;
  assign n3095 = ~n3093;
  assign n3099 = ~n3105;
  assign n1731 = n3135 ^ n3136;
  assign n3137 = ~n3136;
  assign n2579 = ~n1186;
  assign n3038 = ~n3035;
  assign n3032 = n3072 ^ n3073;
  assign n3060 = n3079 ^ n3080;
  assign n3081 = ~n3079;
  assign n3087 = n3095 & n3096;
  assign n3083 = ~n3097;
  assign n3042 = ~n3098;
  assign n3088 = n3099 & n3100;
  assign n1775 = n3112 ^ n1731;
  assign n78349 = n3116 ^ n1731;
  assign n3113 = n1731 & n3124;
  assign n3101 = n1731 & n1722;
  assign n3110 = ~n1731;
  assign n3126 = n3137 & n3138;
  assign n3036 = n75 ^ n3060;
  assign n3057 = n3032 & n74;
  assign n3055 = ~n3032;
  assign n3074 = n3081 & n3082;
  assign n3075 = n3083 & n3073;
  assign n3064 = ~n3087;
  assign n3018 = ~n3088;
  assign n3084 = n3101 ^ n1756;
  assign n3054 = n3110 & n3111;
  assign n1777 = ~n3113;
  assign n3107 = n3110 & n3112;
  assign n3114 = ~n3126;
  assign n1093 = n3035 ^ n3036;
  assign n3037 = ~n3036;
  assign n3045 = n3055 & n3056;
  assign n3011 = ~n3057;
  assign n3061 = ~n3074;
  assign n3063 = ~n3075;
  assign n3039 = n3042 & n3018;
  assign n3076 = n3084 & n3085;
  assign n3077 = ~n3084;
  assign n1758 = ~n3107;
  assign n3089 = n3114 & n3115;
  assign n2497 = ~n1093;
  assign n2985 = n3037 & n3038;
  assign n3030 = ~n3045;
  assign n3058 = n3061 & n3062;
  assign n3040 = n3063 & n3064;
  assign n2998 = ~n3076;
  assign n3065 = n3077 & n3078;
  assign n3067 = n3089 ^ n3023;
  assign n3090 = ~n3089;
  assign n2994 = ~n2985;
  assign n2970 = n3039 ^ n3040;
  assign n3031 = ~n3058;
  assign n3041 = ~n3040;
  assign n2978 = ~n3065;
  assign n1698 = n3066 ^ n3067;
  assign n3086 = n3090 & n3091;
  assign n3015 = n2970 & n3021;
  assign n3020 = n3030 & n3031;
  assign n3009 = n3031 ^ n3032;
  assign n3016 = ~n2970;
  assign n3033 = n3041 & n3042;
  assign n78364 = n3054 ^ n1698;
  assign n3046 = n2998 & n2978;
  assign n3048 = n1698 & n3059;
  assign n3029 = n1698 & n3054;
  assign n3047 = ~n1698;
  assign n3068 = ~n3086;
  assign n2986 = n74 ^ n3009;
  assign n2989 = ~n3015;
  assign n3012 = n3016 & n73;
  assign n3010 = ~n3020;
  assign n3017 = ~n3033;
  assign n2996 = ~n3046;
  assign n3022 = n3047 & n1591;
  assign n1714 = ~n3048;
  assign n3043 = n3047 & n3049;
  assign n3034 = ~n3029;
  assign n3051 = n3068 & n3069;
  assign n1032 = n2985 ^ n2986;
  assign n2944 = n2986 & n2994;
  assign n2987 = n3010 & n3011;
  assign n2972 = ~n3012;
  assign n2995 = n3017 & n3018;
  assign n2935 = n3022 ^ n3023;
  assign n1735 = ~n3043;
  assign n1640 = n3050 ^ n3051;
  assign n3052 = ~n3051;
  assign n2456 = ~n1032;
  assign n2947 = ~n2944;
  assign n2969 = n73 ^ n2987;
  assign n2949 = n2995 ^ n2996;
  assign n2988 = ~n2987;
  assign n2997 = ~n2995;
  assign n3004 = n2935 & n3013;
  assign n3003 = ~n2935;
  assign n1732 = n1735 & n1714;
  assign n78363 = n3029 ^ n1640;
  assign n2960 = n1640 & n3034;
  assign n3014 = n1640 & n1528;
  assign n3026 = n1640 & n1691;
  assign n3024 = ~n1640;
  assign n3044 = n3052 & n3053;
  assign n2945 = n2969 ^ n2970;
  assign n2976 = n2949 & n72;
  assign n2979 = n2988 & n2989;
  assign n2974 = ~n2949;
  assign n2990 = n2997 & n2998;
  assign n2999 = n3003 & n2955;
  assign n2937 = ~n3004;
  assign n3000 = n3014 ^ n1659;
  assign n2962 = ~n2960;
  assign n3019 = n3024 & n3025;
  assign n1693 = ~n3026;
  assign n3027 = ~n3044;
  assign n2349 = n2944 ^ n2945;
  assign n2946 = ~n2945;
  assign n2973 = n2974 & n2975;
  assign n2930 = ~n2976;
  assign n2971 = ~n2979;
  assign n2977 = ~n2990;
  assign n2957 = ~n2999;
  assign n2993 = n3000 & n3001;
  assign n2991 = ~n3000;
  assign n1673 = ~n3019;
  assign n3005 = n3027 & n3028;
  assign n2329 = ~n2349;
  assign n2905 = n2946 & n2947;
  assign n2948 = n2971 & n2972;
  assign n2951 = ~n2973;
  assign n2954 = n2977 & n2978;
  assign n2980 = n2991 & n2992;
  assign n2915 = ~n2993;
  assign n2982 = n3005 ^ n3006;
  assign n3007 = ~n3005;
  assign n2928 = n2948 ^ n2949;
  assign n2934 = n2954 ^ n2955;
  assign n2950 = ~n2948;
  assign n2956 = ~n2954;
  assign n2899 = ~n2980;
  assign n1582 = n2981 ^ n2982;
  assign n3002 = n3007 & n3008;
  assign n2906 = n72 ^ n2928;
  assign n2918 = n2934 ^ n2935;
  assign n2939 = n2950 & n2951;
  assign n2952 = n2956 & n2957;
  assign n78362 = n2960 ^ n1582;
  assign n2963 = n2915 & n2899;
  assign n2953 = n1582 & n1551;
  assign n2965 = n1582 & n1625;
  assign n2961 = ~n1582;
  assign n2983 = ~n3002;
  assign n909 = n2905 ^ n2906;
  assign n2843 = n2906 & n2905;
  assign n2911 = n2918 & n87;
  assign n2909 = ~n2918;
  assign n2929 = ~n2939;
  assign n2936 = ~n2952;
  assign n2938 = n2953 ^ n1610;
  assign n2926 = n2961 & n2962;
  assign n2913 = ~n2963;
  assign n2958 = n2961 & n2964;
  assign n1649 = ~n2965;
  assign n2966 = n2983 & n2984;
  assign n2264 = ~n909;
  assign n2907 = n2909 & n2910;
  assign n2871 = ~n2911;
  assign n2869 = n2929 & n2930;
  assign n2912 = n2936 & n2937;
  assign n2931 = n2938 & n2873;
  assign n2855 = ~n2938;
  assign n1628 = ~n2958;
  assign n2941 = n2966 ^ n1583;
  assign n2967 = ~n2966;
  assign n2893 = ~n2907;
  assign n2900 = n2912 ^ n2913;
  assign n2894 = ~n2869;
  assign n2914 = ~n2912;
  assign n2875 = ~n2931;
  assign n2919 = n2855 & n2932;
  assign n2927 = n2940 ^ n2941;
  assign n2959 = n2967 & n2968;
  assign n2888 = n2893 & n2894;
  assign n2868 = n2893 & n2871;
  assign n2897 = n2900 & n86;
  assign n2895 = ~n2900;
  assign n2908 = n2914 & n2915;
  assign n2858 = ~n2919;
  assign n78361 = n2926 ^ n2927;
  assign n2921 = n2927 & n2933;
  assign n2887 = n2927 & n2926;
  assign n1544 = ~n2927;
  assign n2942 = ~n2959;
  assign n2852 = n2868 ^ n2869;
  assign n2870 = ~n2888;
  assign n2889 = n2895 & n2896;
  assign n2824 = ~n2897;
  assign n2898 = ~n2908;
  assign n2901 = n1544 & n1523;
  assign n2916 = n1544 & n2920;
  assign n1568 = ~n2921;
  assign n2891 = ~n2887;
  assign n2922 = n2942 & n2943;
  assign n2185 = n2843 ^ n2852;
  assign n2816 = n2852 & n2843;
  assign n2844 = ~n2852;
  assign n2845 = n2870 & n2871;
  assign n2854 = ~n2889;
  assign n2872 = n2898 & n2899;
  assign n2890 = n2901 ^ n1583;
  assign n1599 = ~n2916;
  assign n2902 = n2922 ^ n2923;
  assign n2924 = ~n2922;
  assign n2164 = n2843 ^ n2844;
  assign n2853 = ~n2845;
  assign n2865 = n2854 & n2824;
  assign n2856 = n2872 ^ n2873;
  assign n2874 = ~n2872;
  assign n2880 = n2890 & n2829;
  assign n2803 = ~n2890;
  assign n1596 = n1599 & n1568;
  assign n1485 = n1515 ^ n2902;
  assign n2917 = n2924 & n2925;
  assign n2847 = n2853 & n2854;
  assign n2836 = n2855 ^ n2856;
  assign n2846 = ~n2865;
  assign n2866 = n2874 & n2875;
  assign n2876 = n2803 & n2879;
  assign n2831 = ~n2880;
  assign n78360 = n2887 ^ n1485;
  assign n2834 = n1485 & n2891;
  assign n2867 = n1485 & n1471;
  assign n2881 = n1485 & n2892;
  assign n2882 = ~n1485;
  assign n2903 = ~n2917;
  assign n2827 = n2836 & n85;
  assign n2817 = n2845 ^ n2846;
  assign n2823 = ~n2847;
  assign n2825 = ~n2836;
  assign n2857 = ~n2866;
  assign n2859 = n2867 ^ n1515;
  assign n2806 = ~n2876;
  assign n1535 = ~n2881;
  assign n2877 = n2882 & n2883;
  assign n2884 = n2903 & n2904;
  assign n2796 = n2816 ^ n2817;
  assign n2779 = n2823 & n2824;
  assign n2819 = n2825 & n2826;
  assign n2781 = ~n2827;
  assign n2818 = ~n2817;
  assign n2828 = n2857 & n2858;
  assign n2848 = n2859 & n2860;
  assign n2849 = ~n2859;
  assign n1504 = ~n2877;
  assign n2862 = n2884 ^ n1415;
  assign n2885 = ~n2884;
  assign n78316 = n2796 ^ n78348;
  assign n2659 = n2796 & n78348;
  assign n2753 = n2818 & n2816;
  assign n2802 = ~n2779;
  assign n2801 = ~n2819;
  assign n2804 = n2828 ^ n2829;
  assign n2830 = ~n2828;
  assign n2788 = ~n2848;
  assign n2837 = n2849 & n2850;
  assign n1532 = n1535 & n1504;
  assign n1393 = n2861 ^ n2862;
  assign n2878 = n2885 & n2886;
  assign n2772 = ~n78316;
  assign n2797 = n2801 & n2802;
  assign n2778 = n2801 & n2781;
  assign n2756 = n2803 ^ n2804;
  assign n2820 = n2830 & n2831;
  assign n2762 = ~n2837;
  assign n2821 = n1393 & n1327;
  assign n2838 = n1393 & n2851;
  assign n2815 = n1393 & n2834;
  assign n2835 = ~n1393;
  assign n2863 = ~n2878;
  assign n2747 = n2772 & n2773;
  assign n2754 = n2778 ^ n2779;
  assign n2784 = n2756 & n84;
  assign n2780 = ~n2797;
  assign n2782 = ~n2756;
  assign n2805 = ~n2820;
  assign n2785 = n2788 & n2762;
  assign n2736 = n2821 ^ n1415;
  assign n78359 = n2834 ^ n2835;
  assign n2832 = n2835 & n1444;
  assign n1479 = ~n2838;
  assign n2810 = ~n2815;
  assign n2840 = n2863 & n2864;
  assign n2727 = n2747 ^ n2748;
  assign n2720 = n2747 ^ n2749;
  assign n2742 = n2753 ^ n2754;
  assign n2699 = n2754 & n2753;
  assign n2755 = n2780 & n2781;
  assign n2774 = n2782 & n2783;
  assign n2734 = ~n2784;
  assign n2786 = n2805 & n2806;
  assign n2799 = n2736 & n2807;
  assign n2798 = ~n2736;
  assign n1447 = ~n2832;
  assign n1375 = n2839 ^ n2840;
  assign n2841 = ~n2840;
  assign n627 = n295 ^ n2720;
  assign n2694 = n2727 & n2728;
  assign n2473 = n2720 & n295;
  assign n2731 = n2742 & n78347;
  assign n2729 = ~n2742;
  assign n2702 = ~n2699;
  assign n2732 = n2755 ^ n2756;
  assign n2758 = ~n2755;
  assign n2757 = ~n2774;
  assign n2669 = n2785 ^ n2786;
  assign n2787 = ~n2786;
  assign n2791 = n2798 & n2709;
  assign n2738 = ~n2799;
  assign n78358 = n2815 ^ n1375;
  assign n2800 = n1375 & n1349;
  assign n2812 = n1375 & n2822;
  assign n2809 = ~n1375;
  assign n2833 = n2841 & n2842;
  assign n2580 = n2694 ^ n2695;
  assign n2698 = n2694 & n2695;
  assign n633 = ~n627;
  assign n2696 = ~n2694;
  assign n2721 = n2729 & n2730;
  assign n2704 = ~n2731;
  assign n2700 = n84 ^ n2732;
  assign n2750 = n2757 & n2758;
  assign n2759 = n2669 & n2766;
  assign n2760 = ~n2669;
  assign n2775 = n2787 & n2788;
  assign n2711 = ~n2791;
  assign n2789 = n2800 ^ n1395;
  assign n2764 = n2809 & n2810;
  assign n2808 = n2809 & n2811;
  assign n1420 = ~n2812;
  assign n2813 = ~n2833;
  assign n2690 = n2696 & n2697;
  assign n2567 = ~n2698;
  assign n2681 = n2699 ^ n2700;
  assign n2703 = n2704 & n2659;
  assign n2684 = ~n2721;
  assign n2701 = ~n2700;
  assign n2733 = ~n2750;
  assign n2707 = ~n2759;
  assign n2751 = n2760 & n83;
  assign n2761 = ~n2775;
  assign n2776 = n2789 & n2676;
  assign n2647 = ~n2789;
  assign n1384 = ~n2808;
  assign n2793 = n2813 & n2814;
  assign n2666 = n2681 & n2682;
  assign n2597 = ~n2690;
  assign n2667 = ~n2681;
  assign n2639 = n2701 & n2702;
  assign n2683 = ~n2703;
  assign n2691 = n2684 & n2704;
  assign n2705 = n2733 & n2734;
  assign n2671 = ~n2751;
  assign n2735 = n2761 & n2762;
  assign n2678 = ~n2776;
  assign n2767 = n2647 & n2777;
  assign n1417 = n1420 & n1384;
  assign n1292 = n2792 ^ n2793;
  assign n2794 = ~n2793;
  assign n2613 = ~n2666;
  assign n2658 = n2667 & n2565;
  assign n2610 = n2683 & n2684;
  assign n2642 = ~n2639;
  assign n2660 = ~n2691;
  assign n2668 = n83 ^ n2705;
  assign n2706 = ~n2705;
  assign n2708 = n2735 ^ n2736;
  assign n2737 = ~n2735;
  assign n2650 = ~n2767;
  assign n2752 = n1292 & n1205;
  assign n2768 = n1292 & n1331;
  assign n2765 = ~n1292;
  assign n2790 = n2794 & n2795;
  assign n2637 = ~n2658;
  assign n78315 = n2659 ^ n2660;
  assign n2636 = ~n2610;
  assign n2640 = n2668 ^ n2669;
  assign n2692 = n2706 & n2707;
  assign n2644 = n2708 ^ n2709;
  assign n2722 = n2737 & n2738;
  assign n2739 = n2752 ^ n1320;
  assign n78357 = n2764 ^ n2765;
  assign n1353 = ~n2768;
  assign n2763 = n2765 & n2769;
  assign n2713 = n2765 & n2764;
  assign n2770 = ~n2790;
  assign n2633 = n2636 & n2637;
  assign n2609 = n2637 & n2613;
  assign n2611 = n78315 & n2638;
  assign n2547 = n2639 ^ n2640;
  assign n1652 = ~n78315;
  assign n2641 = ~n2640;
  assign n2674 = n2644 & n82;
  assign n2670 = ~n2692;
  assign n2672 = ~n2644;
  assign n2710 = ~n2722;
  assign n2725 = n2739 & n2740;
  assign n2723 = ~n2739;
  assign n1334 = ~n2763;
  assign n2744 = n2770 & n2771;
  assign n1585 = n2609 ^ n2610;
  assign n2581 = n2611 ^ n78347;
  assign n2614 = n2547 & n2503;
  assign n2612 = ~n2633;
  assign n2615 = ~n2547;
  assign n2586 = n2641 & n2642;
  assign n2643 = n2670 & n2671;
  assign n2661 = n2672 & n2673;
  assign n2619 = ~n2674;
  assign n2675 = n2710 & n2711;
  assign n2715 = n2723 & n2724;
  assign n2626 = ~n2725;
  assign n1256 = n2743 ^ n2744;
  assign n2745 = ~n2744;
  assign n2563 = n2580 ^ n2581;
  assign n2582 = n2581 & n2597;
  assign n2564 = n1585 & n2598;
  assign n2513 = n1585 & n78315;
  assign n1613 = ~n1585;
  assign n2583 = n2612 & n2613;
  assign n2584 = ~n2614;
  assign n2604 = n2615 & n2616;
  assign n2589 = ~n2586;
  assign n2617 = n2643 ^ n2644;
  assign n2645 = ~n2643;
  assign n2646 = ~n2661;
  assign n2648 = n2675 ^ n2676;
  assign n2677 = ~n2675;
  assign n2596 = ~n2715;
  assign n2693 = n1256 & n1228;
  assign n2717 = n1256 & n2726;
  assign n2714 = ~n1256;
  assign n2741 = n2745 & n2746;
  assign n2546 = n2563 & n294;
  assign n2535 = n2564 ^ n2565;
  assign n2544 = ~n2563;
  assign n78314 = n1613 ^ n78315;
  assign n2566 = ~n2582;
  assign n2548 = n2583 ^ n2503;
  assign n2585 = ~n2583;
  assign n2550 = ~n2604;
  assign n2587 = n82 ^ n2617;
  assign n2634 = n2645 & n2646;
  assign n2629 = n2647 ^ n2648;
  assign n2662 = n2677 & n2678;
  assign n2685 = n2626 & n2596;
  assign n2679 = n2693 ^ n1293;
  assign n78372 = n2713 ^ n2714;
  assign n2712 = n2714 & n2716;
  assign n2652 = n2714 & n2713;
  assign n1310 = ~n2717;
  assign n2718 = ~n2741;
  assign n2530 = n2535 & n2536;
  assign n2537 = n2544 & n2545;
  assign n2495 = ~n2546;
  assign n1487 = n2547 ^ n2548;
  assign n2528 = ~n2535;
  assign n2463 = n2566 & n2567;
  assign n2575 = n2584 & n2585;
  assign n2568 = n2586 ^ n2587;
  assign n2588 = ~n2587;
  assign n2622 = n2629 & n81;
  assign n2618 = ~n2634;
  assign n2620 = ~n2629;
  assign n2649 = ~n2662;
  assign n2663 = n2679 & n2556;
  assign n2624 = ~n2685;
  assign n2523 = ~n2679;
  assign n1277 = ~n2712;
  assign n2687 = n2718 & n2719;
  assign n2516 = n2528 & n2529;
  assign n2465 = ~n2530;
  assign n2502 = n1487 & n2531;
  assign n2429 = n1487 & n2513;
  assign n2527 = ~n2537;
  assign n1549 = ~n1487;
  assign n2505 = ~n2463;
  assign n2552 = n2568 & n2569;
  assign n2549 = ~n2575;
  assign n2551 = ~n2568;
  assign n2508 = n2588 & n2589;
  assign n2539 = n2618 & n2619;
  assign n2605 = n2620 & n2621;
  assign n2554 = ~n2622;
  assign n2623 = n2649 & n2650;
  assign n2558 = ~n2663;
  assign n2654 = n2523 & n2664;
  assign n1307 = n1310 & n1277;
  assign n1157 = n2686 ^ n2687;
  assign n2688 = ~n2687;
  assign n2363 = n2502 ^ n2503;
  assign n78313 = n2513 ^ n1549;
  assign n2504 = ~n2516;
  assign n2514 = n2527 & n2473;
  assign n2515 = n2527 & n2495;
  assign n2466 = n2549 & n2550;
  assign n2538 = n2551 & n2392;
  assign n2476 = ~n2552;
  assign n2511 = ~n2508;
  assign n2590 = ~n2539;
  assign n2591 = ~n2605;
  assign n2520 = n2623 ^ n2624;
  assign n2625 = ~n2623;
  assign n2526 = ~n2654;
  assign n2635 = n1157 & n1140;
  assign n2655 = n1157 & n2665;
  assign n2653 = ~n1157;
  assign n2680 = n2688 & n2689;
  assign n2460 = n2363 & n2472;
  assign n2461 = ~n2363;
  assign n2493 = n2504 & n2505;
  assign n2462 = n2465 & n2504;
  assign n2494 = ~n2514;
  assign n2474 = ~n2515;
  assign n2517 = ~n2466;
  assign n2518 = ~n2538;
  assign n2576 = n2590 & n2591;
  assign n2577 = n2591 & n2554;
  assign n2594 = n2520 & n80;
  assign n2592 = ~n2520;
  assign n2606 = n2625 & n2626;
  assign n2627 = n2635 ^ n1183;
  assign n78371 = n2652 ^ n2653;
  assign n1239 = ~n2655;
  assign n2651 = n2653 & n1237;
  assign n2561 = n2653 & n2652;
  assign n2656 = ~n2680;
  assign n2381 = ~n2460;
  assign n2446 = n2461 & n2410;
  assign n2421 = n2462 ^ n2463;
  assign n2431 = n2473 ^ n2474;
  assign n2464 = ~n2493;
  assign n2420 = n2494 & n2495;
  assign n2506 = n2517 & n2518;
  assign n2507 = n2518 & n2476;
  assign n2553 = ~n2576;
  assign n2540 = ~n2577;
  assign n2578 = n2592 & n2593;
  assign n2481 = ~n2594;
  assign n2595 = ~n2606;
  assign n2607 = n2627 & n2486;
  assign n2441 = ~n2627;
  assign n1211 = ~n2651;
  assign n2630 = n2656 & n2657;
  assign n2379 = n2420 ^ n2421;
  assign n2423 = n2421 & n2430;
  assign n616 = n2431 ^ n627;
  assign n2422 = ~n2446;
  assign n2424 = ~n2421;
  assign n2447 = n2464 & n2465;
  assign n2432 = ~n2431;
  assign n2390 = ~n2420;
  assign n2475 = ~n2506;
  assign n2467 = ~n2507;
  assign n2509 = n2539 ^ n2540;
  assign n2519 = n2553 & n2554;
  assign n2522 = ~n2578;
  assign n2555 = n2595 & n2596;
  assign n2488 = ~n2607;
  assign n2599 = n2441 & n2608;
  assign n2601 = n2630 ^ n1125;
  assign n2631 = ~n2630;
  assign n2337 = n293 ^ n2379;
  assign n2389 = ~n2423;
  assign n2408 = n2424 & n293;
  assign n1381 = ~n616;
  assign n2336 = n2432 & n627;
  assign n2409 = ~n2447;
  assign n1428 = n2466 ^ n2467;
  assign n2448 = n2475 & n2476;
  assign n2477 = n2508 ^ n2509;
  assign n2479 = n2519 ^ n2520;
  assign n2510 = ~n2509;
  assign n2521 = ~n2519;
  assign n2524 = n2555 ^ n2556;
  assign n2557 = ~n2555;
  assign n2443 = ~n2599;
  assign n1092 = n2600 ^ n2601;
  assign n2628 = n2631 & n2632;
  assign n603 = n2336 ^ n2337;
  assign n2223 = n2337 & n2336;
  assign n2382 = n2389 & n2390;
  assign n2352 = ~n2408;
  assign n2362 = n2409 ^ n2410;
  assign n2407 = n2422 & n2409;
  assign n78312 = n2429 ^ n1428;
  assign n1521 = ~n1428;
  assign n2450 = ~n2448;
  assign n2468 = n2477 & n2478;
  assign n2436 = n80 ^ n2479;
  assign n2449 = ~n2477;
  assign n2435 = n2510 & n2511;
  assign n2512 = n2521 & n2522;
  assign n2394 = n2523 ^ n2524;
  assign n2541 = n2557 & n2558;
  assign n2542 = n1092 & n1074;
  assign n2570 = n1092 & n2579;
  assign n2562 = ~n1092;
  assign n2602 = ~n2628;
  assign n1321 = ~n603;
  assign n2268 = n2362 ^ n2363;
  assign n2351 = ~n2382;
  assign n2380 = ~n2407;
  assign n2391 = n1521 & n2433;
  assign n2350 = n1521 & n2429;
  assign n2367 = n2435 ^ n2436;
  assign n2411 = n2448 ^ n2449;
  assign n2370 = n2436 & n2435;
  assign n2451 = ~n2468;
  assign n2452 = n2449 & n2340;
  assign n2484 = n2394 & n95;
  assign n2480 = ~n2512;
  assign n2482 = ~n2394;
  assign n2525 = ~n2541;
  assign n2359 = n2542 ^ n2543;
  assign n78370 = n2561 ^ n2562;
  assign n2559 = n2562 & n1186;
  assign n1188 = ~n2570;
  assign n2491 = n2562 & n2561;
  assign n2571 = n2602 & n2603;
  assign n2314 = n2268 & n2338;
  assign n2304 = n2351 & n2352;
  assign n2315 = ~n2268;
  assign n2253 = n2380 & n2381;
  assign n2364 = n2391 ^ n2392;
  assign n1401 = n2411 ^ n2340;
  assign n2343 = ~n2367;
  assign n2373 = ~n2370;
  assign n2434 = n2450 & n2451;
  assign n2413 = ~n2452;
  assign n2437 = n2480 & n2481;
  assign n2469 = n2482 & n2483;
  assign n2396 = ~n2484;
  assign n2485 = n2525 & n2526;
  assign n1161 = ~n2559;
  assign n2532 = n2571 ^ n2572;
  assign n2573 = ~n2571;
  assign n2267 = n292 ^ n2304;
  assign n2292 = ~n2314;
  assign n2305 = n2315 & n292;
  assign n2293 = ~n2304;
  assign n2306 = ~n2253;
  assign n2353 = n2364 & n2365;
  assign n2339 = n1401 & n2383;
  assign n2278 = n1401 & n2350;
  assign n2354 = ~n2364;
  assign n1437 = ~n1401;
  assign n2412 = ~n2434;
  assign n2393 = n95 ^ n2437;
  assign n2438 = ~n2437;
  assign n2439 = ~n2469;
  assign n2440 = n2485 ^ n2486;
  assign n2487 = ~n2485;
  assign n1042 = n2532 ^ n1076;
  assign n2560 = n2573 & n2574;
  assign n2224 = n2267 ^ n2268;
  assign n2279 = n2292 & n2293;
  assign n2252 = ~n2305;
  assign n2226 = n2339 ^ n2340;
  assign n78311 = n2350 ^ n1437;
  assign n2270 = ~n2353;
  assign n2341 = n2354 & n2355;
  assign n2371 = n2393 ^ n2394;
  assign n2366 = n2412 & n2413;
  assign n2425 = n2438 & n2439;
  assign n2414 = n2440 ^ n2441;
  assign n2470 = n2487 & n2488;
  assign n2471 = n1042 & n1020;
  assign n2496 = n1042 & n1093;
  assign n2492 = ~n1042;
  assign n2533 = ~n2560;
  assign n591 = n2223 ^ n2224;
  assign n2084 = n2224 & n2223;
  assign n2251 = ~n2279;
  assign n2296 = n2226 & n2188;
  assign n2294 = ~n2226;
  assign n2307 = ~n2341;
  assign n2316 = n2366 ^ n2367;
  assign n2344 = n2370 ^ n2371;
  assign n2369 = n2366 & n2384;
  assign n2372 = ~n2371;
  assign n2368 = ~n2366;
  assign n2399 = n2414 & n94;
  assign n2395 = ~n2425;
  assign n2397 = ~n2414;
  assign n2442 = ~n2470;
  assign n2444 = n2471 ^ n1076;
  assign n78369 = n2491 ^ n2492;
  assign n1130 = ~n2496;
  assign n2489 = n2492 & n2497;
  assign n2459 = n2492 & n2491;
  assign n2499 = n2533 & n2534;
  assign n1294 = ~n591;
  assign n2088 = ~n2084;
  assign n2118 = n2251 & n2252;
  assign n2280 = n2294 & n2295;
  assign n2227 = ~n2296;
  assign n2297 = n2306 & n2307;
  assign n2298 = n2270 & n2307;
  assign n1368 = n2316 ^ n2237;
  assign n2318 = n2344 & n2345;
  assign n2319 = ~n2344;
  assign n2356 = n2368 & n2237;
  assign n2342 = ~n2369;
  assign n2271 = n2372 & n2373;
  assign n2309 = n2395 & n2396;
  assign n2385 = n2397 & n2398;
  assign n2321 = ~n2399;
  assign n2400 = n2442 & n2443;
  assign n2427 = n2444 & n2285;
  assign n2257 = ~n2444;
  assign n1096 = ~n2489;
  assign n2453 = ~n2459;
  assign n976 = n2498 ^ n2499;
  assign n2500 = ~n2499;
  assign n2167 = ~n2118;
  assign n78310 = n2278 ^ n1368;
  assign n2190 = ~n2280;
  assign n2269 = ~n2297;
  assign n2254 = ~n2298;
  assign n1378 = ~n1368;
  assign n2214 = ~n2318;
  assign n2308 = n2319 & n2169;
  assign n2317 = n2342 & n2343;
  assign n2300 = ~n2356;
  assign n2274 = ~n2271;
  assign n2357 = ~n2309;
  assign n2358 = ~n2385;
  assign n2360 = n2400 ^ n2401;
  assign n2404 = n2400 & n2401;
  assign n2402 = ~n2400;
  assign n2415 = n2257 & n2426;
  assign n2287 = ~n2427;
  assign n2335 = n976 & n2453;
  assign n78368 = n2459 ^ n976;
  assign n2428 = n976 & n957;
  assign n2454 = n976 & n1032;
  assign n2455 = ~n976;
  assign n2490 = n2500 & n2501;
  assign n2229 = n2253 ^ n2254;
  assign n2225 = n2269 & n2270;
  assign n2236 = n1378 & n2281;
  assign n2186 = n1378 & n2278;
  assign n2256 = ~n2308;
  assign n2299 = ~n2317;
  assign n2347 = n2357 & n2358;
  assign n2348 = n2358 & n2321;
  assign n2346 = n2359 ^ n2360;
  assign n2386 = n2402 & n2403;
  assign n2374 = ~n2404;
  assign n2260 = ~n2415;
  assign n2405 = n2428 ^ n1010;
  assign n2328 = ~n2335;
  assign n1068 = ~n2454;
  assign n2445 = n2455 & n2456;
  assign n2457 = ~n2490;
  assign n2187 = n2225 ^ n2226;
  assign n2211 = n2229 & n291;
  assign n2147 = n2236 ^ n2237;
  assign n2209 = ~n2229;
  assign n2228 = ~n2225;
  assign n2238 = n2256 & n2214;
  assign n2239 = n2299 & n2300;
  assign n2324 = n2346 & n93;
  assign n2320 = ~n2347;
  assign n2310 = ~n2348;
  assign n2322 = ~n2346;
  assign n2361 = n2374 & n2359;
  assign n2326 = ~n2386;
  assign n2387 = n2405 & n2220;
  assign n2177 = ~n2405;
  assign n1035 = ~n2445;
  assign n2416 = n2457 & n2458;
  assign n2051 = n2187 ^ n2188;
  assign n2196 = n2147 & n2207;
  assign n2197 = n2209 & n2210;
  assign n2127 = ~n2211;
  assign n2208 = n2227 & n2228;
  assign n2195 = ~n2147;
  assign n1241 = n2238 ^ n2239;
  assign n2255 = ~n2239;
  assign n2272 = n2309 ^ n2310;
  assign n2242 = n2320 & n2321;
  assign n2311 = n2322 & n2323;
  assign n2244 = ~n2324;
  assign n2325 = ~n2361;
  assign n2222 = ~n2387;
  assign n2375 = n2177 & n2388;
  assign n2376 = n2416 ^ n2417;
  assign n2418 = ~n2416;
  assign n2072 = ~n2051;
  assign n2191 = n2195 & n2108;
  assign n2149 = ~n2196;
  assign n2166 = ~n2197;
  assign n2189 = ~n2208;
  assign n2168 = n1241 & n2212;
  assign n2093 = n1241 & n2186;
  assign n1314 = ~n1241;
  assign n2240 = n2255 & n2256;
  assign n2132 = n2271 ^ n2272;
  assign n2273 = ~n2272;
  assign n2282 = ~n2242;
  assign n2283 = ~n2311;
  assign n2284 = n2325 & n2326;
  assign n2180 = ~n2375;
  assign n941 = n2376 ^ n977;
  assign n2406 = n2418 & n2419;
  assign n2157 = n2166 & n2167;
  assign n2158 = n2166 & n2127;
  assign n2150 = n2168 ^ n2169;
  assign n78309 = n2186 ^ n1314;
  assign n2146 = n2189 & n2190;
  assign n2111 = ~n2191;
  assign n2097 = ~n2093;
  assign n2213 = ~n2240;
  assign n2230 = n2132 & n2074;
  assign n2231 = ~n2132;
  assign n2198 = n2273 & n2274;
  assign n2275 = n2282 & n2283;
  assign n2241 = n2283 & n2244;
  assign n2258 = n2284 ^ n2285;
  assign n2286 = ~n2284;
  assign n78367 = n2335 ^ n941;
  assign n2301 = n941 & n844;
  assign n2330 = n941 & n2349;
  assign n2327 = ~n941;
  assign n2377 = ~n2406;
  assign n2107 = n2146 ^ n2147;
  assign n2131 = n2150 & n2151;
  assign n2126 = ~n2157;
  assign n2119 = ~n2158;
  assign n2129 = ~n2150;
  assign n2148 = ~n2146;
  assign n2170 = n2213 & n2214;
  assign n2172 = ~n2230;
  assign n2215 = n2231 & n2232;
  assign n2199 = n2241 ^ n2242;
  assign n2201 = ~n2198;
  assign n2192 = n2257 ^ n2258;
  assign n2243 = ~n2275;
  assign n2276 = n2286 & n2287;
  assign n2142 = n2301 ^ n977;
  assign n2250 = n2327 & n2328;
  assign n2312 = n2327 & n2329;
  assign n1004 = ~n2330;
  assign n2331 = n2377 & n2378;
  assign n2083 = n2107 ^ n2108;
  assign n2085 = n2118 ^ n2119;
  assign n2094 = n2126 & n2127;
  assign n2120 = n2129 & n2130;
  assign n2041 = ~n2131;
  assign n2128 = n2148 & n2149;
  assign n2133 = n2170 ^ n2074;
  assign n2171 = ~n2170;
  assign n2173 = n2198 ^ n2199;
  assign n2135 = ~n2215;
  assign n2218 = n2192 & n92;
  assign n2200 = ~n2199;
  assign n2233 = n2243 & n2244;
  assign n2216 = ~n2192;
  assign n2259 = ~n2276;
  assign n2263 = n2142 & n2104;
  assign n2261 = ~n2142;
  assign n965 = ~n2312;
  assign n2288 = n2331 ^ n2332;
  assign n2334 = n2331 & n2290;
  assign n2333 = ~n2331;
  assign n2070 = n2083 & n289;
  assign n587 = n2084 ^ n2085;
  assign n2068 = ~n2083;
  assign n2050 = n290 ^ n2094;
  assign n2096 = n2094 & n2109;
  assign n2087 = ~n2085;
  assign n2095 = ~n2094;
  assign n2076 = ~n2120;
  assign n2110 = ~n2128;
  assign n1246 = n2132 ^ n2133;
  assign n2159 = n2171 & n2172;
  assign n2161 = n2173 & n2174;
  assign n2160 = ~n2173;
  assign n2113 = n2200 & n2201;
  assign n2202 = n2216 & n2217;
  assign n2137 = ~n2218;
  assign n2176 = ~n2233;
  assign n2219 = n2259 & n2260;
  assign n2245 = n2261 & n2262;
  assign n2144 = ~n2263;
  assign n1001 = n1004 & n965;
  assign n931 = n877 ^ n2288;
  assign n2313 = n2333 & n2303;
  assign n2302 = ~n2334;
  assign n2015 = n2050 ^ n2051;
  assign n2052 = n2068 & n2069;
  assign n1973 = ~n2070;
  assign n1194 = ~n587;
  assign n2014 = n2087 & n2088;
  assign n78324 = n2093 ^ n1246;
  assign n2086 = n2095 & n290;
  assign n2071 = ~n2096;
  assign n2089 = n2041 & n2076;
  assign n2046 = n2110 & n2111;
  assign n2073 = n1246 & n2112;
  assign n1258 = ~n1246;
  assign n2134 = ~n2159;
  assign n2152 = n2160 & n2005;
  assign n2056 = ~n2161;
  assign n2116 = ~n2113;
  assign n2153 = n2176 ^ n2192;
  assign n2175 = ~n2202;
  assign n2178 = n2219 ^ n2220;
  assign n2221 = ~n2219;
  assign n2106 = ~n2245;
  assign n78366 = n2250 ^ n931;
  assign n2246 = n931 & n2264;
  assign n2155 = n931 & n2250;
  assign n848 = ~n931;
  assign n2291 = n2302 & n2303;
  assign n2289 = ~n2313;
  assign n578 = n2014 ^ n2015;
  assign n2001 = ~n2052;
  assign n2053 = n2071 & n2072;
  assign n2044 = n2073 ^ n2074;
  assign n2034 = ~n2014;
  assign n2036 = ~n2086;
  assign n2047 = ~n2089;
  assign n2075 = ~n2046;
  assign n2033 = n1258 & n2097;
  assign n2077 = n2134 & n2135;
  assign n2099 = ~n2152;
  assign n2114 = n92 ^ n2153;
  assign n2162 = n2175 & n2176;
  assign n2059 = n2177 ^ n2178;
  assign n2203 = n2221 & n2222;
  assign n2204 = n848 & n785;
  assign n897 = ~n2246;
  assign n2234 = n848 & n909;
  assign n2277 = n2289 & n2290;
  assign n2265 = ~n2291;
  assign n1141 = ~n578;
  assign n1952 = n2015 & n2034;
  assign n2016 = n2001 & n1973;
  assign n2037 = n2044 & n2045;
  assign n2018 = n2046 ^ n2047;
  assign n2035 = ~n2053;
  assign n2038 = ~n2044;
  assign n2054 = n2075 & n2076;
  assign n2091 = n2113 ^ n2114;
  assign n2098 = ~n2077;
  assign n2117 = n2099 & n2056;
  assign n2115 = ~n2114;
  assign n2140 = n2059 & n91;
  assign n2136 = ~n2162;
  assign n2138 = ~n2059;
  assign n2179 = ~n2203;
  assign n2193 = n2204 ^ n877;
  assign n912 = ~n2234;
  assign n2249 = n2265 & n2266;
  assign n2247 = ~n2277;
  assign n1985 = ~n2016;
  assign n2010 = n2018 & n288;
  assign n1984 = n2035 & n2036;
  assign n1971 = ~n2037;
  assign n2017 = n2038 & n2039;
  assign n2008 = ~n2018;
  assign n2040 = ~n2054;
  assign n2081 = n2091 & n1947;
  assign n2090 = n2098 & n2099;
  assign n2079 = ~n2091;
  assign n2021 = n2115 & n2116;
  assign n2078 = ~n2117;
  assign n2100 = n2136 & n2137;
  assign n2121 = n2138 & n2139;
  assign n2061 = ~n2140;
  assign n2141 = n2179 & n2180;
  assign n2183 = n2193 & n2194;
  assign n2181 = ~n2193;
  assign n2235 = n2247 & n2248;
  assign n2206 = ~n2249;
  assign n1953 = n1984 ^ n1985;
  assign n2003 = n2008 & n2009;
  assign n1911 = ~n2010;
  assign n2002 = ~n1984;
  assign n1999 = ~n2017;
  assign n1954 = n2040 & n2041;
  assign n1143 = n2077 ^ n2078;
  assign n2057 = n2079 & n2080;
  assign n2020 = ~n2081;
  assign n2055 = ~n2090;
  assign n2024 = ~n2021;
  assign n2058 = n91 ^ n2100;
  assign n2102 = ~n2100;
  assign n2101 = ~n2121;
  assign n2103 = n2141 ^ n2142;
  assign n2143 = ~n2141;
  assign n2163 = n2181 & n2182;
  assign n2067 = ~n2183;
  assign n2205 = ~n2235;
  assign n555 = n1952 ^ n1953;
  assign n1904 = n1953 & n1952;
  assign n1987 = n2001 & n2002;
  assign n1988 = n1971 & n1999;
  assign n1944 = ~n2003;
  assign n2000 = ~n1954;
  assign n78323 = n2033 ^ n1143;
  assign n1969 = n1143 & n2033;
  assign n2007 = n2055 & n2056;
  assign n1226 = ~n1143;
  assign n1990 = ~n2057;
  assign n2022 = n2058 ^ n2059;
  assign n2092 = n2101 & n2102;
  assign n1994 = n2103 ^ n2104;
  assign n2122 = n2143 & n2144;
  assign n2032 = ~n2163;
  assign n800 = n2205 & n2206;
  assign n1077 = ~n555;
  assign n1907 = ~n1904;
  assign n1974 = n1944 & n1911;
  assign n1972 = ~n1987;
  assign n1955 = ~n1988;
  assign n1986 = n1999 & n2000;
  assign n1929 = n2021 ^ n2022;
  assign n1980 = ~n1969;
  assign n2004 = n1226 & n2042;
  assign n2006 = n1990 & n2020;
  assign n2019 = ~n2007;
  assign n2023 = ~n2022;
  assign n2062 = n1994 & n2082;
  assign n2060 = ~n2092;
  assign n2063 = ~n1994;
  assign n2105 = ~n2122;
  assign n2123 = n2067 & n2032;
  assign n2145 = n800 & n2184;
  assign n2165 = n800 & n2185;
  assign n2156 = ~n800;
  assign n1882 = n1954 ^ n1955;
  assign n1939 = n1972 & n1973;
  assign n1940 = ~n1974;
  assign n1970 = ~n1986;
  assign n1978 = n2004 ^ n2005;
  assign n1992 = n1929 & n1958;
  assign n1134 = n2006 ^ n2007;
  assign n1991 = ~n1929;
  assign n2011 = n2019 & n2020;
  assign n1961 = n2023 & n2024;
  assign n2025 = n2060 & n2061;
  assign n2027 = ~n2062;
  assign n2048 = n2063 & n90;
  assign n2064 = n2105 & n2106;
  assign n2065 = ~n2123;
  assign n1967 = n2145 ^ n832;
  assign n78365 = n2155 ^ n2156;
  assign n2154 = n2156 & n2164;
  assign n2125 = ~n2165;
  assign n1923 = n1882 & n303;
  assign n1905 = n1939 ^ n1940;
  assign n1921 = ~n1882;
  assign n1943 = ~n1939;
  assign n78322 = n1969 ^ n1134;
  assign n1896 = n1970 & n1971;
  assign n1977 = n1978 & n1979;
  assign n1891 = n1134 & n1980;
  assign n1946 = n1134 & n1981;
  assign n1975 = ~n1978;
  assign n1982 = n1991 & n1889;
  assign n1932 = ~n1992;
  assign n1109 = ~n1134;
  assign n1989 = ~n2011;
  assign n1964 = ~n1961;
  assign n1993 = n90 ^ n2025;
  assign n2026 = ~n2025;
  assign n1996 = ~n2048;
  assign n2043 = n2064 ^ n2065;
  assign n2066 = ~n2064;
  assign n2124 = ~n2154;
  assign n546 = n1904 ^ n1905;
  assign n1914 = n1921 & n1922;
  assign n1864 = ~n1923;
  assign n1906 = ~n1905;
  assign n1925 = n1943 & n1944;
  assign n1926 = n1946 ^ n1947;
  assign n1941 = ~n1896;
  assign n1956 = n1975 & n1976;
  assign n1909 = ~n1977;
  assign n1960 = ~n1982;
  assign n1957 = n1989 & n1990;
  assign n1962 = n1993 ^ n1994;
  assign n2012 = n2026 & n2027;
  assign n2030 = n2043 & n89;
  assign n2028 = ~n2043;
  assign n2049 = n2066 & n2067;
  assign n880 = n2124 & n2125;
  assign n999 = ~n546;
  assign n1837 = n1906 & n1907;
  assign n1885 = ~n1914;
  assign n1910 = ~n1925;
  assign n1915 = n1926 & n1927;
  assign n1916 = ~n1926;
  assign n1942 = ~n1956;
  assign n1928 = n1957 ^ n1958;
  assign n1945 = n1961 ^ n1962;
  assign n1959 = ~n1957;
  assign n1963 = ~n1962;
  assign n1995 = ~n2012;
  assign n2013 = n2028 & n2029;
  assign n1938 = ~n2030;
  assign n2031 = ~n2049;
  assign n868 = ~n880;
  assign n1881 = n1910 & n1911;
  assign n1862 = ~n1915;
  assign n1913 = n1916 & n1917;
  assign n1012 = n1928 ^ n1929;
  assign n1924 = n1941 & n1942;
  assign n1930 = n1942 & n1909;
  assign n1934 = n1945 & n1832;
  assign n1899 = ~n1945;
  assign n1948 = n1959 & n1960;
  assign n1919 = n1963 & n1964;
  assign n1949 = n1995 & n1996;
  assign n1966 = ~n2013;
  assign n1997 = n2031 & n2032;
  assign n1860 = n1881 ^ n1882;
  assign n1886 = ~n1881;
  assign n1888 = n1012 & n1912;
  assign n1850 = n1012 & n1891;
  assign n1884 = ~n1913;
  assign n1083 = ~n1012;
  assign n1908 = ~n1924;
  assign n1897 = ~n1930;
  assign n1918 = n1899 & n1933;
  assign n1900 = ~n1934;
  assign n1931 = ~n1948;
  assign n1935 = ~n1919;
  assign n1965 = ~n1949;
  assign n1983 = n1966 & n1938;
  assign n1968 = n1997 ^ n1998;
  assign n1838 = n303 ^ n1860;
  assign n1872 = n1885 & n1886;
  assign n1819 = n1888 ^ n1889;
  assign n78321 = n1891 ^ n1083;
  assign n1868 = n1862 & n1884;
  assign n1887 = n1896 ^ n1897;
  assign n1869 = n1908 & n1909;
  assign n1878 = ~n1918;
  assign n1898 = n1931 & n1932;
  assign n1951 = n1965 & n1966;
  assign n1936 = n1967 ^ n1968;
  assign n1950 = ~n1983;
  assign n978 = n1837 ^ n1838;
  assign n1808 = n1838 & n1837;
  assign n1866 = n1819 & n1867;
  assign n1800 = n1868 ^ n1869;
  assign n1863 = ~n1872;
  assign n1865 = ~n1819;
  assign n1875 = n1887 & n302;
  assign n1873 = ~n1887;
  assign n1883 = ~n1869;
  assign n1876 = n1898 ^ n1899;
  assign n1901 = ~n1898;
  assign n1903 = n88 ^ n1936;
  assign n1920 = n1949 ^ n1950;
  assign n1937 = ~n1951;
  assign n962 = ~n978;
  assign n1846 = n1800 & n1851;
  assign n1828 = n1863 & n1864;
  assign n1852 = n1865 & n1840;
  assign n1821 = ~n1866;
  assign n1847 = ~n1800;
  assign n1870 = n1873 & n1874;
  assign n1823 = ~n1875;
  assign n980 = n1876 ^ n1832;
  assign n1871 = n1883 & n1884;
  assign n1892 = n1900 & n1901;
  assign n1833 = n1919 ^ n1920;
  assign n1879 = n1920 & n1935;
  assign n1902 = n1937 & n1938;
  assign n1802 = ~n1846;
  assign n1845 = n1847 & n301;
  assign n78320 = n1850 ^ n980;
  assign n1843 = ~n1828;
  assign n1841 = ~n1852;
  assign n1844 = ~n1870;
  assign n1023 = ~n980;
  assign n1861 = ~n1871;
  assign n1877 = ~n1892;
  assign n1895 = n1833 & n1804;
  assign n1880 = n1902 ^ n1903;
  assign n1893 = ~n1833;
  assign n1830 = n1843 & n1844;
  assign n1781 = ~n1845;
  assign n1827 = n1844 & n1823;
  assign n1831 = n1023 & n1853;
  assign n1817 = n1023 & n1850;
  assign n1839 = n1861 & n1862;
  assign n1854 = n1877 & n1878;
  assign n1793 = n1879 ^ n1880;
  assign n1890 = n1893 & n1894;
  assign n1856 = ~n1895;
  assign n1809 = n1827 ^ n1828;
  assign n1822 = ~n1830;
  assign n1824 = n1831 ^ n1832;
  assign n1818 = n1839 ^ n1840;
  assign n1813 = ~n1817;
  assign n1842 = ~n1839;
  assign n1834 = n1854 ^ n1804;
  assign n1859 = n1793 & n1766;
  assign n1855 = ~n1854;
  assign n1857 = ~n1793;
  assign n1836 = ~n1890;
  assign n522 = n1808 ^ n1809;
  assign n1746 = n1809 & n1808;
  assign n1805 = n1818 ^ n1819;
  assign n1799 = n1822 & n1823;
  assign n1810 = n1824 & n1825;
  assign n1811 = ~n1824;
  assign n955 = n1833 ^ n1834;
  assign n1829 = n1841 & n1842;
  assign n1848 = n1855 & n1856;
  assign n1849 = n1857 & n1858;
  assign n1795 = ~n1859;
  assign n1779 = n1799 ^ n1800;
  assign n1798 = n1805 & n300;
  assign n892 = ~n522;
  assign n1767 = ~n1746;
  assign n1796 = ~n1805;
  assign n1801 = ~n1799;
  assign n1772 = ~n1810;
  assign n1806 = n1811 & n1812;
  assign n78319 = n1817 ^ n955;
  assign n1803 = n955 & n1826;
  assign n882 = ~n955;
  assign n1820 = ~n1829;
  assign n1835 = ~n1848;
  assign n1816 = ~n1849;
  assign n1759 = n301 ^ n1779;
  assign n1788 = n1796 & n1797;
  assign n1740 = ~n1798;
  assign n1791 = n1801 & n1802;
  assign n1726 = n1803 ^ n1804;
  assign n1790 = ~n1806;
  assign n1778 = n882 & n1813;
  assign n1770 = n1820 & n1821;
  assign n1814 = n1835 & n1836;
  assign n833 = n1746 ^ n1759;
  assign n1736 = n1759 & n1767;
  assign n1747 = ~n1759;
  assign n1782 = n1726 & n1786;
  assign n1762 = ~n1788;
  assign n1780 = ~n1791;
  assign n1769 = n1790 & n1772;
  assign n1783 = ~n1726;
  assign n1784 = ~n1778;
  assign n1789 = ~n1770;
  assign n1792 = n1814 ^ n1766;
  assign n1815 = ~n1814;
  assign n821 = n1746 ^ n1747;
  assign n1719 = n1769 ^ n1770;
  assign n1760 = n1762 & n1740;
  assign n1761 = n1780 & n1781;
  assign n1728 = ~n1782;
  assign n1773 = n1783 & n1752;
  assign n1787 = n1789 & n1790;
  assign n852 = n1792 ^ n1793;
  assign n1807 = n1815 & n1816;
  assign n1737 = n1760 ^ n1761;
  assign n1749 = n1719 & n1764;
  assign n1750 = ~n1719;
  assign n1763 = ~n1761;
  assign n1753 = ~n1773;
  assign n78318 = n1778 ^ n852;
  assign n1755 = n852 & n1784;
  assign n1765 = n852 & n1785;
  assign n1771 = ~n1787;
  assign n886 = ~n852;
  assign n1794 = ~n1807;
  assign n1716 = n1736 ^ n1737;
  assign n1738 = ~n1737;
  assign n1721 = ~n1749;
  assign n1744 = n1750 & n299;
  assign n1748 = n1762 & n1763;
  assign n1707 = n1765 ^ n1766;
  assign n1751 = n1771 & n1772;
  assign n1774 = n1794 & n1795;
  assign n78284 = n1716 ^ n78316;
  assign n1717 = ~n1716;
  assign n1674 = n1738 & n1736;
  assign n1696 = ~n1744;
  assign n1741 = n1707 & n1687;
  assign n1739 = ~n1748;
  assign n1725 = n1751 ^ n1752;
  assign n1742 = ~n1707;
  assign n1754 = ~n1751;
  assign n804 = n1774 ^ n1775;
  assign n1776 = ~n1774;
  assign n1572 = ~n78284;
  assign n1587 = n1717 & n78316;
  assign n1677 = ~n1674;
  assign n1655 = n1725 ^ n1726;
  assign n1718 = n1739 & n1740;
  assign n1708 = ~n1741;
  assign n1729 = n1742 & n1743;
  assign n1745 = n1753 & n1754;
  assign n78317 = n1755 ^ n804;
  assign n827 = ~n804;
  assign n1768 = n1776 & n1777;
  assign n1704 = n1655 & n298;
  assign n1694 = n1718 ^ n1719;
  assign n1702 = ~n1655;
  assign n1720 = ~n1718;
  assign n1689 = ~n1729;
  assign n1727 = ~n1745;
  assign n1715 = n827 & n1755;
  assign n1730 = n827 & n1756;
  assign n1757 = ~n1768;
  assign n1675 = n299 ^ n1694;
  assign n1699 = n1702 & n1703;
  assign n1657 = ~n1704;
  assign n1705 = n1720 & n1721;
  assign n1706 = n1727 & n1728;
  assign n1644 = n1730 ^ n1731;
  assign n1712 = ~n1715;
  assign n1733 = n1757 & n1758;
  assign n1660 = n1674 ^ n1675;
  assign n1676 = ~n1675;
  assign n1680 = ~n1699;
  assign n1695 = ~n1705;
  assign n1686 = n1706 ^ n1707;
  assign n1710 = n1644 & n1722;
  assign n1709 = ~n1706;
  assign n1711 = ~n1644;
  assign n774 = n1732 ^ n1733;
  assign n1734 = ~n1733;
  assign n1653 = n1660 & n78315;
  assign n1651 = ~n1660;
  assign n1631 = n1676 & n1677;
  assign n1604 = n1686 ^ n1687;
  assign n1679 = n1695 & n1696;
  assign n1700 = n1708 & n1709;
  assign n1646 = ~n1710;
  assign n1701 = n1711 & n1667;
  assign n78332 = n1715 ^ n774;
  assign n1697 = n774 & n1723;
  assign n778 = ~n774;
  assign n1724 = n1734 & n1735;
  assign n1642 = n1651 & n1652;
  assign n1630 = ~n1653;
  assign n1634 = ~n1631;
  assign n1663 = n1604 & n1678;
  assign n1654 = n298 ^ n1679;
  assign n1664 = ~n1604;
  assign n1681 = ~n1679;
  assign n1622 = n1697 ^ n1698;
  assign n1688 = ~n1700;
  assign n1669 = ~n1701;
  assign n1650 = n778 & n1712;
  assign n1713 = ~n1724;
  assign n1629 = n1630 & n1587;
  assign n1612 = ~n1642;
  assign n1632 = n1654 ^ n1655;
  assign n1637 = ~n1663;
  assign n1661 = n1664 & n297;
  assign n1665 = n1680 & n1681;
  assign n1682 = n1622 & n1684;
  assign n1666 = n1688 & n1689;
  assign n1683 = ~n1622;
  assign n1658 = ~n1650;
  assign n1690 = n1713 & n1714;
  assign n1611 = ~n1629;
  assign n1616 = n1612 & n1630;
  assign n1554 = n1631 ^ n1632;
  assign n1633 = ~n1632;
  assign n1606 = ~n1661;
  assign n1656 = ~n1665;
  assign n1643 = n1666 ^ n1667;
  assign n1624 = ~n1682;
  assign n1670 = n1683 & n1591;
  assign n1668 = ~n1666;
  assign n1671 = n1690 ^ n1691;
  assign n1692 = ~n1690;
  assign n1584 = n1611 & n1612;
  assign n1601 = n1554 & n1613;
  assign n1588 = ~n1616;
  assign n1602 = ~n1554;
  assign n1575 = n1633 & n1634;
  assign n1635 = n1643 ^ n1644;
  assign n1636 = n1656 & n1657;
  assign n1662 = n1668 & n1669;
  assign n1593 = ~n1670;
  assign n735 = n1671 ^ n1640;
  assign n1685 = n1692 & n1693;
  assign n1553 = n1584 ^ n1585;
  assign n1569 = n1587 ^ n1588;
  assign n1573 = ~n1584;
  assign n1546 = ~n1601;
  assign n1589 = n1602 & n1585;
  assign n1578 = ~n1575;
  assign n1619 = n1635 & n296;
  assign n1603 = n297 ^ n1636;
  assign n1617 = ~n1635;
  assign n1638 = ~n1636;
  assign n78331 = n1650 ^ n735;
  assign n1600 = n735 & n1658;
  assign n1639 = n735 & n1659;
  assign n1645 = ~n1662;
  assign n739 = ~n735;
  assign n1672 = ~n1685;
  assign n1526 = n1553 ^ n1554;
  assign n78283 = n1569 ^ n78284;
  assign n1571 = ~n1569;
  assign n1574 = ~n1589;
  assign n1576 = n1603 ^ n1604;
  assign n1614 = n1617 & n1618;
  assign n1540 = ~n1619;
  assign n1620 = n1637 & n1638;
  assign n1563 = n1639 ^ n1640;
  assign n1621 = n1645 & n1646;
  assign n1595 = ~n1600;
  assign n1647 = n1672 & n1673;
  assign n1525 = n1571 & n1572;
  assign n1555 = n1573 & n1574;
  assign n1517 = n1575 ^ n1576;
  assign n1577 = ~n1576;
  assign n1580 = ~n1614;
  assign n1609 = n1563 & n1528;
  assign n1605 = ~n1620;
  assign n1590 = n1621 ^ n1622;
  assign n1607 = ~n1563;
  assign n1623 = ~n1621;
  assign n1626 = n1647 ^ n1582;
  assign n1648 = ~n1647;
  assign n78282 = n1525 ^ n1526;
  assign n1453 = n1526 & n1525;
  assign n1547 = n1517 & n1487;
  assign n1545 = ~n1555;
  assign n1548 = ~n1517;
  assign n1537 = n1577 & n1578;
  assign n1556 = n1580 & n1540;
  assign n1509 = n1590 ^ n1591;
  assign n1557 = n1605 & n1606;
  assign n1594 = n1607 & n1608;
  assign n1530 = ~n1609;
  assign n1615 = n1623 & n1624;
  assign n673 = n1625 ^ n1626;
  assign n1641 = n1648 & n1649;
  assign n1473 = ~n1453;
  assign n1516 = n1545 & n1546;
  assign n1519 = ~n1547;
  assign n1536 = n1548 & n1549;
  assign n1538 = n1556 ^ n1557;
  assign n1560 = n1509 & n311;
  assign n1558 = ~n1509;
  assign n1579 = ~n1557;
  assign n1565 = ~n1594;
  assign n78330 = n1600 ^ n673;
  assign n1581 = n673 & n1610;
  assign n1592 = ~n1615;
  assign n703 = ~n673;
  assign n1627 = ~n1641;
  assign n1486 = n1516 ^ n1517;
  assign n1518 = ~n1516;
  assign n1489 = ~n1536;
  assign n1520 = n1537 ^ n1538;
  assign n1462 = n1538 & n1537;
  assign n1550 = n1558 & n1559;
  assign n1483 = ~n1560;
  assign n1561 = n1579 & n1580;
  assign n1481 = n1581 ^ n1582;
  assign n1562 = n1592 & n1593;
  assign n1570 = n703 & n1595;
  assign n1597 = n1627 & n1628;
  assign n1454 = n1486 ^ n1487;
  assign n1505 = n1518 & n1519;
  assign n1506 = n1520 & n1521;
  assign n1459 = ~n1520;
  assign n1465 = ~n1462;
  assign n1510 = ~n1550;
  assign n1542 = n1481 & n1551;
  assign n1539 = ~n1561;
  assign n1527 = n1562 ^ n1563;
  assign n1541 = ~n1481;
  assign n1564 = ~n1562;
  assign n1566 = ~n1570;
  assign n678 = n1596 ^ n1597;
  assign n1598 = ~n1597;
  assign n78281 = n1453 ^ n1454;
  assign n1396 = n1454 & n1473;
  assign n1488 = ~n1505;
  assign n1460 = ~n1506;
  assign n1494 = n1459 & n1428;
  assign n1467 = n1527 ^ n1528;
  assign n1508 = n1539 & n1540;
  assign n1531 = n1541 & n1499;
  assign n1475 = ~n1542;
  assign n1552 = n1564 & n1565;
  assign n1493 = n678 & n1566;
  assign n78329 = n1570 ^ n678;
  assign n1543 = n678 & n1583;
  assign n682 = ~n678;
  assign n1586 = n1598 & n1599;
  assign n1399 = ~n1396;
  assign n1458 = n1488 & n1489;
  assign n1430 = ~n1494;
  assign n1495 = n1467 & n1507;
  assign n1490 = n1508 ^ n1509;
  assign n1496 = ~n1467;
  assign n1511 = ~n1508;
  assign n1501 = ~n1531;
  assign n1522 = n1543 ^ n1544;
  assign n1529 = ~n1552;
  assign n1567 = ~n1586;
  assign n1427 = n1458 ^ n1459;
  assign n1461 = ~n1458;
  assign n1463 = n311 ^ n1490;
  assign n1469 = ~n1495;
  assign n1491 = n1496 & n310;
  assign n1497 = n1510 & n1511;
  assign n1514 = n1522 & n1523;
  assign n1498 = n1529 & n1530;
  assign n1512 = ~n1522;
  assign n1533 = n1567 & n1568;
  assign n1397 = n1427 ^ n1428;
  assign n1448 = n1460 & n1461;
  assign n1363 = n1462 ^ n1463;
  assign n1464 = ~n1463;
  assign n1435 = ~n1491;
  assign n1482 = ~n1497;
  assign n1480 = n1498 ^ n1499;
  assign n1502 = n1512 & n1513;
  assign n1426 = ~n1514;
  assign n1500 = ~n1498;
  assign n647 = n1532 ^ n1533;
  assign n1534 = ~n1533;
  assign n78280 = n1396 ^ n1397;
  assign n1398 = ~n1397;
  assign n1432 = n1363 & n1437;
  assign n1429 = ~n1448;
  assign n1431 = ~n1363;
  assign n1404 = n1464 & n1465;
  assign n1409 = n1480 ^ n1481;
  assign n1466 = n1482 & n1483;
  assign n1492 = n1500 & n1501;
  assign n1442 = ~n1502;
  assign n1484 = n647 & n1515;
  assign n1416 = n647 & n1493;
  assign n666 = ~n647;
  assign n1524 = n1534 & n1535;
  assign n1335 = n1398 & n1399;
  assign n1400 = n1429 & n1430;
  assign n1421 = n1431 & n1401;
  assign n1366 = ~n1432;
  assign n1407 = ~n1404;
  assign n1451 = n1409 & n309;
  assign n1433 = n1466 ^ n1467;
  assign n1449 = ~n1409;
  assign n1468 = ~n1466;
  assign n1476 = n1442 & n1426;
  assign n1470 = n1484 ^ n1485;
  assign n1474 = ~n1492;
  assign n78328 = n1493 ^ n666;
  assign n1503 = ~n1524;
  assign n1364 = n1400 ^ n1401;
  assign n1402 = ~n1400;
  assign n1403 = ~n1421;
  assign n1405 = n310 ^ n1433;
  assign n1438 = n1449 & n1450;
  assign n1372 = ~n1451;
  assign n1452 = n1468 & n1469;
  assign n1457 = n1470 & n1471;
  assign n1439 = n1474 & n1475;
  assign n1440 = ~n1476;
  assign n1455 = ~n1470;
  assign n1477 = n1503 & n1504;
  assign n1336 = n1363 ^ n1364;
  assign n1386 = n1402 & n1403;
  assign n1377 = n1404 ^ n1405;
  assign n1406 = ~n1405;
  assign n1411 = ~n1438;
  assign n1342 = n1439 ^ n1440;
  assign n1434 = ~n1452;
  assign n1443 = n1455 & n1456;
  assign n1359 = ~n1457;
  assign n1441 = ~n1439;
  assign n1445 = n1477 ^ n1393;
  assign n1478 = ~n1477;
  assign n78279 = n1335 ^ n1336;
  assign n1263 = n1336 & n1335;
  assign n1369 = n1377 & n1378;
  assign n1365 = ~n1386;
  assign n1367 = ~n1377;
  assign n1339 = n1406 & n1407;
  assign n1408 = n1434 & n1435;
  assign n1424 = n1342 & n308;
  assign n1422 = ~n1342;
  assign n1436 = n1441 & n1442;
  assign n1391 = ~n1443;
  assign n641 = n1444 ^ n1445;
  assign n1472 = n1478 & n1479;
  assign n1297 = n1365 & n1366;
  assign n1354 = n1367 & n1368;
  assign n1338 = ~n1369;
  assign n1370 = n1408 ^ n1409;
  assign n78327 = n1416 ^ n641;
  assign n1410 = ~n1408;
  assign n1413 = n1422 & n1423;
  assign n1318 = ~n1424;
  assign n1414 = n1391 & n1359;
  assign n1425 = ~n1436;
  assign n643 = ~n641;
  assign n1446 = ~n1472;
  assign n1337 = ~n1297;
  assign n1312 = ~n1354;
  assign n1340 = n309 ^ n1370;
  assign n1387 = n1410 & n1411;
  assign n1344 = ~n1413;
  assign n1389 = ~n1414;
  assign n1392 = n643 & n1415;
  assign n1385 = n643 & n1416;
  assign n1388 = n1425 & n1426;
  assign n1418 = n1446 & n1447;
  assign n1323 = n1337 & n1338;
  assign n1324 = n1338 & n1312;
  assign n1279 = n1339 ^ n1340;
  assign n1282 = n1340 & n1339;
  assign n1371 = ~n1387;
  assign n1373 = n1388 ^ n1389;
  assign n1302 = n1392 ^ n1393;
  assign n1394 = ~n1385;
  assign n1390 = ~n1388;
  assign n623 = n1417 ^ n1418;
  assign n1419 = ~n1418;
  assign n1315 = n1279 & n1241;
  assign n1311 = ~n1323;
  assign n1298 = ~n1324;
  assign n1313 = ~n1279;
  assign n1285 = ~n1282;
  assign n1341 = n1371 & n1372;
  assign n1357 = n1373 & n307;
  assign n1360 = n1302 & n1327;
  assign n1355 = ~n1373;
  assign n1361 = ~n1302;
  assign n78326 = n1385 ^ n623;
  assign n1379 = n1390 & n1391;
  assign n1374 = n623 & n1395;
  assign n1382 = n623 & n616;
  assign n1380 = ~n623;
  assign n1412 = n1419 & n1420;
  assign n1264 = n1297 ^ n1298;
  assign n1278 = n1311 & n1312;
  assign n1300 = n1313 & n1314;
  assign n1280 = ~n1315;
  assign n1316 = n1341 ^ n1342;
  assign n1343 = ~n1341;
  assign n1348 = n1355 & n1356;
  assign n1251 = ~n1357;
  assign n1304 = ~n1360;
  assign n1350 = n1361 & n1362;
  assign n1232 = n1374 ^ n1375;
  assign n1358 = ~n1379;
  assign n1376 = n1380 & n1381;
  assign n625 = ~n1382;
  assign n1299 = n1380 & n1394;
  assign n1383 = ~n1412;
  assign n78278 = n1263 ^ n1264;
  assign n1220 = n1264 & n1263;
  assign n1240 = n1278 ^ n1279;
  assign n1281 = ~n1278;
  assign n1243 = ~n1300;
  assign n1283 = n308 ^ n1316;
  assign n1325 = n1343 & n1344;
  assign n1290 = ~n1348;
  assign n1345 = n1232 & n1349;
  assign n1329 = ~n1350;
  assign n1326 = n1358 & n1359;
  assign n1346 = ~n1232;
  assign n618 = ~n1376;
  assign n1319 = ~n1299;
  assign n1351 = n1383 & n1384;
  assign n1221 = n1240 ^ n1241;
  assign n1225 = ~n1220;
  assign n1262 = n1280 & n1281;
  assign n1257 = n1282 ^ n1283;
  assign n1284 = ~n1283;
  assign n1317 = ~n1325;
  assign n1287 = n1290 & n1251;
  assign n1301 = n1326 ^ n1327;
  assign n1234 = ~n1345;
  assign n1330 = n1346 & n1270;
  assign n1328 = ~n1326;
  assign n1332 = n1351 ^ n1292;
  assign n1352 = ~n1351;
  assign n78277 = n1220 ^ n1221;
  assign n1147 = n1221 & n1225;
  assign n1244 = n1257 & n1258;
  assign n1242 = ~n1262;
  assign n1245 = ~n1257;
  assign n1247 = n1284 & n1285;
  assign n1217 = n1301 ^ n1302;
  assign n1288 = n1317 & n1318;
  assign n1322 = n1328 & n1329;
  assign n1272 = ~n1330;
  assign n611 = n1331 ^ n1332;
  assign n1347 = n1352 & n1353;
  assign n1174 = n1242 & n1243;
  assign n1190 = ~n1244;
  assign n1230 = n1245 & n1246;
  assign n1266 = n1217 & n1286;
  assign n1248 = n1287 ^ n1288;
  assign n1267 = ~n1217;
  assign n78325 = n1299 ^ n611;
  assign n1289 = ~n1288;
  assign n1265 = n611 & n1319;
  assign n1291 = n611 & n1320;
  assign n1305 = n611 & n1321;
  assign n1303 = ~n1322;
  assign n1306 = ~n611;
  assign n1333 = ~n1347;
  assign n1212 = ~n1174;
  assign n1213 = ~n1230;
  assign n1163 = n1247 ^ n1248;
  assign n1219 = ~n1266;
  assign n1259 = n1267 & n306;
  assign n1249 = ~n1248;
  assign n1268 = n1289 & n1290;
  assign n1177 = n1291 ^ n1292;
  assign n1269 = n1303 & n1304;
  assign n1274 = ~n1265;
  assign n613 = ~n1305;
  assign n1295 = n1306 & n603;
  assign n1308 = n1333 & n1334;
  assign n1197 = n1212 & n1213;
  assign n1198 = n1213 & n1190;
  assign n1215 = n1163 & n1226;
  assign n1214 = ~n1163;
  assign n1166 = n1249 & n1247;
  assign n1193 = ~n1259;
  assign n1252 = n1177 & n1205;
  assign n1250 = ~n1268;
  assign n1231 = n1269 ^ n1270;
  assign n1253 = ~n1177;
  assign n1271 = ~n1269;
  assign n606 = ~n1295;
  assign n599 = n1307 ^ n1308;
  assign n1309 = ~n1308;
  assign n1189 = ~n1197;
  assign n1175 = ~n1198;
  assign n1199 = n1214 & n1143;
  assign n1165 = ~n1215;
  assign n1137 = n1231 ^ n1232;
  assign n1216 = n1250 & n1251;
  assign n1179 = ~n1252;
  assign n1235 = n1253 & n1254;
  assign n78340 = n1265 ^ n599;
  assign n1260 = n1271 & n1272;
  assign n1255 = n599 & n1293;
  assign n1275 = n599 & n1294;
  assign n1273 = ~n599;
  assign n1296 = n1309 & n1310;
  assign n1158 = n1174 ^ n1175;
  assign n1162 = n1189 & n1190;
  assign n1132 = ~n1199;
  assign n1202 = n1137 & n305;
  assign n1191 = n1216 ^ n1217;
  assign n1200 = ~n1137;
  assign n1218 = ~n1216;
  assign n1207 = ~n1235;
  assign n1227 = n1255 ^ n1256;
  assign n1233 = ~n1260;
  assign n1180 = n1273 & n1274;
  assign n1261 = n1273 & n591;
  assign n601 = ~n1275;
  assign n1276 = ~n1296;
  assign n78292 = n1147 ^ n1158;
  assign n1142 = n1162 ^ n1163;
  assign n1146 = ~n1158;
  assign n1164 = ~n1162;
  assign n1167 = n306 ^ n1191;
  assign n1195 = n1200 & n1201;
  assign n1139 = ~n1202;
  assign n1203 = n1218 & n1219;
  assign n1224 = n1227 & n1228;
  assign n1204 = n1233 & n1234;
  assign n1222 = ~n1227;
  assign n594 = ~n1261;
  assign n1236 = n1276 & n1277;
  assign n1106 = n1142 ^ n1143;
  assign n1105 = n1146 & n1147;
  assign n1148 = n1164 & n1165;
  assign n1079 = n1166 ^ n1167;
  assign n1098 = n1167 & n1166;
  assign n1171 = ~n1195;
  assign n1192 = ~n1203;
  assign n1176 = n1204 ^ n1205;
  assign n1208 = n1222 & n1223;
  assign n1121 = ~n1224;
  assign n1206 = ~n1204;
  assign n1209 = n1236 ^ n1237;
  assign n1238 = ~n1236;
  assign n78291 = n1105 ^ n1106;
  assign n1107 = ~n1106;
  assign n1135 = n1079 & n1109;
  assign n1131 = ~n1148;
  assign n1133 = ~n1079;
  assign n1102 = n1176 ^ n1177;
  assign n1169 = n1192 & n1193;
  assign n1196 = n1206 & n1207;
  assign n1155 = ~n1208;
  assign n582 = n1209 ^ n1157;
  assign n1229 = n1238 & n1239;
  assign n1043 = n1107 & n1105;
  assign n1108 = n1131 & n1132;
  assign n1116 = n1133 & n1134;
  assign n1081 = ~n1135;
  assign n1149 = n1102 & n1168;
  assign n1136 = n305 ^ n1169;
  assign n1150 = ~n1102;
  assign n1170 = ~n1169;
  assign n78339 = n1180 ^ n582;
  assign n1181 = n1155 & n1121;
  assign n1184 = n582 & n1194;
  assign n1127 = n582 & n1180;
  assign n1178 = ~n1196;
  assign n1182 = ~n582;
  assign n1210 = ~n1229;
  assign n1046 = ~n1043;
  assign n1078 = n1108 ^ n1109;
  assign n1110 = ~n1108;
  assign n1111 = ~n1116;
  assign n1099 = n1136 ^ n1137;
  assign n1104 = ~n1149;
  assign n1144 = n1150 & n304;
  assign n1151 = n1170 & n1171;
  assign n1152 = n1178 & n1179;
  assign n1153 = ~n1181;
  assign n1156 = n1182 & n1183;
  assign n580 = ~n1184;
  assign n1172 = n1182 & n587;
  assign n1185 = n1210 & n1211;
  assign n1044 = n1078 ^ n1079;
  assign n1048 = n1098 ^ n1099;
  assign n1097 = n1110 & n1111;
  assign n1100 = ~n1099;
  assign n1073 = ~n1144;
  assign n1138 = ~n1151;
  assign n1038 = n1152 ^ n1153;
  assign n1059 = n1156 ^ n1157;
  assign n1154 = ~n1152;
  assign n589 = ~n1172;
  assign n1159 = n1185 ^ n1186;
  assign n1187 = ~n1185;
  assign n78290 = n1043 ^ n1044;
  assign n1045 = ~n1044;
  assign n1084 = n1048 & n1012;
  assign n1082 = ~n1048;
  assign n1080 = ~n1097;
  assign n1051 = n1100 & n1098;
  assign n1101 = n1138 & n1139;
  assign n1119 = n1038 & n319;
  assign n1122 = n1059 & n1140;
  assign n1117 = ~n1038;
  assign n1123 = ~n1059;
  assign n1145 = n1154 & n1155;
  assign n568 = n1159 ^ n1092;
  assign n1173 = n1187 & n1188;
  assign n989 = n1045 & n1046;
  assign n1047 = n1080 & n1081;
  assign n1070 = n1082 & n1083;
  assign n1050 = ~n1084;
  assign n1054 = ~n1051;
  assign n1071 = n1101 ^ n1102;
  assign n1103 = ~n1101;
  assign n1112 = n1117 & n1118;
  assign n1018 = ~n1119;
  assign n1061 = ~n1122;
  assign n1113 = n1123 & n1088;
  assign n78338 = n1127 ^ n568;
  assign n1069 = n568 & n1127;
  assign n1126 = n568 & n1141;
  assign n1120 = ~n1145;
  assign n1124 = ~n568;
  assign n1160 = ~n1173;
  assign n995 = ~n989;
  assign n1011 = n1047 ^ n1048;
  assign n1049 = ~n1047;
  assign n1014 = ~n1070;
  assign n1052 = n304 ^ n1071;
  assign n1086 = n1103 & n1104;
  assign n1040 = ~n1112;
  assign n1090 = ~n1113;
  assign n1087 = n1120 & n1121;
  assign n1091 = n1124 & n1125;
  assign n1075 = ~n1069;
  assign n1114 = n1124 & n578;
  assign n570 = ~n1126;
  assign n1128 = n1160 & n1161;
  assign n990 = n1011 ^ n1012;
  assign n1036 = n1049 & n1050;
  assign n1022 = n1051 ^ n1052;
  assign n1053 = ~n1052;
  assign n1072 = ~n1086;
  assign n1058 = n1087 ^ n1088;
  assign n1007 = n1091 ^ n1092;
  assign n1089 = ~n1087;
  assign n573 = ~n1114;
  assign n1094 = n1128 ^ n1042;
  assign n1129 = ~n1128;
  assign n78289 = n989 ^ n990;
  assign n921 = n990 & n995;
  assign n1015 = n1022 & n1023;
  assign n1013 = ~n1036;
  assign n942 = ~n1022;
  assign n983 = n1053 & n1054;
  assign n986 = n1058 ^ n1059;
  assign n1037 = n1072 & n1073;
  assign n1062 = n1007 & n1074;
  assign n1063 = ~n1007;
  assign n1085 = n1089 & n1090;
  assign n564 = n1093 ^ n1094;
  assign n1115 = n1129 & n1130;
  assign n914 = ~n921;
  assign n979 = n1013 & n1014;
  assign n1005 = n942 & n980;
  assign n982 = ~n1015;
  assign n1026 = n986 & n318;
  assign n1016 = n1037 ^ n1038;
  assign n1024 = ~n986;
  assign n1039 = ~n1037;
  assign n997 = ~n1062;
  assign n1055 = n1063 & n1029;
  assign n78337 = n1069 ^ n564;
  assign n991 = n564 & n1075;
  assign n1041 = n564 & n1076;
  assign n1064 = n564 & n1077;
  assign n1060 = ~n1085;
  assign n1065 = ~n564;
  assign n1095 = ~n1115;
  assign n943 = n979 ^ n980;
  assign n981 = ~n979;
  assign n945 = ~n1005;
  assign n984 = n319 ^ n1016;
  assign n1019 = n1024 & n1025;
  assign n949 = ~n1026;
  assign n1027 = n1039 & n1040;
  assign n936 = n1041 ^ n1042;
  assign n1031 = ~n1055;
  assign n1028 = n1060 & n1061;
  assign n566 = ~n1064;
  assign n1056 = n1065 & n555;
  assign n1066 = n1095 & n1096;
  assign n922 = n942 ^ n943;
  assign n968 = n981 & n982;
  assign n954 = n983 ^ n984;
  assign n919 = n984 & n983;
  assign n988 = ~n1019;
  assign n1008 = n936 & n1020;
  assign n1017 = ~n1027;
  assign n1006 = n1028 ^ n1029;
  assign n1009 = ~n936;
  assign n1030 = ~n1028;
  assign n558 = ~n1056;
  assign n1033 = n1066 ^ n976;
  assign n1067 = ~n1066;
  assign n78288 = n921 ^ n922;
  assign n913 = ~n922;
  assign n946 = n954 & n955;
  assign n944 = ~n968;
  assign n916 = ~n954;
  assign n889 = n1006 ^ n1007;
  assign n938 = ~n1008;
  assign n998 = n1009 & n974;
  assign n985 = n1017 & n1018;
  assign n1021 = n1030 & n1031;
  assign n549 = n1032 ^ n1033;
  assign n1057 = n1067 & n1068;
  assign n862 = n913 & n914;
  assign n915 = n944 & n945;
  assign n918 = ~n946;
  assign n934 = n916 & n882;
  assign n971 = n889 & n317;
  assign n947 = n985 ^ n986;
  assign n969 = ~n889;
  assign n959 = ~n998;
  assign n987 = ~n985;
  assign n975 = n549 & n1010;
  assign n1000 = n549 & n546;
  assign n966 = n549 & n991;
  assign n996 = ~n1021;
  assign n992 = ~n549;
  assign n1034 = ~n1057;
  assign n865 = ~n862;
  assign n881 = n915 ^ n916;
  assign n917 = ~n915;
  assign n884 = ~n934;
  assign n920 = n318 ^ n947;
  assign n956 = n969 & n970;
  assign n891 = ~n971;
  assign n873 = n975 ^ n976;
  assign n972 = n987 & n988;
  assign n78336 = n991 ^ n992;
  assign n973 = n996 & n997;
  assign n993 = n992 & n999;
  assign n551 = ~n1000;
  assign n961 = ~n966;
  assign n1002 = n1034 & n1035;
  assign n863 = n881 ^ n882;
  assign n899 = n917 & n918;
  assign n834 = n919 ^ n920;
  assign n855 = n920 & n919;
  assign n925 = ~n956;
  assign n950 = n873 & n957;
  assign n951 = ~n873;
  assign n948 = ~n972;
  assign n935 = n973 ^ n974;
  assign n958 = ~n973;
  assign n544 = ~n993;
  assign n967 = n1001 ^ n1002;
  assign n1003 = ~n1002;
  assign n78287 = n862 ^ n863;
  assign n797 = n863 & n865;
  assign n887 = n834 & n852;
  assign n883 = ~n899;
  assign n885 = ~n834;
  assign n858 = ~n855;
  assign n829 = n935 ^ n936;
  assign n923 = n948 & n949;
  assign n875 = ~n950;
  assign n939 = n951 & n905;
  assign n952 = n958 & n959;
  assign n78335 = n966 ^ n967;
  assign n940 = n967 & n977;
  assign n963 = n967 & n978;
  assign n960 = ~n967;
  assign n994 = n1003 & n1004;
  assign n802 = ~n797;
  assign n851 = n883 & n884;
  assign n870 = n885 & n886;
  assign n853 = ~n887;
  assign n902 = n829 & n316;
  assign n888 = n317 ^ n923;
  assign n900 = ~n829;
  assign n924 = ~n923;
  assign n907 = ~n939;
  assign n812 = n940 ^ n941;
  assign n937 = ~n952;
  assign n871 = n960 & n961;
  assign n953 = n960 & n962;
  assign n542 = ~n963;
  assign n964 = ~n994;
  assign n835 = n851 ^ n852;
  assign n854 = ~n851;
  assign n824 = ~n870;
  assign n856 = n888 ^ n889;
  assign n894 = n900 & n901;
  assign n831 = ~n902;
  assign n903 = n924 & n925;
  assign n928 = n812 & n844;
  assign n926 = ~n812;
  assign n904 = n937 & n938;
  assign n530 = ~n953;
  assign n930 = n964 & n965;
  assign n798 = n834 ^ n835;
  assign n838 = n853 & n854;
  assign n768 = n855 ^ n856;
  assign n857 = ~n856;
  assign n860 = ~n894;
  assign n890 = ~n903;
  assign n872 = n904 ^ n905;
  assign n908 = n926 & n927;
  assign n814 = ~n928;
  assign n906 = ~n904;
  assign n539 = n542 & n530;
  assign n910 = n930 ^ n931;
  assign n933 = n930 & n897;
  assign n932 = ~n930;
  assign n78286 = n797 ^ n798;
  assign n801 = ~n798;
  assign n825 = n768 & n804;
  assign n823 = ~n838;
  assign n826 = ~n768;
  assign n779 = n857 & n858;
  assign n794 = n872 ^ n873;
  assign n859 = n890 & n891;
  assign n895 = n906 & n907;
  assign n846 = ~n908;
  assign n528 = n909 ^ n910;
  assign n929 = n932 & n912;
  assign n911 = ~n933;
  assign n751 = n801 & n802;
  assign n803 = n823 & n824;
  assign n771 = ~n825;
  assign n810 = n826 & n827;
  assign n807 = ~n779;
  assign n841 = n794 & n315;
  assign n828 = n316 ^ n859;
  assign n839 = ~n794;
  assign n78334 = n871 ^ n528;
  assign n861 = ~n859;
  assign n878 = n528 & n892;
  assign n818 = n528 & n871;
  assign n874 = ~n895;
  assign n876 = ~n528;
  assign n898 = n911 & n912;
  assign n896 = ~n929;
  assign n759 = ~n751;
  assign n769 = n803 ^ n804;
  assign n805 = ~n803;
  assign n806 = ~n810;
  assign n791 = n828 ^ n829;
  assign n836 = n839 & n840;
  assign n767 = ~n841;
  assign n842 = n860 & n861;
  assign n843 = n874 & n875;
  assign n847 = n876 & n877;
  assign n521 = ~n878;
  assign n866 = n876 & n522;
  assign n893 = n896 & n897;
  assign n879 = ~n898;
  assign n752 = n768 ^ n769;
  assign n777 = n779 ^ n791;
  assign n790 = n805 & n806;
  assign n755 = n791 & n807;
  assign n780 = ~n791;
  assign n796 = ~n836;
  assign n830 = ~n842;
  assign n811 = n843 ^ n844;
  assign n761 = n847 ^ n848;
  assign n845 = ~n843;
  assign n526 = ~n866;
  assign n869 = n879 & n880;
  assign n867 = ~n893;
  assign n78285 = n751 ^ n752;
  assign n708 = n752 & n759;
  assign n772 = n777 & n778;
  assign n773 = n779 ^ n780;
  assign n770 = ~n790;
  assign n758 = ~n755;
  assign n748 = n811 ^ n812;
  assign n793 = n830 & n831;
  assign n815 = n761 & n785;
  assign n816 = ~n761;
  assign n837 = n845 & n846;
  assign n864 = n867 & n868;
  assign n850 = ~n869;
  assign n730 = n770 & n771;
  assign n732 = ~n772;
  assign n764 = n773 & n774;
  assign n781 = n748 & n792;
  assign n765 = n793 ^ n794;
  assign n782 = ~n748;
  assign n795 = ~n793;
  assign n763 = ~n815;
  assign n808 = n816 & n817;
  assign n813 = ~n837;
  assign n849 = ~n864;
  assign n754 = ~n730;
  assign n753 = ~n764;
  assign n756 = n315 ^ n765;
  assign n750 = ~n781;
  assign n775 = n782 & n314;
  assign n783 = n795 & n796;
  assign n787 = ~n808;
  assign n784 = n813 & n814;
  assign n819 = n849 & n850;
  assign n745 = n753 & n754;
  assign n729 = n753 & n732;
  assign n738 = n755 ^ n756;
  assign n757 = ~n756;
  assign n728 = ~n775;
  assign n766 = ~n783;
  assign n760 = n784 ^ n785;
  assign n786 = ~n784;
  assign n78333 = n818 ^ n819;
  assign n799 = n819 & n832;
  assign n822 = n819 & n833;
  assign n820 = ~n819;
  assign n723 = n729 ^ n730;
  assign n733 = n738 & n739;
  assign n731 = ~n745;
  assign n734 = ~n738;
  assign n715 = n757 & n758;
  assign n720 = n760 ^ n761;
  assign n747 = n766 & n767;
  assign n776 = n786 & n787;
  assign n744 = n799 ^ n800;
  assign n809 = n820 & n821;
  assign n789 = ~n822;
  assign n693 = n723 & n708;
  assign n709 = ~n723;
  assign n699 = n731 & n732;
  assign n701 = ~n733;
  assign n724 = n734 & n735;
  assign n718 = ~n715;
  assign n740 = n720 & n746;
  assign n736 = n747 ^ n748;
  assign n741 = ~n720;
  assign n749 = ~n747;
  assign n762 = ~n776;
  assign n788 = ~n809;
  assign n78300 = n708 ^ n709;
  assign n684 = ~n693;
  assign n713 = ~n699;
  assign n714 = ~n724;
  assign n716 = n314 ^ n736;
  assign n722 = ~n740;
  assign n737 = n741 & n313;
  assign n742 = n749 & n750;
  assign n743 = n762 & n763;
  assign n514 = n788 & n789;
  assign n710 = n713 & n714;
  assign n698 = n714 & n701;
  assign n687 = n715 ^ n716;
  assign n717 = ~n716;
  assign n707 = ~n737;
  assign n727 = ~n742;
  assign n725 = n743 ^ n744;
  assign n694 = n698 ^ n699;
  assign n704 = n687 & n673;
  assign n700 = ~n710;
  assign n702 = ~n687;
  assign n690 = n717 & n718;
  assign n711 = n725 ^ n726;
  assign n719 = n727 & n728;
  assign n78299 = n693 ^ n694;
  assign n685 = ~n694;
  assign n686 = n700 & n701;
  assign n697 = n702 & n703;
  assign n689 = ~n704;
  assign n696 = n312 ^ n711;
  assign n705 = n719 ^ n720;
  assign n721 = ~n719;
  assign n668 = n684 & n685;
  assign n672 = n686 ^ n687;
  assign n688 = ~n686;
  assign n675 = ~n697;
  assign n691 = n313 ^ n705;
  assign n712 = n721 & n722;
  assign n669 = n672 ^ n673;
  assign n670 = ~n668;
  assign n683 = n688 & n689;
  assign n681 = n690 ^ n691;
  assign n692 = ~n691;
  assign n706 = ~n712;
  assign n78298 = n668 ^ n669;
  assign n649 = n669 & n670;
  assign n676 = n681 & n682;
  assign n674 = ~n683;
  assign n677 = ~n681;
  assign n679 = n692 & n690;
  assign n695 = n706 & n707;
  assign n656 = n674 & n675;
  assign n659 = ~n676;
  assign n671 = n677 & n678;
  assign n680 = n695 ^ n696;
  assign n663 = ~n656;
  assign n664 = ~n671;
  assign n653 = n679 ^ n680;
  assign n660 = n663 & n664;
  assign n662 = n664 & n659;
  assign n667 = n653 & n647;
  assign n665 = ~n653;
  assign n658 = ~n660;
  assign n657 = ~n662;
  assign n661 = n665 & n666;
  assign n655 = ~n667;
  assign n651 = n656 ^ n657;
  assign n652 = n658 & n659;
  assign n645 = ~n661;
  assign n78297 = n649 ^ n651;
  assign n646 = n652 ^ n653;
  assign n648 = ~n651;
  assign n654 = ~n652;
  assign n637 = n646 ^ n647;
  assign n636 = n648 & n649;
  assign n650 = n654 & n655;
  assign n78296 = n636 ^ n637;
  assign n638 = ~n637;
  assign n639 = ~n636;
  assign n644 = ~n650;
  assign n619 = n638 & n639;
  assign n642 = n644 & n645;
  assign n635 = n642 & n643;
  assign n640 = ~n642;
  assign n632 = ~n635;
  assign n634 = n640 & n641;
  assign n631 = n632 & n633;
  assign n629 = ~n634;
  assign n628 = ~n631;
  assign n630 = n629 & n632;
  assign n622 = n628 & n629;
  assign n626 = ~n630;
  assign n615 = n622 ^ n623;
  assign n620 = n626 ^ n627;
  assign n624 = ~n622;
  assign n609 = n615 ^ n616;
  assign n78295 = n619 ^ n620;
  assign n608 = n620 & n619;
  assign n621 = n624 & n625;
  assign n78294 = n608 ^ n609;
  assign n614 = ~n608;
  assign n617 = ~n621;
  assign n597 = n609 & n614;
  assign n610 = n617 & n618;
  assign n604 = n610 ^ n611;
  assign n612 = ~n610;
  assign n602 = n603 ^ n604;
  assign n607 = n612 & n613;
  assign n78293 = n597 ^ n602;
  assign n596 = ~n602;
  assign n605 = ~n607;
  assign n585 = n596 & n597;
  assign n598 = n605 & n606;
  assign n592 = n598 ^ n599;
  assign n600 = ~n598;
  assign n590 = n591 ^ n592;
  assign n595 = n600 & n601;
  assign n78308 = n585 ^ n590;
  assign n584 = ~n590;
  assign n593 = ~n595;
  assign n574 = n584 & n585;
  assign n586 = n593 & n594;
  assign n581 = n586 ^ n587;
  assign n588 = ~n586;
  assign n575 = n581 ^ n582;
  assign n583 = n588 & n589;
  assign n78307 = n574 ^ n575;
  assign n576 = ~n575;
  assign n579 = ~n583;
  assign n561 = n576 & n574;
  assign n577 = n579 & n580;
  assign n567 = n577 ^ n578;
  assign n572 = ~n577;
  assign n562 = n567 ^ n568;
  assign n571 = n572 & n573;
  assign n78306 = n561 ^ n562;
  assign n560 = ~n562;
  assign n569 = ~n571;
  assign n552 = n560 & n561;
  assign n563 = n569 & n570;
  assign n556 = n563 ^ n564;
  assign n565 = ~n563;
  assign n553 = n555 ^ n556;
  assign n559 = n565 & n566;
  assign n78305 = n552 ^ n553;
  assign n554 = ~n553;
  assign n557 = ~n559;
  assign n537 = n554 & n552;
  assign n548 = n557 & n558;
  assign n536 = ~n537;
  assign n545 = n548 ^ n549;
  assign n550 = ~n548;
  assign n538 = n545 ^ n546;
  assign n547 = n550 & n551;
  assign n78304 = n537 ^ n538;
  assign n535 = ~n538;
  assign n543 = ~n547;
  assign n533 = n535 & n536;
  assign n540 = n543 & n544;
  assign n532 = ~n533;
  assign n531 = n539 ^ n540;
  assign n541 = ~n540;
  assign n517 = n531 & n532;
  assign n78303 = n533 ^ n531;
  assign n534 = n541 & n542;
  assign n529 = ~n534;
  assign n527 = n529 & n530;
  assign n523 = n527 ^ n528;
  assign n525 = ~n527;
  assign n518 = n522 ^ n523;
  assign n524 = n525 & n526;
  assign n78302 = n517 ^ n518;
  assign n516 = ~n518;
  assign n520 = ~n524;
  assign n512 = n516 & n517;
  assign n519 = n520 & n521;
  assign n515 = ~n519;
  assign n513 = n514 ^ n515;
  assign n78301 = n512 ^ n513;
endmodule
