module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10;
  wire n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669;
  assign n11 = ~x5 & ~x6;
  assign n20 = ~x0 & x7;
  assign n21 = ~x2 & ~x8;
  assign n22 = x2 & x8;
  assign n23 = ~x9 & n22;
  assign n24 = ~n21 & ~n23;
  assign n25 = n20 & ~n24;
  assign n26 = x0 & x9;
  assign n27 = ~x2 & x8;
  assign n28 = n26 & n27;
  assign n29 = ~n25 & ~n28;
  assign n30 = ~x3 & ~n29;
  assign n31 = x8 & x9;
  assign n32 = x2 & ~x3;
  assign n33 = n31 & n32;
  assign n34 = ~x8 & ~x9;
  assign n35 = ~x2 & x3;
  assign n36 = n34 & n35;
  assign n37 = ~n33 & ~n36;
  assign n38 = ~x0 & ~n37;
  assign n39 = x3 & ~x9;
  assign n40 = x2 & ~n39;
  assign n41 = x0 & ~n35;
  assign n42 = ~n34 & n41;
  assign n43 = ~n40 & n42;
  assign n44 = ~n38 & ~n43;
  assign n45 = ~x7 & ~n44;
  assign n46 = ~n30 & ~n45;
  assign n47 = ~x1 & ~n46;
  assign n12 = ~x7 & ~x8;
  assign n13 = ~x2 & ~x3;
  assign n14 = ~x7 & ~x9;
  assign n15 = n13 & ~n14;
  assign n16 = ~x8 & x9;
  assign n17 = n16 ^ x0;
  assign n18 = n15 & n17;
  assign n19 = ~n12 & ~n18;
  assign n48 = n47 ^ n19;
  assign n49 = n11 & ~n48;
  assign n50 = ~x1 & ~x8;
  assign n51 = ~x3 & ~n50;
  assign n52 = ~x1 & x2;
  assign n53 = x8 & ~n52;
  assign n54 = x0 & ~n53;
  assign n55 = ~n51 & n54;
  assign n56 = ~x5 & ~x9;
  assign n58 = x8 ^ x2;
  assign n57 = x8 ^ x3;
  assign n59 = n58 ^ n57;
  assign n60 = x8 ^ x1;
  assign n61 = n60 ^ n57;
  assign n62 = n57 & ~n61;
  assign n63 = n62 ^ n57;
  assign n64 = n59 & n63;
  assign n65 = n64 ^ n62;
  assign n66 = n65 ^ x8;
  assign n67 = n66 ^ n57;
  assign n68 = ~x0 & ~n67;
  assign n69 = n56 & ~n68;
  assign n70 = ~n55 & n69;
  assign n71 = ~x5 & x8;
  assign n72 = x0 & x1;
  assign n73 = x8 & n72;
  assign n74 = x8 ^ x5;
  assign n75 = n74 ^ x8;
  assign n76 = ~x1 & ~x2;
  assign n77 = n76 ^ x8;
  assign n78 = ~n75 & ~n77;
  assign n79 = n78 ^ x8;
  assign n80 = ~n13 & n79;
  assign n81 = ~n73 & ~n80;
  assign n82 = ~n71 & ~n81;
  assign n83 = ~x5 & ~n35;
  assign n84 = x5 & ~x8;
  assign n85 = ~x0 & ~x1;
  assign n86 = ~n84 & n85;
  assign n87 = ~n83 & n86;
  assign n88 = n31 & ~n32;
  assign n89 = x5 & x9;
  assign n90 = ~n26 & ~n89;
  assign n91 = ~n88 & n90;
  assign n92 = ~n87 & ~n91;
  assign n93 = ~n82 & n92;
  assign n94 = n13 & n85;
  assign n95 = x5 & n34;
  assign n96 = ~n94 & n95;
  assign n97 = x6 & ~x7;
  assign n98 = ~n96 & n97;
  assign n99 = ~n93 & n98;
  assign n100 = ~n70 & n99;
  assign n101 = ~x3 & ~n22;
  assign n102 = x0 & ~x1;
  assign n103 = ~x1 & x9;
  assign n104 = n103 ^ x2;
  assign n105 = n102 & n104;
  assign n106 = n101 & ~n105;
  assign n107 = x0 & ~x2;
  assign n108 = ~x9 & n107;
  assign n109 = x2 & n16;
  assign n110 = ~n108 & ~n109;
  assign n111 = x1 & ~n110;
  assign n112 = x3 & ~n27;
  assign n113 = ~n111 & n112;
  assign n114 = ~n106 & ~n113;
  assign n115 = x9 ^ x0;
  assign n116 = x1 & ~n115;
  assign n117 = x8 & ~n116;
  assign n118 = x5 & ~x6;
  assign n119 = ~x7 & n118;
  assign n120 = ~n117 & n119;
  assign n121 = ~n114 & n120;
  assign n122 = ~n100 & ~n121;
  assign n123 = ~n49 & n122;
  assign n125 = x6 ^ x5;
  assign n124 = n94 ^ x4;
  assign n126 = n125 ^ n124;
  assign n127 = n125 ^ n34;
  assign n128 = n125 & n127;
  assign n129 = n128 ^ n125;
  assign n130 = ~n126 & n129;
  assign n131 = n130 ^ n128;
  assign n132 = n131 ^ n125;
  assign n133 = n132 ^ n34;
  assign n134 = n94 & n133;
  assign n135 = n134 ^ n124;
  assign n136 = ~n123 & ~n135;
  assign n152 = n22 & n102;
  assign n153 = n21 & n85;
  assign n154 = n14 & ~n153;
  assign n155 = ~n152 & n154;
  assign n137 = ~x3 & ~x9;
  assign n138 = ~x0 & x8;
  assign n139 = x1 & ~x2;
  assign n140 = n138 & n139;
  assign n141 = ~x7 & x8;
  assign n142 = ~n21 & ~n141;
  assign n143 = n102 & ~n142;
  assign n144 = ~n140 & ~n143;
  assign n145 = n137 & ~n144;
  assign n146 = ~n85 & ~n107;
  assign n147 = ~x3 & ~n76;
  assign n148 = n31 ^ x7;
  assign n149 = n147 & n148;
  assign n150 = ~n146 & n149;
  assign n151 = ~n145 & ~n150;
  assign n156 = n155 ^ n151;
  assign n157 = n11 & ~n156;
  assign n158 = ~x1 & ~x5;
  assign n159 = x9 ^ x8;
  assign n160 = x3 ^ x0;
  assign n161 = n160 ^ x0;
  assign n162 = ~n115 & n161;
  assign n163 = n162 ^ x0;
  assign n164 = n159 & n163;
  assign n165 = n164 ^ x3;
  assign n166 = n158 & ~n165;
  assign n167 = x9 ^ x3;
  assign n168 = x1 & ~n167;
  assign n169 = ~x9 & ~n71;
  assign n170 = n168 & ~n169;
  assign n171 = x2 & ~n89;
  assign n172 = ~n170 & n171;
  assign n173 = ~n166 & n172;
  assign n174 = n13 & n72;
  assign n175 = ~x2 & ~n56;
  assign n176 = ~n174 & ~n175;
  assign n177 = x1 & ~n138;
  assign n178 = n89 & n177;
  assign n179 = ~n176 & ~n178;
  assign n180 = ~x3 & ~n85;
  assign n181 = n16 & n72;
  assign n182 = n180 & ~n181;
  assign n183 = n16 & n102;
  assign n184 = x3 & ~n89;
  assign n185 = ~n183 & n184;
  assign n186 = ~n182 & ~n185;
  assign n187 = n179 & ~n186;
  assign n188 = n97 & ~n187;
  assign n189 = ~n173 & n188;
  assign n190 = ~x3 & n152;
  assign n191 = x2 & x3;
  assign n192 = n16 & n191;
  assign n193 = ~n137 & ~n192;
  assign n194 = x1 & ~n193;
  assign n195 = ~n190 & ~n194;
  assign n196 = ~n31 & ~n103;
  assign n197 = x9 & ~n13;
  assign n198 = n196 & ~n197;
  assign n199 = ~x0 & n198;
  assign n200 = x1 & ~n27;
  assign n201 = ~x9 & ~n32;
  assign n202 = ~n200 & n201;
  assign n203 = ~n199 & ~n202;
  assign n204 = n195 & n203;
  assign n205 = n119 & ~n204;
  assign n206 = ~n189 & ~n205;
  assign n207 = ~n157 & n206;
  assign n208 = ~x4 & ~n34;
  assign n209 = n94 & n208;
  assign n210 = ~x0 & ~x6;
  assign n211 = ~x9 & ~n210;
  assign n212 = ~x3 & n76;
  assign n213 = ~n211 & n212;
  assign n214 = x4 & ~n213;
  assign n215 = ~n209 & ~n214;
  assign n216 = ~n207 & n215;
  assign n253 = x1 & x9;
  assign n254 = x6 ^ x2;
  assign n255 = x8 ^ x6;
  assign n256 = n254 & n255;
  assign n257 = n256 ^ x2;
  assign n258 = n253 & ~n257;
  assign n259 = ~x0 & ~n258;
  assign n260 = ~x3 & x9;
  assign n261 = x0 & ~n21;
  assign n262 = n260 & ~n261;
  assign n247 = x1 & ~x6;
  assign n263 = x8 & ~x9;
  assign n264 = n247 & ~n263;
  assign n230 = x2 & ~x6;
  assign n265 = ~x3 & ~n230;
  assign n266 = ~n264 & n265;
  assign n267 = ~n262 & ~n266;
  assign n268 = ~n259 & ~n267;
  assign n269 = ~x7 & ~n268;
  assign n217 = x0 & ~n34;
  assign n218 = n139 & n217;
  assign n219 = ~x6 & x8;
  assign n220 = ~x1 & ~n219;
  assign n221 = n108 & n220;
  assign n222 = ~x0 & x2;
  assign n223 = n31 & n222;
  assign n224 = ~n221 & ~n223;
  assign n225 = ~n218 & n224;
  assign n226 = ~x2 & ~x6;
  assign n227 = ~x8 & ~n210;
  assign n228 = ~n226 & ~n227;
  assign n229 = x1 & ~x9;
  assign n231 = x0 & ~n230;
  assign n232 = n229 & ~n231;
  assign n233 = ~n228 & n232;
  assign n234 = ~x9 & ~n22;
  assign n235 = ~x6 & ~n31;
  assign n236 = n85 & ~n235;
  assign n237 = ~n234 & n236;
  assign n238 = ~n233 & ~n237;
  assign n239 = n225 & n238;
  assign n240 = ~x5 & ~x7;
  assign n241 = x0 & n229;
  assign n242 = n11 & ~n16;
  assign n243 = ~n241 & n242;
  assign n244 = ~n240 & ~n243;
  assign n245 = ~x3 & ~n20;
  assign n246 = ~n137 & ~n245;
  assign n248 = ~x0 & n14;
  assign n249 = n247 & n248;
  assign n250 = ~n246 & ~n249;
  assign n251 = ~n244 & n250;
  assign n252 = ~n239 & n251;
  assign n270 = n269 ^ n252;
  assign n276 = ~x1 & x8;
  assign n272 = ~x5 & x6;
  assign n277 = ~x6 & x9;
  assign n278 = ~n272 & ~n277;
  assign n279 = n276 & ~n278;
  assign n280 = ~n23 & n71;
  assign n281 = ~n138 & ~n280;
  assign n282 = ~n279 & n281;
  assign n283 = x2 & ~x5;
  assign n284 = ~n226 & ~n283;
  assign n285 = ~x1 & n284;
  assign n286 = n229 & n283;
  assign n287 = x5 & x6;
  assign n288 = ~x0 & ~n287;
  assign n289 = ~n175 & n288;
  assign n290 = ~n286 & n289;
  assign n291 = ~n285 & n290;
  assign n292 = ~n282 & ~n291;
  assign n293 = x1 & x6;
  assign n294 = n293 ^ x0;
  assign n295 = n293 ^ x9;
  assign n296 = n295 ^ x9;
  assign n297 = n283 ^ x9;
  assign n298 = n296 & n297;
  assign n299 = n298 ^ x9;
  assign n300 = n294 & n299;
  assign n301 = n284 ^ x0;
  assign n302 = n301 ^ x0;
  assign n303 = n302 ^ x8;
  assign n304 = x5 & n229;
  assign n305 = n304 ^ x9;
  assign n306 = ~x0 & n305;
  assign n307 = n306 ^ n304;
  assign n308 = n303 & ~n307;
  assign n309 = n308 ^ n306;
  assign n310 = n309 ^ n304;
  assign n311 = n310 ^ x0;
  assign n312 = ~x8 & n311;
  assign n313 = ~n300 & n312;
  assign n314 = ~n292 & ~n313;
  assign n271 = ~x2 & n85;
  assign n273 = ~x8 & n272;
  assign n274 = n271 & ~n273;
  assign n275 = n274 ^ x4;
  assign n315 = n314 ^ n275;
  assign n316 = n315 ^ n275;
  assign n317 = n275 ^ n274;
  assign n318 = ~n316 & ~n317;
  assign n319 = n318 ^ n275;
  assign n320 = x3 & ~n319;
  assign n321 = n320 ^ n275;
  assign n322 = n270 & ~n321;
  assign n323 = ~x0 & x5;
  assign n324 = ~n219 & n323;
  assign n325 = ~x5 & ~n263;
  assign n326 = x0 & ~n277;
  assign n327 = n325 & n326;
  assign n328 = ~n324 & ~n327;
  assign n329 = x1 & ~n328;
  assign n330 = x0 & x5;
  assign n331 = x1 & ~n330;
  assign n332 = ~x6 & n31;
  assign n333 = ~n331 & n332;
  assign n334 = n102 & ~n118;
  assign n335 = ~n325 & n334;
  assign n336 = ~n333 & ~n335;
  assign n337 = ~n329 & n336;
  assign n338 = ~n104 & ~n287;
  assign n339 = x3 & ~n338;
  assign n340 = ~n337 & n339;
  assign n341 = n34 ^ x2;
  assign n342 = n341 ^ n34;
  assign n343 = n159 ^ n34;
  assign n344 = ~n342 & n343;
  assign n345 = n344 ^ n34;
  assign n346 = x1 & n345;
  assign n347 = n76 ^ x1;
  assign n348 = n347 ^ x1;
  assign n349 = n34 ^ x1;
  assign n350 = n349 ^ x1;
  assign n351 = n348 & n350;
  assign n352 = n351 ^ x1;
  assign n353 = ~x6 & n352;
  assign n354 = n353 ^ x1;
  assign n355 = ~n346 & ~n354;
  assign n356 = n330 & ~n355;
  assign n357 = ~n103 & ~n138;
  assign n358 = x6 & ~n229;
  assign n359 = ~n357 & n358;
  assign n360 = ~x5 & ~n359;
  assign n361 = n31 & n85;
  assign n362 = ~x6 & ~n361;
  assign n363 = ~n230 & ~n362;
  assign n364 = n360 & n363;
  assign n365 = n22 & n253;
  assign n366 = ~x6 & ~n365;
  assign n367 = ~n293 & n323;
  assign n368 = x2 & n272;
  assign n369 = ~n367 & ~n368;
  assign n370 = ~n366 & ~n369;
  assign n371 = ~n138 & n286;
  assign n372 = ~x3 & ~n371;
  assign n373 = ~n370 & n372;
  assign n374 = ~n364 & n373;
  assign n375 = ~n356 & n374;
  assign n376 = ~n125 & n212;
  assign n377 = n376 ^ x4;
  assign n378 = ~x7 & ~n377;
  assign n379 = ~n375 & n378;
  assign n380 = ~n340 & n379;
  assign n381 = ~x7 & n287;
  assign n382 = n85 ^ x2;
  assign n383 = n85 ^ x4;
  assign n384 = n383 ^ x4;
  assign n385 = n212 ^ x4;
  assign n386 = n385 ^ x4;
  assign n387 = n384 & n386;
  assign n388 = n387 ^ x4;
  assign n389 = n382 & ~n388;
  assign n390 = n381 & n389;
  assign n391 = x3 & ~x4;
  assign n392 = ~n271 & n391;
  assign n393 = x4 & n94;
  assign n394 = ~n392 & ~n393;
  assign n395 = n381 & ~n394;
  assign n396 = ~x3 & ~x4;
  assign n456 = ~x2 & n240;
  assign n457 = ~n34 & n456;
  assign n458 = x6 & ~n457;
  assign n459 = x0 & ~n458;
  assign n460 = n365 ^ x5;
  assign n461 = n460 ^ n365;
  assign n462 = n461 ^ x7;
  assign n463 = n277 ^ x2;
  assign n464 = n277 & ~n463;
  assign n465 = n464 ^ n365;
  assign n466 = n465 ^ n277;
  assign n467 = n462 & ~n466;
  assign n468 = n467 ^ n464;
  assign n469 = n468 ^ n277;
  assign n470 = ~x7 & n469;
  assign n471 = n470 ^ x5;
  assign n472 = n459 & ~n471;
  assign n473 = ~x7 & ~n34;
  assign n474 = x2 & ~n473;
  assign n475 = n14 & n71;
  assign n476 = x7 & ~x8;
  assign n477 = x1 & ~n476;
  assign n478 = ~n475 & n477;
  assign n479 = ~n474 & n478;
  assign n480 = ~x2 & ~n14;
  assign n481 = ~n95 & ~n480;
  assign n482 = x7 & n31;
  assign n483 = ~x1 & ~n482;
  assign n484 = n481 & n483;
  assign n485 = ~n479 & ~n484;
  assign n486 = n472 & ~n485;
  assign n432 = n56 & ~n293;
  assign n433 = n141 & ~n432;
  assign n434 = x2 & ~n433;
  assign n435 = x5 & ~n247;
  assign n436 = ~n253 & ~n435;
  assign n437 = ~x7 & ~n436;
  assign n438 = ~x5 & ~n31;
  assign n439 = ~x1 & ~x6;
  assign n440 = ~n141 & n439;
  assign n441 = n438 & n440;
  assign n442 = ~n437 & ~n441;
  assign n443 = n434 & n442;
  assign n444 = n12 & n293;
  assign n445 = ~x2 & ~n381;
  assign n446 = ~n444 & n445;
  assign n447 = n11 ^ x7;
  assign n448 = ~x8 & ~n447;
  assign n449 = x1 & n11;
  assign n450 = n449 ^ x9;
  assign n451 = n448 & ~n450;
  assign n452 = n451 ^ n449;
  assign n453 = ~x9 & n452;
  assign n454 = n446 & ~n453;
  assign n455 = ~n443 & ~n454;
  assign n487 = n486 ^ n455;
  assign n397 = ~n72 & n84;
  assign n398 = ~n139 & n397;
  assign n399 = ~n108 & n398;
  assign n400 = n103 & n222;
  assign n401 = x5 & x8;
  assign n402 = ~n229 & n401;
  assign n403 = ~n400 & n402;
  assign n404 = ~x4 & ~n403;
  assign n405 = ~n399 & n404;
  assign n406 = n405 ^ x5;
  assign n407 = n405 ^ x6;
  assign n408 = n407 ^ x6;
  assign n409 = ~n22 & ~n277;
  assign n410 = x0 & ~n409;
  assign n411 = ~x1 & ~n16;
  assign n412 = ~x2 & x6;
  assign n413 = ~x0 & ~x9;
  assign n414 = n413 ^ n138;
  assign n415 = n412 & n414;
  assign n416 = n415 ^ n413;
  assign n417 = n411 & ~n416;
  assign n418 = ~n410 & n417;
  assign n419 = ~x0 & n31;
  assign n420 = ~n257 & n419;
  assign n421 = ~x2 & ~n138;
  assign n422 = n211 & n421;
  assign n423 = x1 & ~n422;
  assign n424 = ~n420 & n423;
  assign n425 = ~n418 & ~n424;
  assign n426 = n425 ^ x6;
  assign n427 = n408 & n426;
  assign n428 = n427 ^ x6;
  assign n429 = n406 & ~n428;
  assign n430 = n429 ^ x5;
  assign n431 = ~n393 & ~n430;
  assign n488 = n487 ^ n431;
  assign n489 = n488 ^ n487;
  assign n490 = n487 ^ x7;
  assign n491 = n490 ^ n487;
  assign n492 = ~n489 & ~n491;
  assign n493 = n492 ^ n487;
  assign n494 = ~n396 & n493;
  assign n495 = n494 ^ n487;
  assign n496 = ~n51 & ~n276;
  assign n497 = ~n196 & n496;
  assign n498 = x8 & n116;
  assign n499 = ~x3 & ~n498;
  assign n500 = ~n85 & ~n419;
  assign n501 = ~n499 & n500;
  assign n502 = ~n497 & n501;
  assign n503 = ~x2 & ~n502;
  assign n504 = n22 & n167;
  assign n505 = x0 & ~x8;
  assign n506 = ~n260 & n505;
  assign n507 = ~n35 & n506;
  assign n508 = ~n504 & ~n507;
  assign n509 = x1 & ~n508;
  assign n510 = n159 & n439;
  assign n511 = ~x0 & n13;
  assign n512 = n511 ^ x3;
  assign n513 = n510 & ~n512;
  assign n514 = n118 & ~n513;
  assign n515 = ~n509 & n514;
  assign n516 = ~n503 & n515;
  assign n556 = n34 & n180;
  assign n557 = n196 & ~n276;
  assign n558 = ~n556 & n557;
  assign n559 = ~n103 & n217;
  assign n560 = ~n558 & ~n559;
  assign n561 = ~x2 & ~n560;
  assign n562 = x2 & ~n34;
  assign n563 = ~x0 & x3;
  assign n564 = ~n159 & n563;
  assign n565 = ~n562 & ~n564;
  assign n566 = ~x1 & ~n565;
  assign n567 = ~n33 & ~n566;
  assign n568 = ~n561 & n567;
  assign n518 = x2 ^ x0;
  assign n524 = x1 ^ x0;
  assign n525 = n524 ^ n167;
  assign n526 = n525 ^ x3;
  assign n517 = n167 ^ x1;
  assign n519 = n518 ^ n517;
  assign n527 = n526 ^ n519;
  assign n528 = n527 ^ n518;
  assign n529 = n518 & n528;
  assign n530 = n529 ^ n167;
  assign n531 = n530 ^ n519;
  assign n532 = n531 ^ n518;
  assign n533 = n532 ^ x3;
  assign n534 = n519 ^ n518;
  assign n535 = n534 ^ x3;
  assign n536 = n531 & n535;
  assign n537 = n536 ^ n167;
  assign n538 = n537 ^ n519;
  assign n539 = n538 ^ n518;
  assign n540 = n539 ^ x3;
  assign n541 = n533 & n540;
  assign n520 = n519 ^ n167;
  assign n521 = n520 ^ n518;
  assign n522 = n521 ^ x3;
  assign n523 = n521 & n522;
  assign n542 = n541 ^ n523;
  assign n543 = n542 ^ n529;
  assign n544 = n543 ^ n167;
  assign n545 = n544 ^ n519;
  assign n546 = n545 ^ n518;
  assign n547 = n546 ^ x3;
  assign n548 = x8 & n547;
  assign n549 = n32 & n253;
  assign n550 = ~n101 & ~n413;
  assign n551 = x3 & ~n21;
  assign n552 = ~x1 & ~n551;
  assign n553 = ~n550 & n552;
  assign n554 = ~n549 & ~n553;
  assign n555 = ~n548 & n554;
  assign n569 = n568 ^ n555;
  assign n570 = n569 ^ n568;
  assign n571 = n568 ^ x6;
  assign n572 = n571 ^ n568;
  assign n573 = ~n570 & ~n572;
  assign n574 = n573 ^ n568;
  assign n575 = ~x4 & ~n574;
  assign n576 = n575 ^ x6;
  assign n577 = ~x5 & ~n576;
  assign n578 = ~n516 & ~n577;
  assign n579 = x4 & ~n94;
  assign n580 = x7 & ~n513;
  assign n581 = n14 & n27;
  assign n582 = ~n476 & ~n581;
  assign n583 = x0 & n439;
  assign n584 = ~n582 & n583;
  assign n585 = ~n580 & ~n584;
  assign n586 = ~n579 & n585;
  assign n587 = ~n578 & n586;
  assign n588 = n240 & n393;
  assign n589 = ~n11 & ~n235;
  assign n590 = ~n26 & ~n304;
  assign n591 = n102 & ~n263;
  assign n592 = n357 & ~n591;
  assign n593 = n590 & n592;
  assign n594 = ~x2 & ~n593;
  assign n595 = ~x1 & ~n234;
  assign n596 = ~n438 & n595;
  assign n597 = n372 & ~n596;
  assign n598 = ~n594 & n597;
  assign n599 = ~n589 & n598;
  assign n600 = ~n271 & ~n439;
  assign n601 = ~x9 & ~n227;
  assign n602 = ~n600 & n601;
  assign n603 = x9 & n254;
  assign n604 = ~n177 & n603;
  assign n605 = n226 & ~n276;
  assign n606 = x3 & ~x5;
  assign n607 = ~n605 & n606;
  assign n608 = ~n604 & n607;
  assign n609 = ~n602 & n608;
  assign n610 = n35 & n118;
  assign n611 = n557 ^ n85;
  assign n612 = n611 ^ n557;
  assign n613 = n557 ^ n31;
  assign n614 = n612 & n613;
  assign n615 = n614 ^ n557;
  assign n616 = n610 & ~n615;
  assign n617 = ~n609 & ~n616;
  assign n618 = ~n599 & n617;
  assign n619 = n11 & ~n31;
  assign n620 = ~x2 & ~n229;
  assign n621 = n85 & n562;
  assign n622 = ~n620 & ~n621;
  assign n623 = n619 & ~n622;
  assign n624 = x7 & ~n623;
  assign n625 = ~x4 & ~n624;
  assign n626 = ~n618 & n625;
  assign n627 = ~n588 & ~n626;
  assign n628 = ~n360 & ~n362;
  assign n629 = ~x1 & ~n34;
  assign n630 = n500 & ~n629;
  assign n631 = n11 & n630;
  assign n632 = ~n628 & ~n631;
  assign n633 = x5 ^ x2;
  assign n634 = n633 ^ x6;
  assign n635 = n287 & ~n634;
  assign n636 = n635 ^ n634;
  assign n637 = ~n632 & n636;
  assign n638 = x3 & ~x7;
  assign n639 = ~n637 & n638;
  assign n640 = n230 & n557;
  assign n641 = ~n11 & ~n76;
  assign n642 = ~n640 & n641;
  assign n643 = x7 ^ x2;
  assign n644 = n524 ^ x0;
  assign n645 = ~x9 & ~n138;
  assign n646 = n645 ^ x0;
  assign n647 = n644 & ~n646;
  assign n648 = n647 ^ x0;
  assign n649 = n648 ^ x7;
  assign n650 = n643 & ~n649;
  assign n651 = n650 ^ n647;
  assign n652 = n651 ^ x0;
  assign n653 = n652 ^ x2;
  assign n654 = ~x7 & ~n653;
  assign n655 = n654 ^ x7;
  assign n656 = n655 ^ x7;
  assign n657 = ~n621 & ~n656;
  assign n658 = n22 & n103;
  assign n659 = ~x3 & ~n658;
  assign n660 = ~n376 & n659;
  assign n661 = ~n657 & n660;
  assign n662 = ~n642 & n661;
  assign n663 = ~n639 & ~n662;
  assign n664 = ~n385 & ~n663;
  assign n665 = n191 & n630;
  assign n666 = ~x4 & ~n665;
  assign n667 = ~x7 & n11;
  assign n668 = ~n579 & n667;
  assign n669 = ~n666 & n668;
  assign y0 = n136;
  assign y1 = n216;
  assign y2 = n322;
  assign y3 = n380;
  assign y4 = n390;
  assign y5 = n395;
  assign y6 = ~n495;
  assign y7 = ~n587;
  assign y8 = n627;
  assign y9 = n664;
  assign y10 = n669;
endmodule
