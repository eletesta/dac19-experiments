module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, y0, y1, y2, y3, y4, y5, y6);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10;
  output y0, y1, y2, y3, y4, y5, y6;
  wire n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159;
  assign n12 = x1 & x4;
  assign n13 = n12 ^ x0;
  assign n14 = ~x5 & n13;
  assign n15 = x2 ^ x1;
  assign n16 = x5 & n15;
  assign n17 = ~x6 & ~n16;
  assign n18 = ~n14 & n17;
  assign n19 = x3 ^ x2;
  assign n20 = x6 & ~n19;
  assign n21 = ~x7 & ~n20;
  assign n22 = ~n18 & n21;
  assign n23 = x4 ^ x3;
  assign n24 = x7 & n23;
  assign n25 = ~x8 & ~n24;
  assign n26 = ~n22 & n25;
  assign n27 = x5 ^ x4;
  assign n28 = x8 & ~n27;
  assign n29 = ~n26 & ~n28;
  assign n30 = ~x9 & ~n29;
  assign n31 = x6 ^ x5;
  assign n32 = x9 & ~n31;
  assign n33 = ~x10 & ~n32;
  assign n34 = ~n30 & n33;
  assign n35 = x8 & x9;
  assign n36 = x6 & x7;
  assign n37 = ~n35 & n36;
  assign n38 = ~x6 & ~x7;
  assign n39 = x10 & ~n38;
  assign n40 = ~n37 & n39;
  assign n41 = ~n34 & ~n40;
  assign n46 = x2 & x4;
  assign n44 = ~x0 & n12;
  assign n45 = n44 ^ x1;
  assign n47 = n46 ^ n45;
  assign n42 = x1 & x2;
  assign n43 = n42 ^ x3;
  assign n48 = n47 ^ n43;
  assign n49 = x5 & n48;
  assign n50 = n49 ^ n47;
  assign n51 = ~x6 & ~n50;
  assign n52 = x2 & x3;
  assign n53 = n52 ^ x4;
  assign n54 = x6 & ~x9;
  assign n55 = ~n53 & n54;
  assign n56 = ~n51 & ~n55;
  assign n57 = ~x7 & ~x8;
  assign n58 = ~n56 & n57;
  assign n59 = x4 & x5;
  assign n60 = n59 ^ x6;
  assign n61 = x8 & ~n60;
  assign n62 = ~x9 & ~n61;
  assign n63 = x3 & x4;
  assign n64 = n63 ^ x5;
  assign n65 = x7 & ~x8;
  assign n66 = ~n64 & n65;
  assign n67 = n62 & ~n66;
  assign n68 = x5 & x6;
  assign n69 = n68 ^ x7;
  assign n70 = x9 & n69;
  assign n71 = ~n67 & ~n70;
  assign n72 = ~x10 & ~n71;
  assign n73 = ~n58 & n72;
  assign n74 = x8 & n36;
  assign n75 = ~x9 & n74;
  assign n76 = ~x8 & ~n36;
  assign n77 = x10 & ~n76;
  assign n78 = ~n75 & n77;
  assign n79 = ~n73 & ~n78;
  assign n80 = x6 & n59;
  assign n81 = n52 & n80;
  assign n82 = ~x7 & ~n81;
  assign n83 = x3 & ~x6;
  assign n84 = ~x5 & ~n83;
  assign n85 = ~x4 & ~x6;
  assign n86 = ~n84 & ~n85;
  assign n87 = x6 & ~n63;
  assign n88 = x2 & ~n87;
  assign n89 = ~n86 & ~n88;
  assign n90 = n82 & ~n89;
  assign n91 = ~x0 & ~x5;
  assign n92 = x1 & ~n91;
  assign n93 = ~x3 & x5;
  assign n94 = n92 & ~n93;
  assign n96 = ~x4 & n31;
  assign n97 = x4 & ~x5;
  assign n98 = ~x3 & n97;
  assign n99 = ~n96 & ~n98;
  assign n95 = n46 & n83;
  assign n100 = n99 ^ n95;
  assign n101 = n94 & ~n100;
  assign n102 = n101 ^ n99;
  assign n103 = n90 & n102;
  assign n104 = ~x3 & n36;
  assign n105 = ~n103 & ~n104;
  assign n106 = ~x8 & ~n105;
  assign n107 = x7 & ~n80;
  assign n108 = ~n76 & n107;
  assign n109 = ~x7 & x8;
  assign n110 = ~n83 & ~n109;
  assign n111 = ~n38 & n59;
  assign n112 = ~n110 & n111;
  assign n113 = ~n108 & ~n112;
  assign n114 = ~n106 & n113;
  assign n115 = ~x9 & ~x10;
  assign n116 = ~n114 & n115;
  assign n117 = ~x9 & ~n74;
  assign n118 = x10 & ~n117;
  assign n119 = x5 & n36;
  assign n120 = n119 ^ x8;
  assign n121 = x9 & n120;
  assign n122 = ~n118 & ~n121;
  assign n123 = ~n116 & n122;
  assign n124 = ~x5 & ~x6;
  assign n125 = n57 & n124;
  assign n126 = ~x4 & n125;
  assign n127 = ~x2 & n59;
  assign n128 = n74 & n127;
  assign n129 = ~n126 & ~n128;
  assign n130 = ~x3 & n115;
  assign n131 = ~n129 & n130;
  assign n132 = n92 & n124;
  assign n133 = n52 & n132;
  assign n134 = n42 & n63;
  assign n135 = ~x6 & ~n97;
  assign n136 = ~n134 & n135;
  assign n137 = ~n133 & ~n136;
  assign n138 = n82 & n137;
  assign n139 = ~x8 & ~n138;
  assign n140 = ~x2 & ~x3;
  assign n141 = n59 & ~n140;
  assign n142 = n36 & n141;
  assign n143 = ~x9 & ~n142;
  assign n144 = ~n139 & n143;
  assign n145 = x9 ^ x8;
  assign n146 = ~x9 & ~n63;
  assign n147 = ~n145 & n146;
  assign n148 = n147 ^ n145;
  assign n149 = n119 & ~n148;
  assign n150 = ~x10 & ~n149;
  assign n151 = ~n144 & n150;
  assign n152 = n94 & n95;
  assign n153 = n124 & ~n152;
  assign n154 = n57 & ~n81;
  assign n155 = ~n153 & n154;
  assign n156 = x8 & n142;
  assign n157 = n115 & ~n156;
  assign n158 = ~n155 & n157;
  assign n159 = n115 & n154;
  assign y0 = ~n41;
  assign y1 = ~n79;
  assign y2 = ~n123;
  assign y3 = ~n131;
  assign y4 = ~n151;
  assign y5 = ~n158;
  assign y6 = ~n159;
endmodule
