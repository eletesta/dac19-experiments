// Benchmark "square" written by ABC on Mon Nov 19 12:52:13 2018

module square ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47,
    pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45,
    pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57,
    pi58, pi59, pi60, pi61, pi62, pi63;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127;
  wire n195, n197, n198, n199, n200, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n226, n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n245, n246,
    n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
    n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
    n271, n272, n273, n274, n276, n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290, n291, n292, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
    n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
    n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
    n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
    n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n431, n432,
    n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
    n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
    n469, n470, n471, n472, n473, n475, n476, n477, n478, n479, n480, n481,
    n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
    n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
    n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
    n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
    n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
    n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
    n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
    n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n615, n616,
    n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
    n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
    n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
    n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n677,
    n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
    n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
    n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n732, n733, n734, n735, n736, n737, n738,
    n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
    n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
    n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
    n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
    n787, n788, n789, n790, n791, n792, n793, n794, n795, n797, n798, n799,
    n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
    n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
    n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
    n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
    n848, n849, n850, n851, n852, n853, n854, n855, n857, n858, n859, n860,
    n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
    n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
    n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
    n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n924, n925, n927, n928, n929, n930, n931, n932, n933,
    n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
    n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
    n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
    n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
    n994, n995, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
    n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
    n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1146, n1147,
    n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
    n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
    n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
    n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
    n1218, n1219, n1220, n1221, n1222, n1223, n1225, n1226, n1227, n1228,
    n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
    n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
    n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
    n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
    n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
    n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
    n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
    n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
    n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
    n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
    n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
    n1400, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
    n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
    n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
    n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
    n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
    n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
    n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
    n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1491,
    n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
    n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
    n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
    n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
    n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
    n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
    n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
    n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
    n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
    n1582, n1583, n1584, n1585, n1587, n1588, n1589, n1590, n1591, n1592,
    n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
    n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
    n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
    n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
    n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
    n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
    n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
    n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
    n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
    n1683, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
    n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
    n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
    n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
    n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
    n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
    n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1782, n1783, n1784,
    n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
    n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
    n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
    n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
    n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
    n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
    n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
    n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
    n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
    n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1884, n1885,
    n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
    n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
    n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
    n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
    n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
    n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
    n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
    n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
    n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
    n1986, n1987, n1988, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
    n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
    n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
    n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
    n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
    n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
    n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
    n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
    n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
    n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
    n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
    n2097, n2098, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
    n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
    n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
    n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
    n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
    n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
    n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
    n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
    n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
    n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
    n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
    n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2218,
    n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
    n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
    n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
    n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
    n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
    n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
    n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
    n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
    n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
    n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
    n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2328, n2329,
    n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
    n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
    n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
    n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
    n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
    n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
    n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
    n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
    n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
    n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
    n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
    n2440, n2441, n2442, n2443, n2444, n2446, n2447, n2448, n2449, n2450,
    n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
    n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
    n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
    n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
    n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
    n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
    n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
    n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
    n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
    n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
    n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
    n2561, n2562, n2563, n2564, n2565, n2566, n2568, n2569, n2570, n2571,
    n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
    n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
    n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
    n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
    n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
    n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
    n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
    n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
    n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
    n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
    n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
    n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2690, n2691, n2692,
    n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
    n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
    n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
    n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
    n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
    n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
    n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
    n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
    n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
    n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
    n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
    n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2811, n2812, n2813,
    n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
    n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
    n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
    n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
    n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
    n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
    n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
    n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
    n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
    n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
    n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
    n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
    n2944, n2945, n2946, n2947, n2949, n2950, n2951, n2952, n2953, n2954,
    n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
    n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
    n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
    n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
    n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
    n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
    n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
    n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
    n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
    n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
    n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
    n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
    n3075, n3076, n3077, n3078, n3080, n3081, n3082, n3083, n3084, n3085,
    n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
    n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
    n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
    n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
    n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
    n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
    n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
    n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
    n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
    n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
    n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
    n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
    n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
    n3216, n3217, n3218, n3219, n3220, n3222, n3223, n3224, n3225, n3226,
    n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
    n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
    n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
    n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
    n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
    n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
    n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
    n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
    n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
    n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
    n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
    n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
    n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
    n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
    n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
    n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
    n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
    n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
    n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
    n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
    n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
    n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
    n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
    n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
    n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
    n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
    n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
    n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
    n3508, n3509, n3510, n3511, n3512, n3513, n3515, n3516, n3517, n3518,
    n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
    n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
    n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
    n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
    n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
    n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
    n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
    n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
    n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
    n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
    n3659, n3660, n3661, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
    n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
    n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
    n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
    n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
    n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
    n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
    n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
    n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
    n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
    n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
    n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
    n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
    n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
    n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
    n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3820,
    n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
    n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
    n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
    n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
    n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
    n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
    n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
    n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
    n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
    n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
    n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
    n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
    n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
    n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
    n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3969, n3970, n3971,
    n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
    n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
    n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
    n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
    n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
    n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
    n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
    n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
    n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
    n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
    n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
    n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
    n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
    n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
    n4112, n4113, n4114, n4115, n4116, n4117, n4119, n4120, n4121, n4122,
    n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
    n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
    n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
    n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
    n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
    n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
    n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
    n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
    n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
    n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
    n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
    n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
    n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
    n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
    n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
    n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
    n4283, n4284, n4285, n4286, n4287, n4288, n4290, n4291, n4292, n4293,
    n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
    n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
    n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
    n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
    n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
    n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
    n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
    n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
    n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
    n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
    n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
    n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
    n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
    n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
    n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
    n4444, n4445, n4446, n4447, n4448, n4450, n4451, n4452, n4453, n4454,
    n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
    n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
    n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
    n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
    n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
    n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
    n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
    n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
    n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
    n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
    n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
    n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
    n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
    n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
    n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
    n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
    n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
    n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
    n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
    n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
    n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
    n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
    n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
    n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
    n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
    n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
    n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
    n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
    n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
    n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
    n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
    n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
    n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
    n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4794, n4795, n4796,
    n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
    n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
    n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
    n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
    n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
    n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
    n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
    n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
    n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
    n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
    n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
    n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
    n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
    n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
    n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
    n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
    n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
    n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
    n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
    n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
    n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
    n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
    n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
    n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
    n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
    n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
    n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
    n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
    n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
    n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
    n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
    n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
    n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
    n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
    n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
    n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
    n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
    n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
    n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
    n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
    n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
    n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
    n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
    n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
    n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
    n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
    n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
    n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
    n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
    n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
    n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
    n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
    n5319, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
    n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
    n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
    n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
    n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
    n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
    n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
    n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
    n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
    n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
    n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
    n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
    n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
    n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
    n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
    n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
    n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
    n5490, n5491, n5492, n5493, n5494, n5496, n5497, n5498, n5499, n5500,
    n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
    n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
    n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
    n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
    n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
    n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
    n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
    n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
    n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
    n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
    n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
    n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
    n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
    n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
    n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
    n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
    n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
    n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
    n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5689, n5690, n5691,
    n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
    n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
    n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
    n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
    n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
    n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
    n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
    n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
    n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
    n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
    n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
    n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
    n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
    n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
    n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
    n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
    n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
    n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
    n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5882,
    n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
    n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
    n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
    n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
    n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
    n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
    n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
    n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
    n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
    n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
    n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
    n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
    n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
    n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
    n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
    n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
    n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
    n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
    n6063, n6064, n6065, n6066, n6067, n6068, n6070, n6071, n6072, n6073,
    n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
    n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
    n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
    n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
    n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
    n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
    n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
    n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
    n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
    n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
    n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
    n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
    n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
    n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
    n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
    n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
    n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
    n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
    n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
    n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
    n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
    n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
    n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
    n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
    n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
    n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
    n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
    n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
    n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
    n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
    n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
    n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
    n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
    n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
    n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
    n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
    n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
    n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
    n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
    n6465, n6466, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
    n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
    n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
    n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
    n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
    n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
    n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
    n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
    n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
    n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
    n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
    n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
    n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
    n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
    n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
    n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
    n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
    n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
    n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
    n6656, n6657, n6658, n6659, n6660, n6662, n6663, n6664, n6665, n6666,
    n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
    n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
    n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
    n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
    n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
    n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
    n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
    n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
    n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
    n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
    n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
    n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
    n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
    n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
    n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
    n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
    n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
    n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
    n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
    n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
    n6867, n6868, n6869, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
    n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
    n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
    n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
    n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
    n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
    n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
    n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
    n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
    n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
    n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
    n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
    n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
    n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
    n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
    n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
    n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
    n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
    n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
    n7058, n7059, n7060, n7061, n7062, n7063, n7065, n7066, n7067, n7068,
    n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
    n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
    n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
    n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
    n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
    n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
    n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
    n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
    n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
    n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
    n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
    n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
    n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
    n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
    n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
    n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
    n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
    n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
    n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
    n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7267, n7268, n7269,
    n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
    n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
    n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
    n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
    n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
    n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
    n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
    n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
    n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
    n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
    n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
    n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
    n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
    n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
    n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
    n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
    n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
    n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
    n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7460,
    n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
    n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
    n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
    n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
    n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
    n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
    n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
    n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
    n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
    n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
    n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
    n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
    n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
    n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
    n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
    n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
    n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
    n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
    n7641, n7642, n7643, n7644, n7646, n7647, n7648, n7649, n7650, n7651,
    n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
    n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
    n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
    n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
    n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
    n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
    n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
    n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
    n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
    n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
    n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
    n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
    n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
    n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
    n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
    n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
    n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
    n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
    n7832, n7833, n7834, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
    n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
    n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
    n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
    n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
    n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
    n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
    n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
    n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
    n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
    n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
    n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
    n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
    n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
    n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
    n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
    n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
    n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
    n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
    n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
    n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
    n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
    n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
    n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
    n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
    n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
    n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
    n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
    n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
    n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
    n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
    n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
    n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
    n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
    n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
    n8184, n8185, n8186, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
    n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
    n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
    n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
    n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
    n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
    n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
    n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
    n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
    n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
    n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
    n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
    n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
    n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
    n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
    n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
    n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
    n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8364, n8365,
    n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
    n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
    n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
    n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
    n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
    n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
    n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
    n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
    n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
    n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
    n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
    n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
    n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
    n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
    n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
    n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
    n8526, n8527, n8528, n8529, n8530, n8531, n8533, n8534, n8535, n8536,
    n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
    n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
    n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
    n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
    n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
    n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
    n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
    n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
    n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
    n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
    n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
    n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
    n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
    n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
    n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
    n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
    n8697, n8698, n8699, n8700, n8701, n8703, n8704, n8705, n8706, n8707,
    n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
    n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
    n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
    n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
    n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
    n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
    n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
    n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
    n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
    n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
    n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
    n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
    n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
    n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
    n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
    n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8866, n8867, n8868,
    n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
    n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
    n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
    n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
    n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
    n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
    n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
    n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
    n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
    n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
    n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
    n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
    n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
    n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
    n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
    n9019, n9020, n9021, n9022, n9023, n9024, n9026, n9027, n9028, n9029,
    n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
    n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
    n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
    n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
    n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
    n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
    n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
    n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
    n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
    n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
    n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
    n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
    n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
    n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
    n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
    n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
    n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
    n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
    n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
    n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
    n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
    n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
    n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
    n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
    n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
    n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
    n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
    n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
    n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
    n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
    n9331, n9332, n9333, n9334, n9336, n9337, n9338, n9339, n9340, n9341,
    n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
    n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
    n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
    n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
    n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
    n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
    n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
    n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
    n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
    n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
    n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
    n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
    n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
    n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
    n9482, n9483, n9484, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
    n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
    n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
    n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
    n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
    n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
    n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
    n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
    n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
    n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
    n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
    n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
    n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
    n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
    n9623, n9624, n9625, n9626, n9627, n9629, n9630, n9631, n9632, n9633,
    n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
    n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
    n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
    n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
    n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
    n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
    n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
    n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
    n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
    n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
    n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
    n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
    n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
    n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
    n9774, n9775, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
    n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
    n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
    n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
    n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
    n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
    n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
    n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
    n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
    n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
    n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
    n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
    n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
    n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
    n9915, n9916, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
    n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
    n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
    n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
    n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
    n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
    n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
    n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
    n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
    n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
    n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
    n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
    n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
    n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
    n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10059,
    n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
    n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
    n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
    n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
    n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
    n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
    n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
    n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
    n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
    n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
    n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
    n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
    n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
    n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
    n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
    n10195, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
    n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
    n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
    n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
    n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
    n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
    n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
    n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
    n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
    n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
    n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
    n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
    n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
    n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10322,
    n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
    n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
    n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
    n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
    n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
    n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
    n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
    n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
    n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
    n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
    n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
    n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
    n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
    n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
    n10449, n10450, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
    n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
    n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
    n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
    n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
    n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
    n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
    n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
    n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
    n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
    n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
    n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
    n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
    n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
    n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
    n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
    n10594, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
    n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
    n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
    n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
    n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
    n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
    n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
    n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
    n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
    n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
    n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
    n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
    n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
    n10712, n10713, n10714, n10715, n10716, n10718, n10719, n10720, n10721,
    n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
    n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
    n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
    n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
    n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
    n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
    n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
    n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
    n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
    n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
    n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
    n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
    n10830, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
    n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
    n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
    n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
    n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
    n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
    n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
    n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
    n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
    n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
    n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
    n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
    n10939, n10940, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
    n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
    n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
    n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
    n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
    n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
    n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
    n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
    n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
    n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
    n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
    n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11048,
    n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
    n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
    n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
    n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
    n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
    n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
    n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
    n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
    n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
    n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
    n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
    n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
    n11157, n11158, n11159, n11160, n11161, n11162, n11164, n11165, n11166,
    n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
    n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
    n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
    n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
    n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
    n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
    n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
    n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
    n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
    n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
    n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
    n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
    n11275, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
    n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
    n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
    n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
    n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
    n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
    n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
    n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
    n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
    n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
    n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
    n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
    n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
    n11393, n11394, n11395, n11396, n11398, n11399, n11400, n11401, n11402,
    n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
    n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
    n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
    n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
    n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
    n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
    n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
    n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
    n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
    n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
    n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
    n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
    n11511, n11512, n11513, n11515, n11516, n11517, n11518, n11519, n11520,
    n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
    n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
    n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
    n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
    n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
    n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
    n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
    n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
    n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
    n11602, n11603, n11604, n11605, n11606, n11608, n11609, n11610, n11611,
    n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
    n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
    n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
    n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
    n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
    n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
    n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
    n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
    n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
    n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
    n11702, n11703, n11704, n11705, n11707, n11708, n11709, n11710, n11711,
    n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
    n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
    n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
    n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
    n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
    n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
    n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
    n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
    n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
    n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
    n11802, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
    n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
    n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
    n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
    n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
    n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
    n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
    n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
    n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
    n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
    n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
    n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
    n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
    n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
    n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
    n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
    n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
    n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
    n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
    n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
    n11984, n11985, n11986, n11987, n11988, n11989, n11991, n11992, n11993,
    n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
    n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
    n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
    n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
    n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
    n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
    n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
    n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
    n12066, n12067, n12068, n12069, n12070, n12071, n12073, n12074, n12075,
    n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
    n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
    n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
    n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
    n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
    n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
    n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
    n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
    n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12157,
    n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
    n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
    n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
    n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
    n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
    n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
    n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
    n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
    n12230, n12231, n12232, n12234, n12235, n12236, n12237, n12238, n12239,
    n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
    n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
    n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
    n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
    n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
    n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
    n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
    n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
    n12312, n12313, n12314, n12315, n12317, n12318, n12319, n12320, n12321,
    n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
    n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
    n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
    n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
    n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
    n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
    n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
    n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
    n12394, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
    n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
    n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
    n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
    n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
    n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
    n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
    n12458, n12459, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
    n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
    n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
    n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
    n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
    n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
    n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
    n12522, n12523, n12524, n12526, n12527, n12528, n12529, n12530, n12531,
    n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
    n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
    n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
    n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
    n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
    n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
    n12586, n12587, n12588, n12590, n12591, n12592, n12593, n12594, n12595,
    n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
    n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
    n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
    n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
    n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
    n12641, n12642, n12643, n12644, n12645, n12646, n12648, n12649, n12650,
    n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
    n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
    n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
    n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
    n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
    n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
    n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
    n12714, n12715, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
    n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
    n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
    n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
    n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
    n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
    n12769, n12770, n12771, n12772, n12773, n12774, n12776, n12777, n12778,
    n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
    n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
    n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
    n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
    n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
    n12824, n12825, n12826, n12827, n12829, n12830, n12831, n12832, n12833,
    n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
    n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
    n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
    n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
    n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
    n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
    n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
    n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
    n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
    n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
    n12925, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
    n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
    n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
    n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
    n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
    n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
    n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
    n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
    n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
    n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
    n13017, n13018, n13019, n13020, n13021, n13022, n13024, n13025, n13026,
    n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
    n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
    n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
    n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
    n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
    n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
    n13081, n13082, n13083, n13085, n13086, n13087, n13088, n13089, n13090,
    n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
    n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
    n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
    n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
    n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
    n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
    n13146, n13147, n13148, n13149, n13150, n13151, n13153, n13154, n13155,
    n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
    n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
    n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13182, n13183,
    n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
    n13193, n13194, n13195, n13196, n13198, n13199, n13200, n13201, n13202,
    n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
    n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
    n13221, n13222, n13223, n13225, n13226, n13227, n13228, n13229, n13230,
    n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
    n13240, n13241, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
    n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
    n13260, n13261, n13262, n13263, n13264, n13265, n13266;
  assign po002 = ~pi00 & pi01;
  assign n195 = ~pi01 ^ pi02;
  assign po003 = ~n195 & pi00;
  assign n197 = ~pi01 & pi02;
  assign n198 = n197 & ~pi00;
  assign n199 = ~pi02 ^ pi03;
  assign n200 = ~n199 & pi00;
  assign po004 = n198 | n200;
  assign n202 = ~pi02 & pi03;
  assign n203 = pi03 & pi04;
  assign n204 = ~n202 & ~n203;
  assign n205 = ~pi02 & pi04;
  assign n206 = ~n204 & ~n205;
  assign n207 = ~n199 & pi01;
  assign n208 = ~pi03 & ~pi04;
  assign n209 = ~n207 & ~n208;
  assign n210 = ~n206 & n209;
  assign n211 = n210 & pi00;
  assign n212 = pi00 & pi01;
  assign n213 = n212 & pi04;
  assign n214 = n207 & ~n213;
  assign po005 = n211 | n214;
  assign n216 = n210 & pi01;
  assign n217 = ~n216 & n204;
  assign n218 = ~n217 ^ pi05;
  assign n219 = n218 & pi00;
  assign n220 = ~pi03 ^ ~pi04;
  assign n221 = ~n220 & pi01;
  assign n222 = ~n202 & ~pi01;
  assign n223 = ~n221 & ~n222;
  assign n224 = n223 & ~pi00;
  assign po006 = n219 | n224;
  assign n226 = ~pi03 & ~pi05;
  assign n227 = pi02 & pi04;
  assign n228 = n226 & n227;
  assign n229 = pi03 & pi05;
  assign n230 = ~n228 & ~n229;
  assign n231 = ~n230 & n212;
  assign n232 = pi00 & pi05;
  assign n233 = ~n204 & n232;
  assign n234 = po002 & n203;
  assign n235 = ~n233 & ~n234;
  assign n236 = ~n231 & n235;
  assign n237 = n220 & pi02;
  assign n238 = pi00 & pi06;
  assign n239 = pi01 & pi05;
  assign n240 = ~n238 ^ n239;
  assign n241 = ~n237 ^ ~n240;
  assign n242 = n213 & ~n226;
  assign n243 = ~n241 ^ ~n242;
  assign po007 = n236 ^ n243;
  assign n245 = n236 & ~n242;
  assign n246 = pi05 & pi06;
  assign n247 = n203 & n246;
  assign n248 = n241 & ~n247;
  assign n249 = ~n245 & ~n248;
  assign n250 = pi04 & pi06;
  assign n251 = n250 & pi01;
  assign n252 = pi02 & pi05;
  assign n253 = n251 & ~n252;
  assign n254 = pi01 & pi06;
  assign n255 = ~n254 & ~pi04;
  assign n256 = ~n253 & ~n255;
  assign n257 = n227 & ~pi06;
  assign n258 = n257 & n239;
  assign n259 = n256 & ~n258;
  assign n260 = pi03 & pi06;
  assign n261 = n260 & pi00;
  assign n262 = ~n239 ^ ~pi04;
  assign n263 = ~n261 & ~n262;
  assign n264 = ~n238 & ~pi03;
  assign n265 = ~n264 & pi02;
  assign n266 = ~n263 & n265;
  assign n267 = n212 & ~n227;
  assign n268 = n267 & n246;
  assign n269 = ~n266 & ~n268;
  assign n270 = ~n259 ^ n269;
  assign n271 = ~n203 ^ ~n252;
  assign n272 = pi00 & pi07;
  assign n273 = ~n271 ^ n272;
  assign n274 = ~n270 ^ n273;
  assign po008 = ~n249 ^ ~n274;
  assign n276 = n249 & n274;
  assign n277 = n270 & ~n273;
  assign n278 = ~n276 & ~n277;
  assign n279 = n259 & ~n269;
  assign n280 = ~n279 & ~n258;
  assign n281 = ~n251 ^ pi02;
  assign n282 = ~n281 & pi06;
  assign n283 = pi00 & pi08;
  assign n284 = ~n282 ^ ~n283;
  assign n285 = pi01 & pi07;
  assign n286 = ~n229 ^ ~n285;
  assign n287 = ~n284 ^ ~n286;
  assign n288 = n271 & ~n272;
  assign n289 = ~n203 & ~n252;
  assign n290 = ~n288 & ~n289;
  assign n291 = ~n287 ^ ~n290;
  assign n292 = ~n280 ^ n291;
  assign po009 = n278 ^ ~n292;
  assign n294 = ~n280 & n290;
  assign n295 = n278 & ~n294;
  assign n296 = n280 & ~n290;
  assign n297 = ~n295 & ~n296;
  assign n298 = pi03 & pi07;
  assign n299 = pi05 & pi08;
  assign n300 = ~n298 & n299;
  assign n301 = n300 & pi01;
  assign n302 = pi01 & pi08;
  assign n303 = ~n302 & ~pi05;
  assign n304 = ~n301 & ~n303;
  assign n305 = n239 & n298;
  assign n306 = n305 & ~pi08;
  assign n307 = n304 & ~n306;
  assign n308 = pi00 & pi09;
  assign n309 = ~n307 ^ ~n308;
  assign n310 = pi04 & pi08;
  assign n311 = n212 & n310;
  assign n312 = ~n311 & ~pi02;
  assign n313 = n283 & pi06;
  assign n314 = ~n251 & ~n313;
  assign n315 = ~n312 & ~n314;
  assign n316 = pi04 & pi05;
  assign n317 = ~n260 ^ ~n316;
  assign n318 = pi02 & pi07;
  assign n319 = ~n317 ^ ~n318;
  assign n320 = ~n315 ^ ~n319;
  assign n321 = ~n309 ^ ~n320;
  assign n322 = ~n297 ^ ~n321;
  assign n323 = ~po009 & n287;
  assign n324 = n284 & n286;
  assign n325 = ~n323 & ~n324;
  assign po010 = ~n322 ^ n325;
  assign n327 = n322 & ~n325;
  assign n328 = n297 & n321;
  assign n329 = ~n327 & ~n328;
  assign n330 = n309 & n320;
  assign n331 = n315 & n319;
  assign n332 = ~n330 & ~n331;
  assign n333 = n304 & n308;
  assign n334 = ~n333 & ~n306;
  assign n335 = pi02 & pi08;
  assign n336 = ~n298 ^ ~n335;
  assign n337 = pi00 & pi10;
  assign n338 = ~n336 ^ n337;
  assign n339 = ~n334 ^ ~n338;
  assign n340 = n317 & n318;
  assign n341 = ~n340 & ~n247;
  assign n342 = ~n299 ^ pi09;
  assign n343 = ~n342 & pi01;
  assign n344 = ~n343 ^ n250;
  assign n345 = ~n341 ^ ~n344;
  assign n346 = ~n339 ^ ~n345;
  assign n347 = ~n332 ^ n346;
  assign po011 = ~n329 ^ n347;
  assign n349 = ~n332 & n345;
  assign n350 = ~n329 & n349;
  assign n351 = n332 & ~n345;
  assign n352 = n329 & n351;
  assign n353 = ~n350 & ~n352;
  assign n354 = n353 & n339;
  assign n355 = n329 & ~n349;
  assign n356 = ~n355 & ~n351;
  assign n357 = n334 & n338;
  assign n358 = n356 & n357;
  assign n359 = ~n354 & ~n358;
  assign n360 = ~n334 & ~n338;
  assign n361 = ~n356 & n360;
  assign n362 = n359 & ~n361;
  assign n363 = ~n250 ^ pi09;
  assign n364 = ~n363 & n299;
  assign n365 = n341 & ~n364;
  assign n366 = n363 & ~n299;
  assign n367 = ~n366 & pi01;
  assign n368 = ~n365 & n367;
  assign n369 = n250 & ~pi01;
  assign n370 = ~n341 & n369;
  assign n371 = ~n368 & ~n370;
  assign n372 = pi04 & pi07;
  assign n373 = ~n246 ^ ~n372;
  assign n374 = pi00 & pi11;
  assign n375 = ~n373 ^ n374;
  assign n376 = ~n371 ^ ~n375;
  assign n377 = ~n281 & pi09;
  assign n378 = pi03 & pi08;
  assign n379 = ~n377 ^ ~n378;
  assign n380 = n336 & ~n337;
  assign n381 = ~n298 & ~n335;
  assign n382 = ~n380 & ~n381;
  assign n383 = ~n379 ^ ~n382;
  assign n384 = pi01 & pi10;
  assign n385 = ~n384 ^ pi06;
  assign n386 = ~n383 ^ ~n385;
  assign n387 = ~n376 ^ n386;
  assign po012 = ~n362 ^ n387;
  assign n389 = n329 & ~n360;
  assign n390 = ~n349 & ~n387;
  assign n391 = ~n390 & ~n357;
  assign n392 = ~n389 & n391;
  assign n393 = n349 & n387;
  assign n394 = ~n392 & ~n393;
  assign n395 = ~n387 & ~n360;
  assign n396 = ~n395 & ~n351;
  assign n397 = ~po011 & n396;
  assign n398 = n394 & ~n397;
  assign n399 = n376 & ~n386;
  assign n400 = ~n371 & ~n375;
  assign n401 = ~n399 & ~n400;
  assign n402 = n383 & n385;
  assign n403 = ~n379 & ~n382;
  assign n404 = ~n402 & ~n403;
  assign n405 = n378 & pi02;
  assign n406 = ~n251 & ~n405;
  assign n407 = ~n378 & ~pi02;
  assign n408 = ~n407 & pi09;
  assign n409 = ~n406 & n408;
  assign n410 = pi06 & pi10;
  assign n411 = n410 & pi01;
  assign n412 = ~n411 ^ ~n310;
  assign n413 = pi01 & pi11;
  assign n414 = pi05 & pi07;
  assign n415 = ~n413 ^ ~n414;
  assign n416 = ~n412 ^ ~n415;
  assign n417 = ~n409 ^ ~n416;
  assign n418 = n373 & ~n374;
  assign n419 = ~n246 & ~n372;
  assign n420 = ~n418 & ~n419;
  assign n421 = pi03 & pi09;
  assign n422 = pi02 & pi10;
  assign n423 = ~n421 ^ ~n422;
  assign n424 = pi00 & pi12;
  assign n425 = ~n423 ^ n424;
  assign n426 = ~n420 ^ n425;
  assign n427 = ~n417 ^ n426;
  assign n428 = ~n404 ^ n427;
  assign n429 = ~n401 ^ n428;
  assign po013 = n398 ^ ~n429;
  assign n431 = n398 & n429;
  assign n432 = n401 & ~n428;
  assign n433 = ~n431 & ~n432;
  assign n434 = n409 & n416;
  assign n435 = ~n404 & ~n434;
  assign n436 = ~n409 & ~n416;
  assign n437 = ~n435 & ~n436;
  assign n438 = n420 & ~n425;
  assign n439 = ~n437 & n438;
  assign n440 = ~n404 & n436;
  assign n441 = n404 & n434;
  assign n442 = ~n440 & ~n441;
  assign n443 = n442 & n426;
  assign n444 = ~n439 & ~n443;
  assign n445 = ~n420 & n425;
  assign n446 = n437 & n445;
  assign n447 = n444 & ~n446;
  assign n448 = n423 & ~n424;
  assign n449 = ~n421 & ~n422;
  assign n450 = ~n448 & ~n449;
  assign n451 = pi05 & pi11;
  assign n452 = n451 & pi01;
  assign n453 = ~n452 & pi07;
  assign n454 = pi01 & pi12;
  assign n455 = ~n453 ^ ~n454;
  assign n456 = ~n450 ^ ~n455;
  assign n457 = ~n447 ^ n456;
  assign n458 = n412 & n415;
  assign n459 = pi08 & pi10;
  assign n460 = n251 & n459;
  assign n461 = ~n458 & ~n460;
  assign n462 = pi04 & pi09;
  assign n463 = pi03 & pi10;
  assign n464 = ~n462 ^ ~n463;
  assign n465 = pi00 & pi13;
  assign n466 = ~n464 ^ n465;
  assign n467 = pi06 & pi07;
  assign n468 = ~n299 ^ ~n467;
  assign n469 = pi02 & pi11;
  assign n470 = ~n468 ^ n469;
  assign n471 = ~n466 ^ ~n470;
  assign n472 = ~n461 ^ n471;
  assign n473 = ~n457 ^ ~n472;
  assign po014 = n433 ^ n473;
  assign n475 = ~n433 & n473;
  assign n476 = ~n457 & ~n472;
  assign n477 = ~n475 & ~n476;
  assign n478 = ~n457 & n420;
  assign n479 = ~n435 & n456;
  assign n480 = ~n478 & ~n479;
  assign n481 = ~n480 & ~n436;
  assign n482 = ~n434 & ~n456;
  assign n483 = ~n457 & ~n482;
  assign n484 = ~n481 & ~n483;
  assign n485 = n450 & n455;
  assign n486 = n285 & ~pi12;
  assign n487 = n486 & n451;
  assign n488 = ~n485 & ~n487;
  assign n489 = n454 & pi07;
  assign n490 = pi05 & pi09;
  assign n491 = ~n489 ^ ~n490;
  assign n492 = pi04 & pi10;
  assign n493 = ~n491 ^ n492;
  assign n494 = pi03 & pi11;
  assign n495 = pi02 & pi12;
  assign n496 = ~n494 ^ ~n495;
  assign n497 = pi00 & pi14;
  assign n498 = ~n496 ^ n497;
  assign n499 = ~n493 ^ ~n498;
  assign n500 = ~n488 ^ ~n499;
  assign n501 = n464 & ~n465;
  assign n502 = ~n462 & ~n463;
  assign n503 = ~n501 & ~n502;
  assign n504 = n468 & ~n469;
  assign n505 = ~n299 & ~n467;
  assign n506 = ~n504 & ~n505;
  assign n507 = ~n503 ^ ~n506;
  assign n508 = pi06 & pi08;
  assign n509 = pi01 & pi13;
  assign n510 = ~n508 ^ ~n509;
  assign n511 = ~n507 ^ ~n510;
  assign n512 = ~n500 ^ n511;
  assign n513 = ~n461 & n471;
  assign n514 = ~n466 & ~n470;
  assign n515 = ~n513 & ~n514;
  assign n516 = ~n512 ^ ~n515;
  assign n517 = ~n484 ^ n516;
  assign po015 = ~n477 ^ n517;
  assign n519 = n484 & n515;
  assign n520 = n477 & ~n519;
  assign n521 = ~n484 & ~n515;
  assign n522 = ~n520 & ~n521;
  assign n523 = n500 & ~n511;
  assign n524 = ~n522 & n523;
  assign n525 = ~n500 & n511;
  assign n526 = n522 & n525;
  assign n527 = ~n524 & ~n526;
  assign n528 = n477 & n521;
  assign n529 = ~n528 & n512;
  assign n530 = ~n477 & n519;
  assign n531 = n529 & ~n530;
  assign n532 = n527 & ~n531;
  assign n533 = n488 & n499;
  assign n534 = n493 & n498;
  assign n535 = ~n533 & ~n534;
  assign n536 = n491 & ~n492;
  assign n537 = ~n489 & ~n490;
  assign n538 = ~n536 & ~n537;
  assign n539 = n496 & ~n497;
  assign n540 = ~n494 & ~n495;
  assign n541 = ~n539 & ~n540;
  assign n542 = pi05 & pi10;
  assign n543 = pi03 & pi12;
  assign n544 = ~n542 ^ ~n543;
  assign n545 = pi00 & pi15;
  assign n546 = ~n544 ^ n545;
  assign n547 = ~n541 ^ n546;
  assign n548 = ~n538 ^ n547;
  assign n549 = ~n535 ^ n548;
  assign n550 = n507 & n510;
  assign n551 = n503 & n506;
  assign n552 = ~n550 & ~n551;
  assign n553 = n508 & n509;
  assign n554 = ~n553 & pi08;
  assign n555 = pi01 & pi14;
  assign n556 = ~n554 ^ ~n555;
  assign n557 = pi04 & pi11;
  assign n558 = ~n556 ^ ~n557;
  assign n559 = pi07 & pi08;
  assign n560 = pi06 & pi09;
  assign n561 = ~n559 ^ ~n560;
  assign n562 = pi02 & pi13;
  assign n563 = ~n561 ^ n562;
  assign n564 = ~n558 ^ n563;
  assign n565 = ~n552 ^ n564;
  assign n566 = ~n549 ^ n565;
  assign po016 = ~n532 ^ ~n566;
  assign n568 = ~n566 & ~n523;
  assign n569 = n522 & ~n568;
  assign n570 = n566 & n523;
  assign n571 = ~n569 & ~n570;
  assign n572 = ~n530 & ~n566;
  assign n573 = n529 & ~n572;
  assign n574 = n571 & ~n573;
  assign n575 = n549 & ~n565;
  assign n576 = ~n535 & n548;
  assign n577 = ~n575 & ~n576;
  assign n578 = n556 & n557;
  assign n579 = n553 & ~pi14;
  assign n580 = ~n578 & ~n579;
  assign n581 = n544 & ~n545;
  assign n582 = ~n542 & ~n543;
  assign n583 = ~n581 & ~n582;
  assign n584 = ~n410 ^ ~n451;
  assign n585 = pi00 & pi16;
  assign n586 = ~n584 ^ n585;
  assign n587 = ~n583 ^ n586;
  assign n588 = ~n580 ^ n587;
  assign n589 = ~n577 ^ ~n588;
  assign n590 = ~n552 & n564;
  assign n591 = n558 & ~n563;
  assign n592 = ~n590 & ~n591;
  assign n593 = ~n538 & n547;
  assign n594 = ~n541 & n546;
  assign n595 = ~n593 & ~n594;
  assign n596 = n561 & ~n562;
  assign n597 = ~n559 & ~n560;
  assign n598 = ~n596 & ~n597;
  assign n599 = pi08 & pi14;
  assign n600 = ~n599 ^ ~pi15;
  assign n601 = n600 & pi01;
  assign n602 = pi07 & pi09;
  assign n603 = ~n601 ^ n602;
  assign n604 = ~n598 ^ n603;
  assign n605 = pi04 & pi12;
  assign n606 = pi03 & pi13;
  assign n607 = ~n605 ^ ~n606;
  assign n608 = pi02 & pi14;
  assign n609 = ~n607 ^ n608;
  assign n610 = ~n604 ^ n609;
  assign n611 = ~n595 ^ ~n610;
  assign n612 = ~n592 ^ n611;
  assign n613 = ~n589 ^ n612;
  assign po017 = ~n574 ^ n613;
  assign n615 = ~n577 & ~n588;
  assign n616 = n574 & ~n615;
  assign n617 = n577 & n588;
  assign n618 = ~n616 & ~n617;
  assign n619 = ~n592 & n611;
  assign n620 = n618 & n619;
  assign n621 = n574 & n617;
  assign n622 = ~n621 & n612;
  assign n623 = ~n574 & n615;
  assign n624 = n622 & ~n623;
  assign n625 = ~n620 & ~n624;
  assign n626 = n592 & ~n611;
  assign n627 = ~n618 & n626;
  assign n628 = n625 & ~n627;
  assign n629 = ~n580 & n587;
  assign n630 = n583 & ~n586;
  assign n631 = ~n629 & ~n630;
  assign n632 = ~n602 ^ pi15;
  assign n633 = ~n632 & n599;
  assign n634 = ~n598 & ~n633;
  assign n635 = n632 & ~n599;
  assign n636 = ~n635 & pi01;
  assign n637 = ~n634 & n636;
  assign n638 = n602 & ~pi01;
  assign n639 = n598 & n638;
  assign n640 = ~n637 & ~n639;
  assign n641 = n607 & ~n608;
  assign n642 = ~n605 & ~n606;
  assign n643 = ~n641 & ~n642;
  assign n644 = n584 & ~n585;
  assign n645 = ~n410 & ~n451;
  assign n646 = ~n644 & ~n645;
  assign n647 = ~n643 ^ ~n646;
  assign n648 = pi01 & pi16;
  assign n649 = ~n648 ^ ~pi09;
  assign n650 = ~n647 ^ n649;
  assign n651 = ~n640 ^ ~n650;
  assign n652 = ~n631 ^ ~n651;
  assign n653 = n595 & n610;
  assign n654 = n604 & ~n609;
  assign n655 = ~n653 & ~n654;
  assign n656 = ~n652 ^ ~n655;
  assign n657 = pi09 & pi15;
  assign n658 = n285 & n657;
  assign n659 = pi00 & pi17;
  assign n660 = pi05 & pi12;
  assign n661 = ~n659 ^ ~n660;
  assign n662 = ~n658 ^ ~n661;
  assign n663 = pi06 & pi11;
  assign n664 = pi04 & pi13;
  assign n665 = ~n663 ^ ~n664;
  assign n666 = pi02 & pi15;
  assign n667 = ~n665 ^ n666;
  assign n668 = ~n662 ^ n667;
  assign n669 = pi08 & pi09;
  assign n670 = pi07 & pi10;
  assign n671 = ~n669 ^ ~n670;
  assign n672 = pi03 & pi14;
  assign n673 = ~n671 ^ n672;
  assign n674 = ~n668 ^ n673;
  assign n675 = ~n656 ^ n674;
  assign po018 = ~n628 ^ ~n675;
  assign n677 = ~n675 & ~n626;
  assign n678 = n618 & ~n677;
  assign n679 = n675 & n626;
  assign n680 = ~n678 & ~n679;
  assign n681 = ~n623 & ~n675;
  assign n682 = n622 & ~n681;
  assign n683 = n680 & ~n682;
  assign n684 = n656 & ~n674;
  assign n685 = n652 & n655;
  assign n686 = ~n684 & ~n685;
  assign n687 = n631 & n651;
  assign n688 = n640 & n650;
  assign n689 = ~n687 & ~n688;
  assign n690 = n647 & ~n649;
  assign n691 = ~n643 & ~n646;
  assign n692 = ~n690 & ~n691;
  assign n693 = n668 & ~n673;
  assign n694 = n662 & ~n667;
  assign n695 = ~n693 & ~n694;
  assign n696 = ~n692 ^ n695;
  assign n697 = n671 & ~n672;
  assign n698 = ~n669 & ~n670;
  assign n699 = ~n697 & ~n698;
  assign n700 = n665 & ~n666;
  assign n701 = ~n663 & ~n664;
  assign n702 = ~n700 & ~n701;
  assign n703 = ~n699 ^ ~n702;
  assign n704 = n658 & n661;
  assign n705 = pi05 & pi17;
  assign n706 = n424 & n705;
  assign n707 = ~n704 & ~n706;
  assign n708 = ~n703 ^ n707;
  assign n709 = ~n696 ^ n708;
  assign n710 = n648 & pi09;
  assign n711 = pi06 & pi12;
  assign n712 = ~n710 ^ ~n711;
  assign n713 = pi01 & pi17;
  assign n714 = ~n459 ^ n713;
  assign n715 = ~n712 ^ n714;
  assign n716 = pi07 & pi11;
  assign n717 = pi05 & pi13;
  assign n718 = ~n716 ^ ~n717;
  assign n719 = pi00 & pi18;
  assign n720 = ~n718 ^ n719;
  assign n721 = pi04 & pi14;
  assign n722 = pi03 & pi15;
  assign n723 = ~n721 ^ ~n722;
  assign n724 = pi02 & pi16;
  assign n725 = ~n723 ^ n724;
  assign n726 = ~n720 ^ ~n725;
  assign n727 = ~n715 ^ ~n726;
  assign n728 = ~n709 ^ n727;
  assign n729 = ~n689 ^ n728;
  assign n730 = ~n686 ^ n729;
  assign po019 = n683 ^ n730;
  assign n732 = n709 & ~n727;
  assign n733 = n689 & ~n732;
  assign n734 = ~n709 & n727;
  assign n735 = ~n733 & ~n734;
  assign n736 = n686 & ~n735;
  assign n737 = n689 & n734;
  assign n738 = ~n736 & ~n737;
  assign n739 = n683 & ~n738;
  assign n740 = n686 & n737;
  assign n741 = ~n689 & n732;
  assign n742 = ~n686 & n741;
  assign n743 = ~n740 & ~n742;
  assign n744 = ~n739 & n743;
  assign n745 = n686 & ~n741;
  assign n746 = ~n745 & n735;
  assign n747 = ~n683 & n746;
  assign n748 = n744 & ~n747;
  assign n749 = n696 & ~n708;
  assign n750 = ~n692 & n695;
  assign n751 = ~n749 & ~n750;
  assign n752 = n715 & n726;
  assign n753 = ~n720 & ~n725;
  assign n754 = ~n752 & ~n753;
  assign n755 = n723 & ~n724;
  assign n756 = ~n721 & ~n722;
  assign n757 = ~n755 & ~n756;
  assign n758 = pi08 & pi17;
  assign n759 = n384 & n758;
  assign n760 = ~n759 & pi10;
  assign n761 = pi01 & pi18;
  assign n762 = ~n760 ^ ~n761;
  assign n763 = ~n757 ^ ~n762;
  assign n764 = ~n754 ^ n763;
  assign n765 = n712 & ~n714;
  assign n766 = n710 & n711;
  assign n767 = ~n765 & ~n766;
  assign n768 = n718 & ~n719;
  assign n769 = ~n716 & ~n717;
  assign n770 = ~n768 & ~n769;
  assign n771 = pi09 & pi10;
  assign n772 = pi08 & pi11;
  assign n773 = ~n771 ^ ~n772;
  assign n774 = pi03 & pi16;
  assign n775 = ~n773 ^ n774;
  assign n776 = ~n770 ^ n775;
  assign n777 = ~n767 ^ n776;
  assign n778 = ~n764 ^ ~n777;
  assign n779 = n703 & ~n707;
  assign n780 = n699 & n702;
  assign n781 = ~n779 & ~n780;
  assign n782 = pi06 & pi13;
  assign n783 = pi07 & pi12;
  assign n784 = ~n782 ^ ~n783;
  assign n785 = pi05 & pi14;
  assign n786 = ~n784 ^ n785;
  assign n787 = pi04 & pi15;
  assign n788 = pi02 & pi17;
  assign n789 = ~n787 ^ ~n788;
  assign n790 = pi00 & pi19;
  assign n791 = ~n789 ^ n790;
  assign n792 = ~n786 ^ ~n791;
  assign n793 = ~n781 ^ n792;
  assign n794 = ~n778 ^ ~n793;
  assign n795 = ~n751 ^ n794;
  assign po020 = n748 ^ ~n795;
  assign n797 = n738 & n795;
  assign n798 = ~n797 & ~n742;
  assign n799 = n683 & n798;
  assign n800 = ~n740 & n795;
  assign n801 = ~n746 & ~n800;
  assign n802 = ~n799 & ~n801;
  assign n803 = ~n751 & n794;
  assign n804 = ~n778 & ~n793;
  assign n805 = ~n803 & ~n804;
  assign n806 = ~n781 & n792;
  assign n807 = ~n786 & ~n791;
  assign n808 = ~n806 & ~n807;
  assign n809 = n789 & ~n790;
  assign n810 = ~n787 & ~n788;
  assign n811 = ~n809 & ~n810;
  assign n812 = n773 & ~n774;
  assign n813 = ~n771 & ~n772;
  assign n814 = ~n812 & ~n813;
  assign n815 = ~n811 ^ ~n814;
  assign n816 = pi01 & pi19;
  assign n817 = pi09 & pi11;
  assign n818 = ~n816 ^ ~n817;
  assign n819 = ~n815 ^ ~n818;
  assign n820 = ~n808 ^ n819;
  assign n821 = n761 & pi10;
  assign n822 = pi00 & pi20;
  assign n823 = ~n821 ^ ~n822;
  assign n824 = pi07 & pi13;
  assign n825 = ~n823 ^ n824;
  assign n826 = pi08 & pi12;
  assign n827 = pi06 & pi14;
  assign n828 = ~n826 ^ ~n827;
  assign n829 = pi05 & pi15;
  assign n830 = ~n828 ^ n829;
  assign n831 = ~n825 ^ ~n830;
  assign n832 = n784 & ~n785;
  assign n833 = ~n782 & ~n783;
  assign n834 = ~n832 & ~n833;
  assign n835 = ~n831 ^ n834;
  assign n836 = ~n820 ^ ~n835;
  assign n837 = n764 & n777;
  assign n838 = ~n754 & n763;
  assign n839 = ~n837 & ~n838;
  assign n840 = ~n767 & n776;
  assign n841 = n770 & ~n775;
  assign n842 = ~n840 & ~n841;
  assign n843 = n757 & n762;
  assign n844 = n759 & ~pi18;
  assign n845 = ~n843 & ~n844;
  assign n846 = pi04 & pi16;
  assign n847 = pi03 & pi17;
  assign n848 = ~n846 ^ ~n847;
  assign n849 = pi02 & pi18;
  assign n850 = ~n848 ^ n849;
  assign n851 = ~n845 ^ ~n850;
  assign n852 = ~n842 ^ n851;
  assign n853 = ~n839 ^ n852;
  assign n854 = ~n836 ^ ~n853;
  assign n855 = ~n805 ^ n854;
  assign po021 = ~n802 ^ n855;
  assign n857 = n839 & ~n852;
  assign n858 = ~n836 & ~n857;
  assign n859 = ~n839 & n852;
  assign n860 = ~n858 & ~n859;
  assign n861 = ~n836 & n859;
  assign n862 = ~n805 & ~n861;
  assign n863 = ~n860 & ~n862;
  assign n864 = ~n802 & n863;
  assign n865 = n805 & n861;
  assign n866 = n836 & n857;
  assign n867 = ~n805 & n866;
  assign n868 = ~n865 & ~n867;
  assign n869 = ~n864 & n868;
  assign n870 = n805 & ~n866;
  assign n871 = n860 & ~n870;
  assign n872 = n802 & n871;
  assign n873 = n869 & ~n872;
  assign n874 = n820 & n835;
  assign n875 = n808 & ~n819;
  assign n876 = ~n874 & ~n875;
  assign n877 = ~n842 & n851;
  assign n878 = ~n845 & ~n850;
  assign n879 = ~n877 & ~n878;
  assign n880 = pi10 & pi11;
  assign n881 = pi09 & pi12;
  assign n882 = ~n880 ^ ~n881;
  assign n883 = pi04 & pi17;
  assign n884 = ~n882 ^ n883;
  assign n885 = pi08 & pi13;
  assign n886 = pi07 & pi14;
  assign n887 = ~n885 ^ ~n886;
  assign n888 = pi06 & pi15;
  assign n889 = ~n887 ^ n888;
  assign n890 = ~n884 ^ ~n889;
  assign n891 = pi05 & pi16;
  assign n892 = pi03 & pi18;
  assign n893 = ~n891 ^ ~n892;
  assign n894 = pi02 & pi19;
  assign n895 = ~n893 ^ n894;
  assign n896 = ~n890 ^ n895;
  assign n897 = ~n879 ^ n896;
  assign n898 = n823 & ~n824;
  assign n899 = ~n821 & ~n822;
  assign n900 = ~n898 & ~n899;
  assign n901 = n848 & ~n849;
  assign n902 = ~n846 & ~n847;
  assign n903 = ~n901 & ~n902;
  assign n904 = n828 & ~n829;
  assign n905 = ~n826 & ~n827;
  assign n906 = ~n904 & ~n905;
  assign n907 = ~n903 ^ ~n906;
  assign n908 = ~n900 ^ n907;
  assign n909 = ~n897 ^ ~n908;
  assign n910 = ~n876 ^ n909;
  assign n911 = n815 & n818;
  assign n912 = n811 & n814;
  assign n913 = ~n911 & ~n912;
  assign n914 = n816 & n817;
  assign n915 = ~n914 & pi11;
  assign n916 = pi00 & pi21;
  assign n917 = pi01 & pi20;
  assign n918 = ~n916 ^ n917;
  assign n919 = ~n915 ^ ~n918;
  assign n920 = ~n913 ^ ~n919;
  assign n921 = n831 & ~n834;
  assign n922 = n825 & n830;
  assign n923 = ~n921 & ~n922;
  assign n924 = ~n920 ^ ~n923;
  assign n925 = ~n910 ^ ~n924;
  assign po022 = n873 ^ n925;
  assign n927 = ~n805 & n836;
  assign n928 = ~n802 & ~n927;
  assign n929 = n925 & ~n857;
  assign n930 = n805 & ~n836;
  assign n931 = ~n929 & ~n930;
  assign n932 = ~n928 & n931;
  assign n933 = ~n925 & n857;
  assign n934 = ~n932 & ~n933;
  assign n935 = n925 & ~n927;
  assign n936 = ~n935 & ~n859;
  assign n937 = po021 & n936;
  assign n938 = n934 & ~n937;
  assign n939 = n910 & n924;
  assign n940 = n876 & ~n909;
  assign n941 = ~n939 & ~n940;
  assign n942 = n897 & n908;
  assign n943 = n879 & ~n896;
  assign n944 = ~n942 & ~n943;
  assign n945 = ~n900 & n907;
  assign n946 = ~n903 & ~n906;
  assign n947 = ~n945 & ~n946;
  assign n948 = n882 & ~n883;
  assign n949 = ~n880 & ~n881;
  assign n950 = ~n948 & ~n949;
  assign n951 = pi11 & pi20;
  assign n952 = ~n951 ^ ~pi21;
  assign n953 = n952 & pi01;
  assign n954 = pi10 & pi12;
  assign n955 = ~n953 ^ n954;
  assign n956 = ~n950 ^ ~n955;
  assign n957 = ~n947 ^ n956;
  assign n958 = n890 & ~n895;
  assign n959 = ~n884 & ~n889;
  assign n960 = ~n958 & ~n959;
  assign n961 = ~n957 ^ ~n960;
  assign n962 = ~n944 ^ n961;
  assign n963 = n920 & n923;
  assign n964 = ~n913 & ~n919;
  assign n965 = ~n963 & ~n964;
  assign n966 = pi07 & pi15;
  assign n967 = ~n599 ^ ~n966;
  assign n968 = pi00 & pi22;
  assign n969 = ~n967 ^ n968;
  assign n970 = pi09 & pi13;
  assign n971 = pi06 & pi16;
  assign n972 = ~n970 ^ ~n971;
  assign n973 = pi02 & pi20;
  assign n974 = ~n972 ^ n973;
  assign n975 = ~n969 ^ ~n974;
  assign n976 = pi04 & pi18;
  assign n977 = ~n705 ^ ~n976;
  assign n978 = pi03 & pi19;
  assign n979 = ~n977 ^ n978;
  assign n980 = ~n975 ^ n979;
  assign n981 = ~n965 ^ n980;
  assign n982 = n919 & n916;
  assign n983 = n914 & ~pi20;
  assign n984 = ~n982 & ~n983;
  assign n985 = n887 & ~n888;
  assign n986 = ~n885 & ~n886;
  assign n987 = ~n985 & ~n986;
  assign n988 = n893 & ~n894;
  assign n989 = ~n891 & ~n892;
  assign n990 = ~n988 & ~n989;
  assign n991 = ~n987 ^ ~n990;
  assign n992 = ~n984 ^ n991;
  assign n993 = ~n981 ^ ~n992;
  assign n994 = ~n962 ^ ~n993;
  assign n995 = ~n941 ^ n994;
  assign po023 = n938 ^ n995;
  assign n997 = ~po023 & n994;
  assign n998 = n938 & ~n941;
  assign n999 = ~n997 & ~n998;
  assign n1000 = n962 & n993;
  assign n1001 = n944 & ~n961;
  assign n1002 = ~n1000 & ~n1001;
  assign n1003 = n957 & n960;
  assign n1004 = ~n947 & n956;
  assign n1005 = ~n1003 & ~n1004;
  assign n1006 = ~n954 ^ ~pi21;
  assign n1007 = n1006 & n951;
  assign n1008 = ~n950 & ~n1007;
  assign n1009 = ~n1006 & ~n951;
  assign n1010 = ~n1009 & pi01;
  assign n1011 = ~n1008 & n1010;
  assign n1012 = n954 & ~pi01;
  assign n1013 = n950 & n1012;
  assign n1014 = ~n1011 & ~n1013;
  assign n1015 = pi06 & pi17;
  assign n1016 = pi05 & pi18;
  assign n1017 = ~n1015 ^ ~n1016;
  assign n1018 = pi03 & pi20;
  assign n1019 = ~n1017 ^ n1018;
  assign n1020 = ~n1014 ^ ~n1019;
  assign n1021 = pi11 & pi12;
  assign n1022 = pi10 & pi13;
  assign n1023 = ~n1021 ^ ~n1022;
  assign n1024 = pi04 & pi19;
  assign n1025 = ~n1023 ^ n1024;
  assign n1026 = ~n1020 ^ ~n1025;
  assign n1027 = ~n1005 ^ n1026;
  assign n1028 = n967 & ~n968;
  assign n1029 = ~n599 & ~n966;
  assign n1030 = ~n1028 & ~n1029;
  assign n1031 = pi09 & pi14;
  assign n1032 = pi08 & pi15;
  assign n1033 = ~n1031 ^ ~n1032;
  assign n1034 = pi07 & pi16;
  assign n1035 = ~n1033 ^ n1034;
  assign n1036 = ~n1030 ^ n1035;
  assign n1037 = n454 & pi10;
  assign n1038 = ~n1037 ^ pi02;
  assign n1039 = ~n1038 & pi21;
  assign n1040 = pi00 & pi23;
  assign n1041 = ~n1039 ^ n1040;
  assign n1042 = ~n1036 ^ n1041;
  assign n1043 = ~n1027 ^ n1042;
  assign n1044 = ~n984 & n991;
  assign n1045 = n987 & n990;
  assign n1046 = ~n1044 & ~n1045;
  assign n1047 = n975 & ~n979;
  assign n1048 = ~n969 & ~n974;
  assign n1049 = ~n1047 & ~n1048;
  assign n1050 = n977 & ~n978;
  assign n1051 = ~n705 & ~n976;
  assign n1052 = ~n1050 & ~n1051;
  assign n1053 = n972 & ~n973;
  assign n1054 = ~n970 & ~n971;
  assign n1055 = ~n1053 & ~n1054;
  assign n1056 = ~n1052 ^ ~n1055;
  assign n1057 = pi01 & pi22;
  assign n1058 = ~n1057 ^ ~pi12;
  assign n1059 = ~n1056 ^ ~n1058;
  assign n1060 = ~n1049 ^ n1059;
  assign n1061 = ~n1046 ^ n1060;
  assign n1062 = ~n1043 ^ n1061;
  assign n1063 = n981 & n992;
  assign n1064 = ~n965 & n980;
  assign n1065 = ~n1063 & ~n1064;
  assign n1066 = ~n1062 ^ n1065;
  assign n1067 = ~n1002 ^ n1066;
  assign po024 = ~n999 ^ n1067;
  assign n1069 = ~n1002 & ~n1065;
  assign n1070 = ~n1043 & n1061;
  assign n1071 = ~n1069 & ~n1070;
  assign n1072 = n1002 & n1065;
  assign n1073 = n1043 & ~n1061;
  assign n1074 = ~n1072 & ~n1073;
  assign n1075 = ~n1071 & n1074;
  assign n1076 = ~n999 & n1075;
  assign n1077 = n1069 & n1070;
  assign n1078 = n1072 & n1073;
  assign n1079 = ~n1077 & ~n1078;
  assign n1080 = ~n1076 & n1079;
  assign n1081 = n1071 & ~n1074;
  assign n1082 = n999 & n1081;
  assign n1083 = n1080 & ~n1082;
  assign n1084 = n1027 & ~n1042;
  assign n1085 = ~n1005 & n1026;
  assign n1086 = ~n1084 & ~n1085;
  assign n1087 = ~n1046 & n1060;
  assign n1088 = ~n1049 & n1059;
  assign n1089 = ~n1087 & ~n1088;
  assign n1090 = n1056 & n1058;
  assign n1091 = n1052 & n1055;
  assign n1092 = ~n1090 & ~n1091;
  assign n1093 = n454 & pi22;
  assign n1094 = pi01 & pi23;
  assign n1095 = pi11 & pi13;
  assign n1096 = ~n1094 ^ ~n1095;
  assign n1097 = ~n1093 ^ ~n1096;
  assign n1098 = pi00 & pi24;
  assign n1099 = ~n1097 ^ n1098;
  assign n1100 = pi07 & pi17;
  assign n1101 = pi06 & pi18;
  assign n1102 = ~n1100 ^ ~n1101;
  assign n1103 = pi02 & pi22;
  assign n1104 = ~n1102 ^ n1103;
  assign n1105 = ~n1099 ^ ~n1104;
  assign n1106 = ~n1092 ^ n1105;
  assign n1107 = ~n1089 ^ n1106;
  assign n1108 = ~n1038 & n1040;
  assign n1109 = n422 & n454;
  assign n1110 = ~n1108 & ~n1109;
  assign n1111 = ~n1110 & pi21;
  assign n1112 = pi05 & pi19;
  assign n1113 = pi04 & pi20;
  assign n1114 = ~n1112 ^ ~n1113;
  assign n1115 = pi03 & pi21;
  assign n1116 = ~n1114 ^ n1115;
  assign n1117 = pi10 & pi14;
  assign n1118 = ~n657 ^ ~n1117;
  assign n1119 = pi08 & pi16;
  assign n1120 = ~n1118 ^ n1119;
  assign n1121 = ~n1116 ^ ~n1120;
  assign n1122 = ~n1111 ^ n1121;
  assign n1123 = ~n1107 ^ n1122;
  assign n1124 = n1020 & n1025;
  assign n1125 = n1014 & n1019;
  assign n1126 = ~n1124 & ~n1125;
  assign n1127 = n1033 & ~n1034;
  assign n1128 = ~n1031 & ~n1032;
  assign n1129 = ~n1127 & ~n1128;
  assign n1130 = n1017 & ~n1018;
  assign n1131 = ~n1015 & ~n1016;
  assign n1132 = ~n1130 & ~n1131;
  assign n1133 = ~n1129 ^ ~n1132;
  assign n1134 = n1023 & ~n1024;
  assign n1135 = ~n1021 & ~n1022;
  assign n1136 = ~n1134 & ~n1135;
  assign n1137 = ~n1133 ^ ~n1136;
  assign n1138 = ~n1126 ^ ~n1137;
  assign n1139 = n1036 & ~n1041;
  assign n1140 = n1030 & ~n1035;
  assign n1141 = ~n1139 & ~n1140;
  assign n1142 = ~n1138 ^ n1141;
  assign n1143 = ~n1123 ^ ~n1142;
  assign n1144 = ~n1086 ^ n1143;
  assign po025 = ~n1083 ^ n1144;
  assign n1146 = n999 & ~n1069;
  assign n1147 = n1144 & ~n1070;
  assign n1148 = ~n1072 & ~n1147;
  assign n1149 = ~n1146 & n1148;
  assign n1150 = ~n1144 & n1070;
  assign n1151 = ~n1149 & ~n1150;
  assign n1152 = ~n1069 & n1144;
  assign n1153 = ~n1152 & ~n1073;
  assign n1154 = ~po024 & n1153;
  assign n1155 = n1151 & ~n1154;
  assign n1156 = n1138 & ~n1141;
  assign n1157 = n1126 & n1137;
  assign n1158 = ~n1156 & ~n1157;
  assign n1159 = pi10 & pi15;
  assign n1160 = pi02 & pi23;
  assign n1161 = ~n1159 ^ ~n1160;
  assign n1162 = pi00 & pi25;
  assign n1163 = ~n1161 ^ n1162;
  assign n1164 = pi06 & pi19;
  assign n1165 = pi04 & pi21;
  assign n1166 = ~n1164 ^ ~n1165;
  assign n1167 = pi03 & pi22;
  assign n1168 = ~n1166 ^ n1167;
  assign n1169 = ~n1163 ^ ~n1168;
  assign n1170 = pi09 & pi16;
  assign n1171 = ~n1170 ^ ~n758;
  assign n1172 = pi07 & pi18;
  assign n1173 = ~n1171 ^ n1172;
  assign n1174 = ~n1169 ^ n1173;
  assign n1175 = ~n1158 ^ n1174;
  assign n1176 = n1133 & n1136;
  assign n1177 = n1129 & n1132;
  assign n1178 = ~n1176 & ~n1177;
  assign n1179 = n1114 & ~n1115;
  assign n1180 = ~n1112 & ~n1113;
  assign n1181 = ~n1179 & ~n1180;
  assign n1182 = pi11 & pi23;
  assign n1183 = n1182 & pi01;
  assign n1184 = ~n1183 & pi13;
  assign n1185 = pi01 & pi24;
  assign n1186 = ~n1184 ^ n1185;
  assign n1187 = ~n1181 ^ n1186;
  assign n1188 = pi12 & pi13;
  assign n1189 = pi11 & pi14;
  assign n1190 = ~n1188 ^ ~n1189;
  assign n1191 = pi05 & pi20;
  assign n1192 = ~n1190 ^ n1191;
  assign n1193 = ~n1187 ^ n1192;
  assign n1194 = ~n1178 ^ ~n1193;
  assign n1195 = ~n1175 ^ n1194;
  assign n1196 = n1107 & ~n1122;
  assign n1197 = ~n1089 & n1106;
  assign n1198 = ~n1196 & ~n1197;
  assign n1199 = ~n1195 ^ n1198;
  assign n1200 = ~n1086 & n1143;
  assign n1201 = ~n1123 & ~n1142;
  assign n1202 = ~n1200 & ~n1201;
  assign n1203 = ~n1092 & n1105;
  assign n1204 = ~n1099 & ~n1104;
  assign n1205 = ~n1203 & ~n1204;
  assign n1206 = ~n1111 & n1121;
  assign n1207 = n1116 & n1120;
  assign n1208 = ~n1206 & ~n1207;
  assign n1209 = ~n1205 ^ n1208;
  assign n1210 = n1099 & n1096;
  assign n1211 = n1093 & n1098;
  assign n1212 = ~n1210 & ~n1211;
  assign n1213 = n1118 & ~n1119;
  assign n1214 = ~n657 & ~n1117;
  assign n1215 = ~n1213 & ~n1214;
  assign n1216 = n1102 & ~n1103;
  assign n1217 = ~n1100 & ~n1101;
  assign n1218 = ~n1216 & ~n1217;
  assign n1219 = ~n1215 ^ ~n1218;
  assign n1220 = ~n1212 ^ n1219;
  assign n1221 = ~n1209 ^ n1220;
  assign n1222 = ~n1202 ^ n1221;
  assign n1223 = ~n1199 ^ n1222;
  assign po026 = ~n1155 ^ ~n1223;
  assign n1225 = n1195 & ~n1198;
  assign n1226 = n1155 & ~n1225;
  assign n1227 = ~n1195 & n1198;
  assign n1228 = ~n1226 & ~n1227;
  assign n1229 = n1202 & ~n1221;
  assign n1230 = n1228 & n1229;
  assign n1231 = ~n1202 & n1221;
  assign n1232 = n1225 & ~n1231;
  assign n1233 = ~n1155 & n1232;
  assign n1234 = n1227 & n1231;
  assign n1235 = ~n1233 & ~n1234;
  assign n1236 = ~n1225 & n1231;
  assign n1237 = n1227 & ~n1229;
  assign n1238 = ~n1236 & ~n1237;
  assign n1239 = n1155 & ~n1238;
  assign n1240 = n1235 & ~n1239;
  assign n1241 = ~n1230 & n1240;
  assign n1242 = n1175 & ~n1194;
  assign n1243 = ~n1158 & n1174;
  assign n1244 = ~n1242 & ~n1243;
  assign n1245 = n1209 & ~n1220;
  assign n1246 = n1205 & ~n1208;
  assign n1247 = ~n1245 & ~n1246;
  assign n1248 = n1181 & pi24;
  assign n1249 = n1182 & pi13;
  assign n1250 = ~n1248 & ~n1249;
  assign n1251 = pi13 & pi24;
  assign n1252 = ~n1251 & pi01;
  assign n1253 = ~n1250 & n1252;
  assign n1254 = ~n1182 & n1185;
  assign n1255 = ~n1254 & pi13;
  assign n1256 = n1181 & n1255;
  assign n1257 = ~n1253 & ~n1256;
  assign n1258 = n1171 & ~n1172;
  assign n1259 = ~n1170 & ~n758;
  assign n1260 = ~n1258 & ~n1259;
  assign n1261 = n1161 & ~n1162;
  assign n1262 = ~n1159 & ~n1160;
  assign n1263 = ~n1261 & ~n1262;
  assign n1264 = ~n1260 ^ ~n1263;
  assign n1265 = n509 & pi24;
  assign n1266 = pi00 & pi26;
  assign n1267 = pi08 & pi18;
  assign n1268 = ~n1266 ^ ~n1267;
  assign n1269 = ~n1265 ^ ~n1268;
  assign n1270 = ~n1264 ^ n1269;
  assign n1271 = ~n1257 ^ ~n1270;
  assign n1272 = ~n1212 & n1219;
  assign n1273 = n1215 & n1218;
  assign n1274 = ~n1272 & ~n1273;
  assign n1275 = ~n1271 ^ n1274;
  assign n1276 = ~n1247 ^ ~n1275;
  assign n1277 = pi07 & pi19;
  assign n1278 = pi03 & pi23;
  assign n1279 = ~n1277 ^ ~n1278;
  assign n1280 = pi02 & pi24;
  assign n1281 = ~n1279 ^ n1280;
  assign n1282 = pi06 & pi20;
  assign n1283 = pi05 & pi21;
  assign n1284 = ~n1282 ^ ~n1283;
  assign n1285 = pi04 & pi22;
  assign n1286 = ~n1284 ^ n1285;
  assign n1287 = ~n1281 ^ ~n1286;
  assign n1288 = pi11 & pi15;
  assign n1289 = pi10 & pi16;
  assign n1290 = ~n1288 ^ ~n1289;
  assign n1291 = pi09 & pi17;
  assign n1292 = ~n1290 ^ n1291;
  assign n1293 = ~n1287 ^ n1292;
  assign n1294 = ~n1276 ^ n1293;
  assign n1295 = ~n1244 ^ ~n1294;
  assign n1296 = n1178 & n1193;
  assign n1297 = ~n1187 & n1192;
  assign n1298 = ~n1296 & ~n1297;
  assign n1299 = n1190 & ~n1191;
  assign n1300 = ~n1188 & ~n1189;
  assign n1301 = ~n1299 & ~n1300;
  assign n1302 = n1166 & ~n1167;
  assign n1303 = ~n1164 & ~n1165;
  assign n1304 = ~n1302 & ~n1303;
  assign n1305 = ~n1301 ^ ~n1304;
  assign n1306 = pi01 & pi25;
  assign n1307 = pi12 & pi14;
  assign n1308 = ~n1306 ^ ~n1307;
  assign n1309 = ~n1305 ^ ~n1308;
  assign n1310 = ~n1298 ^ ~n1309;
  assign n1311 = n1169 & ~n1173;
  assign n1312 = ~n1163 & ~n1168;
  assign n1313 = ~n1311 & ~n1312;
  assign n1314 = ~n1310 ^ ~n1313;
  assign n1315 = ~n1295 ^ n1314;
  assign po027 = ~n1241 ^ ~n1315;
  assign n1317 = n1315 & ~n1231;
  assign n1318 = ~n1228 & ~n1317;
  assign n1319 = n1315 & ~n1227;
  assign n1320 = ~n1319 & ~n1229;
  assign n1321 = po026 & n1320;
  assign n1322 = ~n1315 & n1231;
  assign n1323 = ~n1321 & ~n1322;
  assign n1324 = ~n1318 & n1323;
  assign n1325 = n1295 & ~n1314;
  assign n1326 = ~n1244 & ~n1294;
  assign n1327 = ~n1325 & ~n1326;
  assign n1328 = n1276 & ~n1293;
  assign n1329 = ~n1247 & ~n1275;
  assign n1330 = ~n1328 & ~n1329;
  assign n1331 = n1271 & ~n1274;
  assign n1332 = ~n1257 & ~n1270;
  assign n1333 = ~n1331 & ~n1332;
  assign n1334 = n1279 & ~n1280;
  assign n1335 = ~n1277 & ~n1278;
  assign n1336 = ~n1334 & ~n1335;
  assign n1337 = n1290 & ~n1291;
  assign n1338 = ~n1288 & ~n1289;
  assign n1339 = ~n1337 & ~n1338;
  assign n1340 = ~n1336 ^ ~n1339;
  assign n1341 = n1284 & ~n1285;
  assign n1342 = ~n1282 & ~n1283;
  assign n1343 = ~n1341 & ~n1342;
  assign n1344 = ~n1340 ^ n1343;
  assign n1345 = ~n1333 ^ ~n1344;
  assign n1346 = pi13 & pi14;
  assign n1347 = pi12 & pi15;
  assign n1348 = ~n1346 ^ ~n1347;
  assign n1349 = pi05 & pi22;
  assign n1350 = ~n1348 ^ n1349;
  assign n1351 = pi06 & pi21;
  assign n1352 = pi04 & pi23;
  assign n1353 = ~n1351 ^ ~n1352;
  assign n1354 = pi03 & pi24;
  assign n1355 = ~n1353 ^ n1354;
  assign n1356 = ~n1350 ^ ~n1355;
  assign n1357 = pi14 & pi25;
  assign n1358 = n454 & n1357;
  assign n1359 = ~n1358 & pi14;
  assign n1360 = pi00 & pi27;
  assign n1361 = pi01 & pi26;
  assign n1362 = ~n1360 ^ n1361;
  assign n1363 = ~n1359 ^ ~n1362;
  assign n1364 = ~n1356 ^ n1363;
  assign n1365 = ~n1345 ^ n1364;
  assign n1366 = n1310 & n1313;
  assign n1367 = ~n1298 & ~n1309;
  assign n1368 = ~n1366 & ~n1367;
  assign n1369 = n1305 & n1308;
  assign n1370 = n1301 & n1304;
  assign n1371 = ~n1369 & ~n1370;
  assign n1372 = n1264 & ~n1269;
  assign n1373 = ~n1260 & ~n1263;
  assign n1374 = ~n1372 & ~n1373;
  assign n1375 = ~n1371 ^ n1374;
  assign n1376 = n1287 & ~n1292;
  assign n1377 = ~n1281 & ~n1286;
  assign n1378 = ~n1376 & ~n1377;
  assign n1379 = ~n1375 ^ n1378;
  assign n1380 = n1265 & n1268;
  assign n1381 = pi18 & pi26;
  assign n1382 = n283 & n1381;
  assign n1383 = ~n1380 & ~n1382;
  assign n1384 = pi10 & pi17;
  assign n1385 = pi09 & pi18;
  assign n1386 = ~n1384 ^ ~n1385;
  assign n1387 = pi08 & pi19;
  assign n1388 = ~n1386 ^ n1387;
  assign n1389 = pi11 & pi16;
  assign n1390 = pi07 & pi20;
  assign n1391 = ~n1389 ^ ~n1390;
  assign n1392 = pi02 & pi25;
  assign n1393 = ~n1391 ^ n1392;
  assign n1394 = ~n1388 ^ ~n1393;
  assign n1395 = ~n1383 ^ n1394;
  assign n1396 = ~n1379 ^ ~n1395;
  assign n1397 = ~n1368 ^ n1396;
  assign n1398 = ~n1365 ^ n1397;
  assign n1399 = ~n1330 ^ n1398;
  assign n1400 = ~n1327 ^ n1399;
  assign po028 = n1324 ^ n1400;
  assign n1402 = n1327 & ~n1399;
  assign n1403 = n1324 & ~n1402;
  assign n1404 = ~n1327 & n1399;
  assign n1405 = ~n1403 & ~n1404;
  assign n1406 = ~n1365 & n1368;
  assign n1407 = ~n1330 & ~n1406;
  assign n1408 = n1365 & ~n1368;
  assign n1409 = ~n1407 & ~n1408;
  assign n1410 = ~n1379 & ~n1395;
  assign n1411 = n1409 & n1410;
  assign n1412 = ~n1330 & ~n1408;
  assign n1413 = n1330 & ~n1406;
  assign n1414 = ~n1412 & ~n1413;
  assign n1415 = ~n1414 & n1396;
  assign n1416 = ~n1411 & ~n1415;
  assign n1417 = n1379 & n1395;
  assign n1418 = ~n1409 & n1417;
  assign n1419 = n1416 & ~n1418;
  assign n1420 = n1375 & ~n1378;
  assign n1421 = ~n1371 & n1374;
  assign n1422 = ~n1420 & ~n1421;
  assign n1423 = n1340 & ~n1343;
  assign n1424 = ~n1336 & ~n1339;
  assign n1425 = ~n1423 & ~n1424;
  assign n1426 = pi09 & pi19;
  assign n1427 = pi10 & pi18;
  assign n1428 = ~n1426 ^ ~n1427;
  assign n1429 = pi02 & pi26;
  assign n1430 = ~n1428 ^ n1429;
  assign n1431 = pi12 & pi16;
  assign n1432 = pi11 & pi17;
  assign n1433 = ~n1431 ^ ~n1432;
  assign n1434 = pi00 & pi28;
  assign n1435 = ~n1433 ^ n1434;
  assign n1436 = ~n1430 ^ ~n1435;
  assign n1437 = ~n1425 ^ n1436;
  assign n1438 = ~n1422 ^ ~n1437;
  assign n1439 = n1353 & ~n1354;
  assign n1440 = ~n1351 & ~n1352;
  assign n1441 = ~n1439 & ~n1440;
  assign n1442 = n1391 & ~n1392;
  assign n1443 = ~n1389 & ~n1390;
  assign n1444 = ~n1442 & ~n1443;
  assign n1445 = ~n1441 ^ ~n1444;
  assign n1446 = n1386 & ~n1387;
  assign n1447 = ~n1384 & ~n1385;
  assign n1448 = ~n1446 & ~n1447;
  assign n1449 = ~n1445 ^ ~n1448;
  assign n1450 = ~n1438 ^ n1449;
  assign n1451 = ~n1419 ^ ~n1450;
  assign n1452 = n1345 & ~n1364;
  assign n1453 = n1333 & n1344;
  assign n1454 = ~n1452 & ~n1453;
  assign n1455 = ~n1383 & n1394;
  assign n1456 = ~n1388 & ~n1393;
  assign n1457 = ~n1455 & ~n1456;
  assign n1458 = n1348 & ~n1349;
  assign n1459 = ~n1346 & ~n1347;
  assign n1460 = ~n1458 & ~n1459;
  assign n1461 = pi14 & pi26;
  assign n1462 = ~n1461 ^ ~pi27;
  assign n1463 = n1462 & pi01;
  assign n1464 = pi13 & pi15;
  assign n1465 = ~n1463 ^ n1464;
  assign n1466 = ~n1460 ^ n1465;
  assign n1467 = ~n1457 ^ n1466;
  assign n1468 = n1356 & ~n1363;
  assign n1469 = ~n1350 & ~n1355;
  assign n1470 = ~n1468 & ~n1469;
  assign n1471 = ~n1467 ^ n1470;
  assign n1472 = n1363 & n1360;
  assign n1473 = n1358 & ~pi26;
  assign n1474 = ~n1472 & ~n1473;
  assign n1475 = pi08 & pi20;
  assign n1476 = pi04 & pi24;
  assign n1477 = ~n1475 ^ ~n1476;
  assign n1478 = pi03 & pi25;
  assign n1479 = ~n1477 ^ n1478;
  assign n1480 = pi07 & pi21;
  assign n1481 = pi06 & pi22;
  assign n1482 = ~n1480 ^ ~n1481;
  assign n1483 = pi05 & pi23;
  assign n1484 = ~n1482 ^ n1483;
  assign n1485 = ~n1479 ^ ~n1484;
  assign n1486 = ~n1474 ^ n1485;
  assign n1487 = ~n1471 ^ ~n1486;
  assign n1488 = ~n1454 ^ n1487;
  assign n1489 = ~n1451 ^ n1488;
  assign po029 = ~n1405 ^ n1489;
  assign n1491 = n1451 & ~n1488;
  assign n1492 = n1405 & ~n1491;
  assign n1493 = ~n1451 & n1488;
  assign n1494 = ~n1492 & ~n1493;
  assign n1495 = ~n1451 & n1330;
  assign n1496 = ~n1408 & ~n1450;
  assign n1497 = ~n1495 & ~n1496;
  assign n1498 = ~n1497 & n1396;
  assign n1499 = ~n1451 & n1409;
  assign n1500 = ~n1450 & n1417;
  assign n1501 = ~n1499 & ~n1500;
  assign n1502 = ~n1498 & n1501;
  assign n1503 = n1438 & ~n1449;
  assign n1504 = n1422 & n1437;
  assign n1505 = ~n1503 & ~n1504;
  assign n1506 = ~n1425 & n1436;
  assign n1507 = n1430 & n1435;
  assign n1508 = ~n1506 & ~n1507;
  assign n1509 = ~n1474 & n1485;
  assign n1510 = ~n1479 & ~n1484;
  assign n1511 = ~n1509 & ~n1510;
  assign n1512 = n1428 & ~n1429;
  assign n1513 = ~n1426 & ~n1427;
  assign n1514 = ~n1512 & ~n1513;
  assign n1515 = n1433 & ~n1434;
  assign n1516 = ~n1431 & ~n1432;
  assign n1517 = ~n1515 & ~n1516;
  assign n1518 = ~n1514 ^ ~n1517;
  assign n1519 = n1464 & pi01;
  assign n1520 = ~n1519 ^ ~pi02;
  assign n1521 = n1520 & pi27;
  assign n1522 = pi00 & pi29;
  assign n1523 = ~n1521 ^ ~n1522;
  assign n1524 = ~n1518 ^ ~n1523;
  assign n1525 = ~n1511 ^ n1524;
  assign n1526 = ~n1508 ^ ~n1525;
  assign n1527 = ~n1505 ^ ~n1526;
  assign n1528 = n1467 & ~n1470;
  assign n1529 = ~n1457 & n1466;
  assign n1530 = ~n1528 & ~n1529;
  assign n1531 = ~n1527 ^ ~n1530;
  assign n1532 = ~n1464 ^ pi27;
  assign n1533 = ~n1532 & n1461;
  assign n1534 = ~n1460 & ~n1533;
  assign n1535 = n1532 & ~n1461;
  assign n1536 = ~n1535 & pi01;
  assign n1537 = ~n1534 & n1536;
  assign n1538 = n1464 & ~pi01;
  assign n1539 = n1460 & n1538;
  assign n1540 = ~n1537 & ~n1539;
  assign n1541 = n1445 & n1448;
  assign n1542 = n1441 & n1444;
  assign n1543 = ~n1541 & ~n1542;
  assign n1544 = ~n1540 ^ ~n1543;
  assign n1545 = pi14 & pi15;
  assign n1546 = pi13 & pi16;
  assign n1547 = ~n1545 ^ ~n1546;
  assign n1548 = pi06 & pi23;
  assign n1549 = ~n1547 ^ n1548;
  assign n1550 = ~n1544 ^ ~n1549;
  assign n1551 = n1477 & ~n1478;
  assign n1552 = ~n1475 & ~n1476;
  assign n1553 = ~n1551 & ~n1552;
  assign n1554 = n1482 & ~n1483;
  assign n1555 = ~n1480 & ~n1481;
  assign n1556 = ~n1554 & ~n1555;
  assign n1557 = ~n1553 ^ ~n1556;
  assign n1558 = pi01 & pi28;
  assign n1559 = ~n1558 ^ ~pi15;
  assign n1560 = ~n1557 ^ n1559;
  assign n1561 = ~n1550 ^ ~n1560;
  assign n1562 = pi12 & pi17;
  assign n1563 = pi08 & pi21;
  assign n1564 = ~n1562 ^ ~n1563;
  assign n1565 = pi03 & pi26;
  assign n1566 = ~n1564 ^ n1565;
  assign n1567 = pi11 & pi18;
  assign n1568 = pi10 & pi19;
  assign n1569 = ~n1567 ^ ~n1568;
  assign n1570 = pi09 & pi20;
  assign n1571 = ~n1569 ^ n1570;
  assign n1572 = ~n1566 ^ ~n1571;
  assign n1573 = pi07 & pi22;
  assign n1574 = pi05 & pi24;
  assign n1575 = ~n1573 ^ ~n1574;
  assign n1576 = pi04 & pi25;
  assign n1577 = ~n1575 ^ n1576;
  assign n1578 = ~n1572 ^ n1577;
  assign n1579 = ~n1561 ^ ~n1578;
  assign n1580 = ~n1531 ^ n1579;
  assign n1581 = ~n1454 & n1487;
  assign n1582 = ~n1471 & ~n1486;
  assign n1583 = ~n1581 & ~n1582;
  assign n1584 = ~n1580 ^ ~n1583;
  assign n1585 = ~n1502 ^ n1584;
  assign po030 = ~n1494 ^ ~n1585;
  assign n1587 = ~n1502 & n1583;
  assign n1588 = ~n1587 & ~n1579;
  assign n1589 = n1502 & ~n1583;
  assign n1590 = ~n1588 & ~n1589;
  assign n1591 = ~n1590 & n1531;
  assign n1592 = n1589 & ~n1579;
  assign n1593 = ~n1591 & ~n1592;
  assign n1594 = ~n1494 & ~n1593;
  assign n1595 = n1587 & n1579;
  assign n1596 = ~n1595 & ~n1592;
  assign n1597 = ~n1596 & ~n1580;
  assign n1598 = ~n1594 & ~n1597;
  assign n1599 = ~n1595 & n1531;
  assign n1600 = n1590 & ~n1599;
  assign n1601 = n1494 & n1600;
  assign n1602 = n1598 & ~n1601;
  assign n1603 = n1527 & n1530;
  assign n1604 = ~n1505 & ~n1526;
  assign n1605 = ~n1603 & ~n1604;
  assign n1606 = n1508 & n1525;
  assign n1607 = ~n1511 & n1524;
  assign n1608 = ~n1606 & ~n1607;
  assign n1609 = n1544 & n1549;
  assign n1610 = n1540 & n1543;
  assign n1611 = ~n1609 & ~n1610;
  assign n1612 = pi08 & pi22;
  assign n1613 = pi04 & pi26;
  assign n1614 = ~n1612 ^ ~n1613;
  assign n1615 = pi03 & pi27;
  assign n1616 = ~n1614 ^ n1615;
  assign n1617 = pi12 & pi18;
  assign n1618 = pi11 & pi19;
  assign n1619 = ~n1617 ^ ~n1618;
  assign n1620 = pi10 & pi20;
  assign n1621 = ~n1619 ^ n1620;
  assign n1622 = ~n1616 ^ ~n1621;
  assign n1623 = pi07 & pi23;
  assign n1624 = pi06 & pi24;
  assign n1625 = ~n1623 ^ ~n1624;
  assign n1626 = pi05 & pi25;
  assign n1627 = ~n1625 ^ n1626;
  assign n1628 = ~n1622 ^ n1627;
  assign n1629 = ~n1611 ^ ~n1628;
  assign n1630 = ~n1608 ^ ~n1629;
  assign n1631 = ~n1605 ^ n1630;
  assign n1632 = n1561 & n1578;
  assign n1633 = ~n1550 & ~n1560;
  assign n1634 = ~n1632 & ~n1633;
  assign n1635 = n1557 & ~n1559;
  assign n1636 = ~n1553 & ~n1556;
  assign n1637 = ~n1635 & ~n1636;
  assign n1638 = n1558 & pi15;
  assign n1639 = pi00 & pi30;
  assign n1640 = ~n1638 ^ ~n1639;
  assign n1641 = pi01 & pi29;
  assign n1642 = pi14 & pi16;
  assign n1643 = ~n1641 ^ ~n1642;
  assign n1644 = ~n1640 ^ ~n1643;
  assign n1645 = ~n1637 ^ ~n1644;
  assign n1646 = n1518 & n1523;
  assign n1647 = n1514 & n1517;
  assign n1648 = ~n1646 & ~n1647;
  assign n1649 = ~n1645 ^ ~n1648;
  assign n1650 = ~n1634 ^ ~n1649;
  assign n1651 = n1575 & ~n1576;
  assign n1652 = ~n1573 & ~n1574;
  assign n1653 = ~n1651 & ~n1652;
  assign n1654 = pi13 & pi17;
  assign n1655 = pi09 & pi21;
  assign n1656 = ~n1654 ^ ~n1655;
  assign n1657 = pi02 & pi28;
  assign n1658 = ~n1656 ^ n1657;
  assign n1659 = ~n1653 ^ n1658;
  assign n1660 = n1547 & ~n1548;
  assign n1661 = ~n1545 & ~n1546;
  assign n1662 = ~n1660 & ~n1661;
  assign n1663 = ~n1659 ^ ~n1662;
  assign n1664 = ~n1522 & ~pi02;
  assign n1665 = n1519 & ~n1664;
  assign n1666 = n1522 & pi02;
  assign n1667 = ~n1665 & ~n1666;
  assign n1668 = ~n1667 & pi27;
  assign n1669 = n1564 & ~n1565;
  assign n1670 = ~n1562 & ~n1563;
  assign n1671 = ~n1669 & ~n1670;
  assign n1672 = n1569 & ~n1570;
  assign n1673 = ~n1567 & ~n1568;
  assign n1674 = ~n1672 & ~n1673;
  assign n1675 = ~n1671 ^ ~n1674;
  assign n1676 = ~n1668 ^ n1675;
  assign n1677 = ~n1663 ^ n1676;
  assign n1678 = n1572 & ~n1577;
  assign n1679 = ~n1566 & ~n1571;
  assign n1680 = ~n1678 & ~n1679;
  assign n1681 = ~n1677 ^ n1680;
  assign n1682 = ~n1650 ^ n1681;
  assign n1683 = ~n1631 ^ n1682;
  assign po031 = n1602 ^ n1683;
  assign n1685 = ~n1595 & ~n1683;
  assign n1686 = ~n1685 & ~n1592;
  assign n1687 = n1686 & ~n1531;
  assign n1688 = n1590 & n1683;
  assign n1689 = ~n1687 & ~n1688;
  assign n1690 = ~n1494 & n1689;
  assign n1691 = ~n1686 & n1531;
  assign n1692 = ~n1590 & ~n1683;
  assign n1693 = ~n1691 & ~n1692;
  assign n1694 = ~n1690 & n1693;
  assign n1695 = n1631 & ~n1682;
  assign n1696 = n1605 & ~n1630;
  assign n1697 = ~n1695 & ~n1696;
  assign n1698 = n1650 & ~n1681;
  assign n1699 = n1634 & n1649;
  assign n1700 = ~n1698 & ~n1699;
  assign n1701 = n1677 & ~n1680;
  assign n1702 = n1663 & ~n1676;
  assign n1703 = ~n1701 & ~n1702;
  assign n1704 = n1640 & n1643;
  assign n1705 = n1638 & n1639;
  assign n1706 = ~n1704 & ~n1705;
  assign n1707 = pi12 & pi19;
  assign n1708 = pi13 & pi18;
  assign n1709 = ~n1707 ^ ~n1708;
  assign n1710 = ~n1709 ^ n951;
  assign n1711 = pi10 & pi21;
  assign n1712 = pi09 & pi22;
  assign n1713 = ~n1711 ^ ~n1712;
  assign n1714 = pi00 & pi31;
  assign n1715 = ~n1713 ^ n1714;
  assign n1716 = ~n1710 ^ ~n1715;
  assign n1717 = ~n1706 ^ n1716;
  assign n1718 = pi08 & pi23;
  assign n1719 = pi07 & pi24;
  assign n1720 = ~n1718 ^ ~n1719;
  assign n1721 = pi05 & pi26;
  assign n1722 = ~n1720 ^ n1721;
  assign n1723 = pi04 & pi27;
  assign n1724 = pi03 & pi28;
  assign n1725 = ~n1723 ^ ~n1724;
  assign n1726 = pi02 & pi29;
  assign n1727 = ~n1725 ^ n1726;
  assign n1728 = ~n1722 ^ ~n1727;
  assign n1729 = pi15 & pi16;
  assign n1730 = pi14 & pi17;
  assign n1731 = ~n1729 ^ ~n1730;
  assign n1732 = pi06 & pi25;
  assign n1733 = ~n1731 ^ n1732;
  assign n1734 = ~n1728 ^ ~n1733;
  assign n1735 = ~n1717 ^ n1734;
  assign n1736 = ~n1703 ^ n1735;
  assign n1737 = ~n1700 ^ ~n1736;
  assign n1738 = n1608 & n1629;
  assign n1739 = ~n1611 & ~n1628;
  assign n1740 = ~n1738 & ~n1739;
  assign n1741 = n1645 & n1648;
  assign n1742 = ~n1637 & ~n1644;
  assign n1743 = ~n1741 & ~n1742;
  assign n1744 = n1622 & ~n1627;
  assign n1745 = ~n1616 & ~n1621;
  assign n1746 = ~n1744 & ~n1745;
  assign n1747 = ~n1743 ^ n1746;
  assign n1748 = n1614 & ~n1615;
  assign n1749 = ~n1612 & ~n1613;
  assign n1750 = ~n1748 & ~n1749;
  assign n1751 = n1656 & ~n1657;
  assign n1752 = ~n1654 & ~n1655;
  assign n1753 = ~n1751 & ~n1752;
  assign n1754 = ~n1750 ^ ~n1753;
  assign n1755 = n1619 & ~n1620;
  assign n1756 = ~n1617 & ~n1618;
  assign n1757 = ~n1755 & ~n1756;
  assign n1758 = ~n1754 ^ ~n1757;
  assign n1759 = ~n1747 ^ n1758;
  assign n1760 = n1659 & n1662;
  assign n1761 = n1653 & ~n1658;
  assign n1762 = ~n1760 & ~n1761;
  assign n1763 = n1625 & ~n1626;
  assign n1764 = ~n1623 & ~n1624;
  assign n1765 = ~n1763 & ~n1764;
  assign n1766 = pi14 & pi29;
  assign n1767 = n1766 & pi01;
  assign n1768 = ~n1767 & pi16;
  assign n1769 = pi01 & pi30;
  assign n1770 = ~n1768 ^ n1769;
  assign n1771 = ~n1765 ^ n1770;
  assign n1772 = ~n1762 ^ n1771;
  assign n1773 = ~n1668 & n1675;
  assign n1774 = ~n1671 & ~n1674;
  assign n1775 = ~n1773 & ~n1774;
  assign n1776 = ~n1772 ^ n1775;
  assign n1777 = ~n1759 ^ ~n1776;
  assign n1778 = ~n1740 ^ n1777;
  assign n1779 = ~n1737 ^ n1778;
  assign n1780 = ~n1697 ^ n1779;
  assign po032 = ~n1694 ^ ~n1780;
  assign n1782 = n1697 & ~n1779;
  assign n1783 = n1694 & ~n1782;
  assign n1784 = ~n1697 & n1779;
  assign n1785 = ~n1783 & ~n1784;
  assign n1786 = n1737 & ~n1778;
  assign n1787 = n1700 & n1736;
  assign n1788 = ~n1786 & ~n1787;
  assign n1789 = n1747 & ~n1758;
  assign n1790 = ~n1743 & n1746;
  assign n1791 = ~n1789 & ~n1790;
  assign n1792 = ~n648 & ~pi02;
  assign n1793 = ~n1792 & pi30;
  assign n1794 = n648 & pi02;
  assign n1795 = n1793 & ~n1794;
  assign n1796 = pi00 & pi32;
  assign n1797 = ~n1795 ^ ~n1796;
  assign n1798 = pi13 & pi19;
  assign n1799 = pi12 & pi20;
  assign n1800 = ~n1798 ^ ~n1799;
  assign n1801 = pi11 & pi21;
  assign n1802 = ~n1800 ^ n1801;
  assign n1803 = pi14 & pi18;
  assign n1804 = pi10 & pi22;
  assign n1805 = ~n1803 ^ ~n1804;
  assign n1806 = pi03 & pi29;
  assign n1807 = ~n1805 ^ n1806;
  assign n1808 = ~n1802 ^ ~n1807;
  assign n1809 = ~n1797 ^ ~n1808;
  assign n1810 = ~n1791 ^ ~n1809;
  assign n1811 = n1765 & pi30;
  assign n1812 = n1766 & pi16;
  assign n1813 = ~n1811 & ~n1812;
  assign n1814 = pi16 & pi30;
  assign n1815 = ~n1814 & pi01;
  assign n1816 = ~n1813 & n1815;
  assign n1817 = ~n1766 & n1769;
  assign n1818 = ~n1817 & pi16;
  assign n1819 = n1765 & n1818;
  assign n1820 = ~n1816 & ~n1819;
  assign n1821 = pi09 & pi23;
  assign n1822 = pi05 & pi27;
  assign n1823 = ~n1821 ^ ~n1822;
  assign n1824 = pi04 & pi28;
  assign n1825 = ~n1823 ^ n1824;
  assign n1826 = pi08 & pi24;
  assign n1827 = pi07 & pi25;
  assign n1828 = ~n1826 ^ ~n1827;
  assign n1829 = pi06 & pi26;
  assign n1830 = ~n1828 ^ n1829;
  assign n1831 = ~n1825 ^ ~n1830;
  assign n1832 = ~n1820 ^ n1831;
  assign n1833 = ~n1810 ^ n1832;
  assign n1834 = n1772 & ~n1775;
  assign n1835 = n1762 & ~n1771;
  assign n1836 = ~n1834 & ~n1835;
  assign n1837 = n1731 & ~n1732;
  assign n1838 = ~n1729 & ~n1730;
  assign n1839 = ~n1837 & ~n1838;
  assign n1840 = n1720 & ~n1721;
  assign n1841 = ~n1718 & ~n1719;
  assign n1842 = ~n1840 & ~n1841;
  assign n1843 = ~n1839 ^ ~n1842;
  assign n1844 = pi01 & pi31;
  assign n1845 = pi15 & pi17;
  assign n1846 = ~n1844 ^ ~n1845;
  assign n1847 = ~n1843 ^ ~n1846;
  assign n1848 = ~n1836 ^ ~n1847;
  assign n1849 = n1725 & ~n1726;
  assign n1850 = ~n1723 & ~n1724;
  assign n1851 = ~n1849 & ~n1850;
  assign n1852 = n1709 & ~n951;
  assign n1853 = ~n1707 & ~n1708;
  assign n1854 = ~n1852 & ~n1853;
  assign n1855 = ~n1851 ^ ~n1854;
  assign n1856 = n1713 & ~n1714;
  assign n1857 = ~n1711 & ~n1712;
  assign n1858 = ~n1856 & ~n1857;
  assign n1859 = ~n1855 ^ ~n1858;
  assign n1860 = ~n1848 ^ n1859;
  assign n1861 = ~n1706 & n1716;
  assign n1862 = ~n1710 & ~n1715;
  assign n1863 = ~n1861 & ~n1862;
  assign n1864 = n1728 & n1733;
  assign n1865 = n1722 & n1727;
  assign n1866 = ~n1864 & ~n1865;
  assign n1867 = ~n1863 ^ n1866;
  assign n1868 = n1754 & n1757;
  assign n1869 = n1750 & n1753;
  assign n1870 = ~n1868 & ~n1869;
  assign n1871 = ~n1867 ^ ~n1870;
  assign n1872 = ~n1860 ^ ~n1871;
  assign n1873 = ~n1703 & n1735;
  assign n1874 = n1717 & ~n1734;
  assign n1875 = ~n1873 & ~n1874;
  assign n1876 = ~n1872 ^ n1875;
  assign n1877 = ~n1833 ^ ~n1876;
  assign n1878 = ~n1740 & n1777;
  assign n1879 = n1759 & n1776;
  assign n1880 = ~n1878 & ~n1879;
  assign n1881 = ~n1877 ^ n1880;
  assign n1882 = ~n1788 ^ n1881;
  assign po033 = n1785 ^ ~n1882;
  assign n1884 = ~n1833 & n1876;
  assign n1885 = ~n1884 & ~n1880;
  assign n1886 = n1833 & ~n1876;
  assign n1887 = ~n1885 & ~n1886;
  assign n1888 = n1788 & ~n1887;
  assign n1889 = n1886 & ~n1880;
  assign n1890 = ~n1888 & ~n1889;
  assign n1891 = n1884 & n1880;
  assign n1892 = ~n1788 & n1891;
  assign n1893 = n1890 & ~n1892;
  assign n1894 = n1785 & n1893;
  assign n1895 = n1788 & ~n1891;
  assign n1896 = ~n1895 & n1887;
  assign n1897 = n1788 & n1889;
  assign n1898 = ~n1896 & ~n1897;
  assign n1899 = ~n1785 & n1898;
  assign n1900 = ~n1894 & ~n1899;
  assign n1901 = n1810 & ~n1832;
  assign n1902 = ~n1791 & ~n1809;
  assign n1903 = ~n1901 & ~n1902;
  assign n1904 = ~n1794 & ~n1796;
  assign n1905 = n1793 & ~n1904;
  assign n1906 = n1800 & ~n1801;
  assign n1907 = ~n1798 & ~n1799;
  assign n1908 = ~n1906 & ~n1907;
  assign n1909 = ~n1905 ^ ~n1908;
  assign n1910 = n1805 & ~n1806;
  assign n1911 = ~n1803 & ~n1804;
  assign n1912 = ~n1910 & ~n1911;
  assign n1913 = ~n1909 ^ n1912;
  assign n1914 = pi09 & pi24;
  assign n1915 = pi04 & pi29;
  assign n1916 = ~n1914 ^ ~n1915;
  assign n1917 = pi03 & pi30;
  assign n1918 = ~n1916 ^ n1917;
  assign n1919 = pi08 & pi25;
  assign n1920 = pi06 & pi27;
  assign n1921 = ~n1919 ^ ~n1920;
  assign n1922 = pi05 & pi28;
  assign n1923 = ~n1921 ^ n1922;
  assign n1924 = ~n1918 ^ ~n1923;
  assign n1925 = pi16 & pi17;
  assign n1926 = pi15 & pi18;
  assign n1927 = ~n1925 ^ ~n1926;
  assign n1928 = pi07 & pi26;
  assign n1929 = ~n1927 ^ n1928;
  assign n1930 = ~n1924 ^ ~n1929;
  assign n1931 = ~n1913 ^ ~n1930;
  assign n1932 = n1828 & ~n1829;
  assign n1933 = ~n1826 & ~n1827;
  assign n1934 = ~n1932 & ~n1933;
  assign n1935 = pi11 & pi22;
  assign n1936 = pi02 & pi31;
  assign n1937 = ~n1935 ^ ~n1936;
  assign n1938 = pi00 & pi33;
  assign n1939 = ~n1937 ^ n1938;
  assign n1940 = ~n1934 ^ n1939;
  assign n1941 = n1823 & ~n1824;
  assign n1942 = ~n1821 & ~n1822;
  assign n1943 = ~n1941 & ~n1942;
  assign n1944 = ~n1940 ^ ~n1943;
  assign n1945 = ~n1931 ^ ~n1944;
  assign n1946 = ~n1903 ^ ~n1945;
  assign n1947 = ~n1820 & n1831;
  assign n1948 = ~n1825 & ~n1830;
  assign n1949 = ~n1947 & ~n1948;
  assign n1950 = n1797 & n1808;
  assign n1951 = ~n1802 & ~n1807;
  assign n1952 = ~n1950 & ~n1951;
  assign n1953 = ~n1949 ^ ~n1952;
  assign n1954 = n1855 & n1858;
  assign n1955 = n1851 & n1854;
  assign n1956 = ~n1954 & ~n1955;
  assign n1957 = ~n1953 ^ n1956;
  assign n1958 = ~n1946 ^ ~n1957;
  assign n1959 = n1872 & ~n1875;
  assign n1960 = ~n1860 & ~n1871;
  assign n1961 = ~n1959 & ~n1960;
  assign n1962 = ~n1958 ^ n1961;
  assign n1963 = n1848 & ~n1859;
  assign n1964 = ~n1836 & ~n1847;
  assign n1965 = ~n1963 & ~n1964;
  assign n1966 = n1867 & n1870;
  assign n1967 = n1863 & ~n1866;
  assign n1968 = ~n1966 & ~n1967;
  assign n1969 = n1843 & n1846;
  assign n1970 = n1839 & n1842;
  assign n1971 = ~n1969 & ~n1970;
  assign n1972 = pi14 & pi19;
  assign n1973 = pi13 & pi20;
  assign n1974 = ~n1972 ^ ~n1973;
  assign n1975 = pi12 & pi21;
  assign n1976 = ~n1974 ^ n1975;
  assign n1977 = ~n1971 ^ ~n1976;
  assign n1978 = pi15 & pi31;
  assign n1979 = n1978 & pi01;
  assign n1980 = ~n1979 & pi17;
  assign n1981 = pi10 & pi23;
  assign n1982 = pi01 & pi32;
  assign n1983 = ~n1981 ^ n1982;
  assign n1984 = ~n1980 ^ ~n1983;
  assign n1985 = ~n1977 ^ n1984;
  assign n1986 = ~n1968 ^ ~n1985;
  assign n1987 = ~n1965 ^ ~n1986;
  assign n1988 = ~n1962 ^ ~n1987;
  assign po034 = ~n1900 ^ n1988;
  assign n1990 = n1988 & ~n1897;
  assign n1991 = ~n1990 & ~n1896;
  assign n1992 = ~n1785 & ~n1991;
  assign n1993 = n1988 & n1890;
  assign n1994 = ~n1993 & ~n1892;
  assign n1995 = ~n1992 & n1994;
  assign n1996 = n1962 & n1987;
  assign n1997 = n1958 & ~n1961;
  assign n1998 = ~n1996 & ~n1997;
  assign n1999 = n1946 & n1957;
  assign n2000 = n1903 & n1945;
  assign n2001 = ~n1999 & ~n2000;
  assign n2002 = n1965 & n1986;
  assign n2003 = n1968 & n1985;
  assign n2004 = ~n2002 & ~n2003;
  assign n2005 = n1977 & ~n1984;
  assign n2006 = ~n1971 & ~n1976;
  assign n2007 = ~n2005 & ~n2006;
  assign n2008 = pi10 & pi32;
  assign n2009 = n2008 & pi23;
  assign n2010 = pi17 & pi31;
  assign n2011 = n2010 & pi15;
  assign n2012 = ~n2009 & ~n2011;
  assign n2013 = pi17 & pi32;
  assign n2014 = ~n2013 & pi01;
  assign n2015 = ~n2012 & n2014;
  assign n2016 = ~n1978 & n1982;
  assign n2017 = pi17 & pi23;
  assign n2018 = n2017 & pi10;
  assign n2019 = ~n2016 & n2018;
  assign n2020 = ~n2015 & ~n2019;
  assign n2021 = n1974 & ~n1975;
  assign n2022 = ~n1972 & ~n1973;
  assign n2023 = ~n2021 & ~n2022;
  assign n2024 = pi12 & pi22;
  assign n2025 = ~n1182 ^ ~n2024;
  assign n2026 = pi02 & pi32;
  assign n2027 = ~n2025 ^ n2026;
  assign n2028 = ~n2023 ^ n2027;
  assign n2029 = ~n2020 ^ n2028;
  assign n2030 = pi10 & pi24;
  assign n2031 = pi09 & pi25;
  assign n2032 = ~n2030 ^ ~n2031;
  assign n2033 = pi05 & pi29;
  assign n2034 = ~n2032 ^ n2033;
  assign n2035 = pi15 & pi19;
  assign n2036 = pi14 & pi20;
  assign n2037 = ~n2035 ^ ~n2036;
  assign n2038 = pi13 & pi21;
  assign n2039 = ~n2037 ^ n2038;
  assign n2040 = ~n2034 ^ ~n2039;
  assign n2041 = pi08 & pi26;
  assign n2042 = pi07 & pi27;
  assign n2043 = ~n2041 ^ ~n2042;
  assign n2044 = pi06 & pi28;
  assign n2045 = ~n2043 ^ n2044;
  assign n2046 = ~n2040 ^ n2045;
  assign n2047 = ~n2029 ^ ~n2046;
  assign n2048 = ~n2007 ^ n2047;
  assign n2049 = n1937 & ~n1938;
  assign n2050 = ~n1935 & ~n1936;
  assign n2051 = ~n2049 & ~n2050;
  assign n2052 = n1921 & ~n1922;
  assign n2053 = ~n1919 & ~n1920;
  assign n2054 = ~n2052 & ~n2053;
  assign n2055 = ~n2051 ^ ~n2054;
  assign n2056 = n1916 & ~n1917;
  assign n2057 = ~n1914 & ~n1915;
  assign n2058 = ~n2056 & ~n2057;
  assign n2059 = ~n2055 ^ ~n2058;
  assign n2060 = n1927 & ~n1928;
  assign n2061 = ~n1925 & ~n1926;
  assign n2062 = ~n2060 & ~n2061;
  assign n2063 = ~n2013 ^ ~pi33;
  assign n2064 = n2063 & pi01;
  assign n2065 = pi16 & pi18;
  assign n2066 = ~n2064 ^ n2065;
  assign n2067 = ~n2062 ^ ~n2066;
  assign n2068 = ~n2059 ^ n2067;
  assign n2069 = n1924 & n1929;
  assign n2070 = n1918 & n1923;
  assign n2071 = ~n2069 & ~n2070;
  assign n2072 = ~n2068 ^ n2071;
  assign n2073 = ~n2048 ^ n2072;
  assign n2074 = ~n2004 ^ n2073;
  assign n2075 = n1953 & ~n1956;
  assign n2076 = ~n1949 & ~n1952;
  assign n2077 = ~n2075 & ~n2076;
  assign n2078 = n1931 & n1944;
  assign n2079 = ~n1913 & ~n1930;
  assign n2080 = ~n2078 & ~n2079;
  assign n2081 = n1909 & ~n1912;
  assign n2082 = ~n1905 & ~n1908;
  assign n2083 = ~n2081 & ~n2082;
  assign n2084 = pi04 & pi30;
  assign n2085 = pi03 & pi31;
  assign n2086 = ~n2084 ^ ~n2085;
  assign n2087 = pi00 & pi34;
  assign n2088 = ~n2086 ^ n2087;
  assign n2089 = ~n2083 ^ n2088;
  assign n2090 = n1940 & n1943;
  assign n2091 = n1934 & ~n1939;
  assign n2092 = ~n2090 & ~n2091;
  assign n2093 = ~n2089 ^ n2092;
  assign n2094 = ~n2080 ^ n2093;
  assign n2095 = ~n2077 ^ ~n2094;
  assign n2096 = ~n2074 ^ ~n2095;
  assign n2097 = ~n2001 ^ n2096;
  assign n2098 = ~n1998 ^ ~n2097;
  assign po035 = n1995 ^ ~n2098;
  assign n2100 = ~n2074 & n2095;
  assign n2101 = n2001 & n2100;
  assign n2102 = ~n1998 & ~n2101;
  assign n2103 = n2074 & ~n2095;
  assign n2104 = n2001 & ~n2103;
  assign n2105 = ~n2104 & ~n2100;
  assign n2106 = ~n2102 & ~n2105;
  assign n2107 = n1995 & n2106;
  assign n2108 = n1998 & n2101;
  assign n2109 = ~n2107 & ~n2108;
  assign n2110 = ~n2001 & n2103;
  assign n2111 = n1998 & ~n2110;
  assign n2112 = ~n2111 & n2105;
  assign n2113 = ~n1995 & n2112;
  assign n2114 = ~n1998 & n2110;
  assign n2115 = ~n2113 & ~n2114;
  assign n2116 = n2109 & n2115;
  assign n2117 = ~n2004 & n2073;
  assign n2118 = n2048 & ~n2072;
  assign n2119 = ~n2117 & ~n2118;
  assign n2120 = n2077 & n2094;
  assign n2121 = n2080 & ~n2093;
  assign n2122 = ~n2120 & ~n2121;
  assign n2123 = n2089 & ~n2092;
  assign n2124 = n2083 & ~n2088;
  assign n2125 = ~n2123 & ~n2124;
  assign n2126 = n761 & pi16;
  assign n2127 = ~n2126 ^ pi02;
  assign n2128 = ~n2127 & pi33;
  assign n2129 = pi00 & pi35;
  assign n2130 = ~n2128 ^ ~n2129;
  assign n2131 = pi12 & pi23;
  assign n2132 = pi11 & pi24;
  assign n2133 = ~n2131 ^ ~n2132;
  assign n2134 = pi03 & pi32;
  assign n2135 = ~n2133 ^ n2134;
  assign n2136 = pi15 & pi20;
  assign n2137 = pi14 & pi21;
  assign n2138 = ~n2136 ^ ~n2137;
  assign n2139 = pi13 & pi22;
  assign n2140 = ~n2138 ^ n2139;
  assign n2141 = ~n2135 ^ ~n2140;
  assign n2142 = ~n2130 ^ n2141;
  assign n2143 = pi17 & pi18;
  assign n2144 = pi16 & pi19;
  assign n2145 = ~n2143 ^ ~n2144;
  assign n2146 = pi07 & pi28;
  assign n2147 = ~n2145 ^ n2146;
  assign n2148 = pi08 & pi27;
  assign n2149 = pi06 & pi29;
  assign n2150 = ~n2148 ^ ~n2149;
  assign n2151 = pi05 & pi30;
  assign n2152 = ~n2150 ^ n2151;
  assign n2153 = ~n2147 ^ ~n2152;
  assign n2154 = pi10 & pi25;
  assign n2155 = pi09 & pi26;
  assign n2156 = ~n2154 ^ ~n2155;
  assign n2157 = pi04 & pi31;
  assign n2158 = ~n2156 ^ n2157;
  assign n2159 = ~n2153 ^ ~n2158;
  assign n2160 = ~n2142 ^ ~n2159;
  assign n2161 = ~n2125 ^ ~n2160;
  assign n2162 = n2040 & ~n2045;
  assign n2163 = ~n2034 & ~n2039;
  assign n2164 = ~n2162 & ~n2163;
  assign n2165 = n2043 & ~n2044;
  assign n2166 = ~n2041 & ~n2042;
  assign n2167 = ~n2165 & ~n2166;
  assign n2168 = n2032 & ~n2033;
  assign n2169 = ~n2030 & ~n2031;
  assign n2170 = ~n2168 & ~n2169;
  assign n2171 = ~n2167 ^ ~n2170;
  assign n2172 = pi01 & pi34;
  assign n2173 = ~n2172 ^ ~pi18;
  assign n2174 = ~n2171 ^ ~n2173;
  assign n2175 = ~n2164 ^ n2174;
  assign n2176 = n2025 & ~n2026;
  assign n2177 = ~n1182 & ~n2024;
  assign n2178 = ~n2176 & ~n2177;
  assign n2179 = n2086 & ~n2087;
  assign n2180 = ~n2084 & ~n2085;
  assign n2181 = ~n2179 & ~n2180;
  assign n2182 = ~n2178 ^ ~n2181;
  assign n2183 = n2037 & ~n2038;
  assign n2184 = ~n2035 & ~n2036;
  assign n2185 = ~n2183 & ~n2184;
  assign n2186 = ~n2182 ^ ~n2185;
  assign n2187 = ~n2175 ^ ~n2186;
  assign n2188 = ~n2161 ^ n2187;
  assign n2189 = ~n2122 ^ n2188;
  assign n2190 = ~n2007 & n2047;
  assign n2191 = n2029 & n2046;
  assign n2192 = ~n2190 & ~n2191;
  assign n2193 = n2068 & ~n2071;
  assign n2194 = ~n2059 & n2067;
  assign n2195 = ~n2193 & ~n2194;
  assign n2196 = ~n2065 ^ pi33;
  assign n2197 = ~n2196 & n2013;
  assign n2198 = ~n2062 & ~n2197;
  assign n2199 = n2196 & ~n2013;
  assign n2200 = ~n2199 & pi01;
  assign n2201 = ~n2198 & n2200;
  assign n2202 = n2065 & ~pi01;
  assign n2203 = n2062 & n2202;
  assign n2204 = ~n2201 & ~n2203;
  assign n2205 = n2055 & n2058;
  assign n2206 = n2051 & n2054;
  assign n2207 = ~n2205 & ~n2206;
  assign n2208 = ~n2204 ^ ~n2207;
  assign n2209 = ~n2020 & n2028;
  assign n2210 = n2023 & ~n2027;
  assign n2211 = ~n2209 & ~n2210;
  assign n2212 = ~n2208 ^ n2211;
  assign n2213 = ~n2195 ^ ~n2212;
  assign n2214 = ~n2192 ^ n2213;
  assign n2215 = ~n2189 ^ ~n2214;
  assign n2216 = ~n2119 ^ n2215;
  assign po036 = ~n2116 ^ n2216;
  assign n2218 = ~n2108 & ~n2216;
  assign n2219 = ~n2112 & ~n2218;
  assign n2220 = ~n1995 & ~n2219;
  assign n2221 = ~n2106 & ~n2216;
  assign n2222 = ~n2221 & ~n2114;
  assign n2223 = ~n2220 & n2222;
  assign n2224 = n2216 & n2214;
  assign n2225 = ~n2119 & ~n2189;
  assign n2226 = ~n2224 & ~n2225;
  assign n2227 = ~n2122 & n2188;
  assign n2228 = n2161 & ~n2187;
  assign n2229 = ~n2227 & ~n2228;
  assign n2230 = ~n2192 & n2213;
  assign n2231 = n2195 & n2212;
  assign n2232 = ~n2230 & ~n2231;
  assign n2233 = n2208 & ~n2211;
  assign n2234 = ~n2204 & ~n2207;
  assign n2235 = ~n2233 & ~n2234;
  assign n2236 = pi16 & pi20;
  assign n2237 = pi15 & pi21;
  assign n2238 = ~n2236 ^ ~n2237;
  assign n2239 = pi14 & pi22;
  assign n2240 = ~n2238 ^ n2239;
  assign n2241 = pi11 & pi25;
  assign n2242 = pi04 & pi32;
  assign n2243 = ~n2241 ^ ~n2242;
  assign n2244 = pi03 & pi33;
  assign n2245 = ~n2243 ^ n2244;
  assign n2246 = ~n2240 ^ ~n2245;
  assign n2247 = n761 & pi34;
  assign n2248 = pi01 & pi35;
  assign n2249 = pi17 & pi19;
  assign n2250 = ~n2248 ^ ~n2249;
  assign n2251 = ~n2247 ^ ~n2250;
  assign n2252 = pi00 & pi36;
  assign n2253 = ~n2251 ^ n2252;
  assign n2254 = ~n2246 ^ ~n2253;
  assign n2255 = ~n2235 ^ ~n2254;
  assign n2256 = pi13 & pi23;
  assign n2257 = pi12 & pi24;
  assign n2258 = ~n2256 ^ ~n2257;
  assign n2259 = pi02 & pi34;
  assign n2260 = ~n2258 ^ n2259;
  assign n2261 = pi10 & pi26;
  assign n2262 = pi09 & pi27;
  assign n2263 = ~n2261 ^ ~n2262;
  assign n2264 = pi05 & pi31;
  assign n2265 = ~n2263 ^ n2264;
  assign n2266 = ~n2260 ^ ~n2265;
  assign n2267 = pi08 & pi28;
  assign n2268 = pi07 & pi29;
  assign n2269 = ~n2267 ^ ~n2268;
  assign n2270 = pi06 & pi30;
  assign n2271 = ~n2269 ^ n2270;
  assign n2272 = ~n2266 ^ n2271;
  assign n2273 = ~n2255 ^ n2272;
  assign n2274 = ~n2126 & ~pi02;
  assign n2275 = ~n2274 & n2129;
  assign n2276 = n724 & n761;
  assign n2277 = ~n2275 & ~n2276;
  assign n2278 = ~n2277 & pi33;
  assign n2279 = n2133 & ~n2134;
  assign n2280 = ~n2131 & ~n2132;
  assign n2281 = ~n2279 & ~n2280;
  assign n2282 = n2138 & ~n2139;
  assign n2283 = ~n2136 & ~n2137;
  assign n2284 = ~n2282 & ~n2283;
  assign n2285 = ~n2281 ^ ~n2284;
  assign n2286 = ~n2278 ^ n2285;
  assign n2287 = n2153 & n2158;
  assign n2288 = n2147 & n2152;
  assign n2289 = ~n2287 & ~n2288;
  assign n2290 = n2150 & ~n2151;
  assign n2291 = ~n2148 & ~n2149;
  assign n2292 = ~n2290 & ~n2291;
  assign n2293 = n2156 & ~n2157;
  assign n2294 = ~n2154 & ~n2155;
  assign n2295 = ~n2293 & ~n2294;
  assign n2296 = ~n2292 ^ ~n2295;
  assign n2297 = n2145 & ~n2146;
  assign n2298 = ~n2143 & ~n2144;
  assign n2299 = ~n2297 & ~n2298;
  assign n2300 = ~n2296 ^ n2299;
  assign n2301 = ~n2289 ^ n2300;
  assign n2302 = ~n2286 ^ ~n2301;
  assign n2303 = ~n2273 ^ ~n2302;
  assign n2304 = ~n2232 ^ n2303;
  assign n2305 = n2125 & n2160;
  assign n2306 = n2142 & n2159;
  assign n2307 = ~n2305 & ~n2306;
  assign n2308 = n2175 & n2186;
  assign n2309 = ~n2164 & n2174;
  assign n2310 = ~n2308 & ~n2309;
  assign n2311 = n2171 & n2173;
  assign n2312 = n2167 & n2170;
  assign n2313 = ~n2311 & ~n2312;
  assign n2314 = n2182 & n2185;
  assign n2315 = n2178 & n2181;
  assign n2316 = ~n2314 & ~n2315;
  assign n2317 = ~n2313 ^ ~n2316;
  assign n2318 = ~n2130 & n2141;
  assign n2319 = n2135 & n2140;
  assign n2320 = ~n2318 & ~n2319;
  assign n2321 = ~n2317 ^ n2320;
  assign n2322 = ~n2310 ^ ~n2321;
  assign n2323 = ~n2307 ^ ~n2322;
  assign n2324 = ~n2304 ^ n2323;
  assign n2325 = ~n2229 ^ n2324;
  assign n2326 = ~n2226 ^ n2325;
  assign po037 = ~n2223 ^ n2326;
  assign n2328 = n2304 & n2323;
  assign n2329 = ~n2229 & ~n2328;
  assign n2330 = ~n2304 & ~n2323;
  assign n2331 = ~n2329 & ~n2330;
  assign n2332 = n2226 & ~n2331;
  assign n2333 = ~n2229 & n2330;
  assign n2334 = ~n2332 & ~n2333;
  assign n2335 = n2223 & ~n2334;
  assign n2336 = n2229 & n2328;
  assign n2337 = ~n2226 & n2336;
  assign n2338 = ~n2335 & ~n2337;
  assign n2339 = n2226 & ~n2336;
  assign n2340 = ~n2339 & n2331;
  assign n2341 = ~n2223 & n2340;
  assign n2342 = n2226 & n2333;
  assign n2343 = ~n2341 & ~n2342;
  assign n2344 = n2338 & n2343;
  assign n2345 = ~n2232 & n2303;
  assign n2346 = ~n2273 & ~n2302;
  assign n2347 = ~n2345 & ~n2346;
  assign n2348 = n2307 & n2322;
  assign n2349 = ~n2310 & ~n2321;
  assign n2350 = ~n2348 & ~n2349;
  assign n2351 = n2253 & n2250;
  assign n2352 = n2247 & n2252;
  assign n2353 = ~n2351 & ~n2352;
  assign n2354 = n2263 & ~n2264;
  assign n2355 = ~n2261 & ~n2262;
  assign n2356 = ~n2354 & ~n2355;
  assign n2357 = pi15 & pi22;
  assign n2358 = pi14 & pi23;
  assign n2359 = ~n2357 ^ ~n2358;
  assign n2360 = ~n2359 ^ n1251;
  assign n2361 = ~n2356 ^ n2360;
  assign n2362 = ~n2353 ^ n2361;
  assign n2363 = n2246 & n2253;
  assign n2364 = n2240 & n2245;
  assign n2365 = ~n2363 & ~n2364;
  assign n2366 = n2243 & ~n2244;
  assign n2367 = ~n2241 & ~n2242;
  assign n2368 = ~n2366 & ~n2367;
  assign n2369 = n2238 & ~n2239;
  assign n2370 = ~n2236 & ~n2237;
  assign n2371 = ~n2369 & ~n2370;
  assign n2372 = ~n2368 ^ ~n2371;
  assign n2373 = n2258 & ~n2259;
  assign n2374 = ~n2256 & ~n2257;
  assign n2375 = ~n2373 & ~n2374;
  assign n2376 = ~n2372 ^ n2375;
  assign n2377 = ~n2365 ^ n2376;
  assign n2378 = ~n2362 ^ ~n2377;
  assign n2379 = ~n2350 ^ n2378;
  assign n2380 = n2317 & ~n2320;
  assign n2381 = n2313 & n2316;
  assign n2382 = ~n2380 & ~n2381;
  assign n2383 = ~n2278 & n2285;
  assign n2384 = ~n2281 & ~n2284;
  assign n2385 = ~n2383 & ~n2384;
  assign n2386 = pi18 & pi19;
  assign n2387 = pi17 & pi20;
  assign n2388 = ~n2386 ^ ~n2387;
  assign n2389 = pi08 & pi29;
  assign n2390 = ~n2388 ^ n2389;
  assign n2391 = pi11 & pi26;
  assign n2392 = pi10 & pi27;
  assign n2393 = ~n2391 ^ ~n2392;
  assign n2394 = pi05 & pi32;
  assign n2395 = ~n2393 ^ n2394;
  assign n2396 = ~n2390 ^ ~n2395;
  assign n2397 = ~n2385 ^ n2396;
  assign n2398 = pi09 & pi28;
  assign n2399 = pi07 & pi30;
  assign n2400 = ~n2398 ^ ~n2399;
  assign n2401 = pi06 & pi31;
  assign n2402 = ~n2400 ^ n2401;
  assign n2403 = pi16 & pi21;
  assign n2404 = pi03 & pi34;
  assign n2405 = ~n2403 ^ ~n2404;
  assign n2406 = pi02 & pi35;
  assign n2407 = ~n2405 ^ n2406;
  assign n2408 = ~n2402 ^ ~n2407;
  assign n2409 = pi12 & pi25;
  assign n2410 = pi04 & pi33;
  assign n2411 = ~n2409 ^ ~n2410;
  assign n2412 = pi00 & pi37;
  assign n2413 = ~n2411 ^ n2412;
  assign n2414 = ~n2408 ^ n2413;
  assign n2415 = ~n2397 ^ n2414;
  assign n2416 = ~n2382 ^ n2415;
  assign n2417 = ~n2379 ^ ~n2416;
  assign n2418 = ~n2347 ^ ~n2417;
  assign n2419 = n2255 & ~n2272;
  assign n2420 = n2235 & n2254;
  assign n2421 = ~n2419 & ~n2420;
  assign n2422 = n2286 & n2301;
  assign n2423 = ~n2289 & n2300;
  assign n2424 = ~n2422 & ~n2423;
  assign n2425 = n2296 & ~n2299;
  assign n2426 = ~n2292 & ~n2295;
  assign n2427 = ~n2425 & ~n2426;
  assign n2428 = n2266 & ~n2271;
  assign n2429 = ~n2260 & ~n2265;
  assign n2430 = ~n2428 & ~n2429;
  assign n2431 = n2269 & ~n2270;
  assign n2432 = ~n2267 & ~n2268;
  assign n2433 = ~n2431 & ~n2432;
  assign n2434 = pi17 & pi35;
  assign n2435 = n2434 & pi01;
  assign n2436 = ~n2435 & pi19;
  assign n2437 = pi01 & pi36;
  assign n2438 = ~n2436 ^ n2437;
  assign n2439 = ~n2433 ^ n2438;
  assign n2440 = ~n2430 ^ n2439;
  assign n2441 = ~n2427 ^ ~n2440;
  assign n2442 = ~n2424 ^ ~n2441;
  assign n2443 = ~n2421 ^ n2442;
  assign n2444 = ~n2418 ^ n2443;
  assign po038 = ~n2344 ^ ~n2444;
  assign n2446 = ~n2337 & ~n2444;
  assign n2447 = n2334 & ~n2446;
  assign n2448 = n2223 & ~n2447;
  assign n2449 = ~n2340 & ~n2444;
  assign n2450 = ~n2449 & ~n2342;
  assign n2451 = ~n2448 & n2450;
  assign n2452 = n2418 & ~n2443;
  assign n2453 = ~n2347 & ~n2417;
  assign n2454 = ~n2452 & ~n2453;
  assign n2455 = n2379 & n2416;
  assign n2456 = n2350 & ~n2378;
  assign n2457 = ~n2455 & ~n2456;
  assign n2458 = ~n2385 & n2396;
  assign n2459 = n2390 & n2395;
  assign n2460 = ~n2458 & ~n2459;
  assign n2461 = pi17 & pi21;
  assign n2462 = pi16 & pi22;
  assign n2463 = ~n2461 ^ ~n2462;
  assign n2464 = pi15 & pi23;
  assign n2465 = ~n2463 ^ n2464;
  assign n2466 = pi10 & pi28;
  assign n2467 = pi06 & pi32;
  assign n2468 = ~n2466 ^ ~n2467;
  assign n2469 = pi05 & pi33;
  assign n2470 = ~n2468 ^ n2469;
  assign n2471 = ~n2465 ^ ~n2470;
  assign n2472 = pi09 & pi29;
  assign n2473 = pi08 & pi30;
  assign n2474 = ~n2472 ^ ~n2473;
  assign n2475 = pi07 & pi31;
  assign n2476 = ~n2474 ^ n2475;
  assign n2477 = ~n2471 ^ n2476;
  assign n2478 = ~n2460 ^ ~n2477;
  assign n2479 = n2359 & ~n1251;
  assign n2480 = ~n2357 & ~n2358;
  assign n2481 = ~n2479 & ~n2480;
  assign n2482 = n2405 & ~n2406;
  assign n2483 = ~n2403 & ~n2404;
  assign n2484 = ~n2482 & ~n2483;
  assign n2485 = ~n2481 ^ ~n2484;
  assign n2486 = n2411 & ~n2412;
  assign n2487 = ~n2409 & ~n2410;
  assign n2488 = ~n2486 & ~n2487;
  assign n2489 = ~n2485 ^ ~n2488;
  assign n2490 = ~n2478 ^ n2489;
  assign n2491 = n2362 & n2377;
  assign n2492 = n2365 & ~n2376;
  assign n2493 = ~n2491 & ~n2492;
  assign n2494 = ~n2490 ^ ~n2493;
  assign n2495 = ~n2382 & n2415;
  assign n2496 = n2397 & ~n2414;
  assign n2497 = ~n2495 & ~n2496;
  assign n2498 = ~n2494 ^ n2497;
  assign n2499 = ~n2457 ^ n2498;
  assign n2500 = ~n2421 & n2442;
  assign n2501 = ~n2424 & ~n2441;
  assign n2502 = ~n2500 & ~n2501;
  assign n2503 = n2433 & pi36;
  assign n2504 = n2434 & pi19;
  assign n2505 = ~n2503 & ~n2504;
  assign n2506 = pi19 & pi36;
  assign n2507 = ~n2506 & pi01;
  assign n2508 = ~n2505 & n2507;
  assign n2509 = ~n2434 & n2437;
  assign n2510 = ~n2509 & pi19;
  assign n2511 = n2433 & n2510;
  assign n2512 = ~n2508 & ~n2511;
  assign n2513 = pi12 & pi26;
  assign n2514 = pi11 & pi27;
  assign n2515 = ~n2513 ^ ~n2514;
  assign n2516 = pi04 & pi34;
  assign n2517 = ~n2515 ^ n2516;
  assign n2518 = ~n2512 ^ ~n2517;
  assign n2519 = n2372 & ~n2375;
  assign n2520 = ~n2368 & ~n2371;
  assign n2521 = ~n2519 & ~n2520;
  assign n2522 = ~n2518 ^ ~n2521;
  assign n2523 = n2427 & n2440;
  assign n2524 = ~n2430 & n2439;
  assign n2525 = ~n2523 & ~n2524;
  assign n2526 = ~n816 & ~pi02;
  assign n2527 = ~n2526 & pi36;
  assign n2528 = n816 & pi02;
  assign n2529 = n2527 & ~n2528;
  assign n2530 = pi00 & pi38;
  assign n2531 = ~n2529 ^ ~n2530;
  assign n2532 = pi14 & pi24;
  assign n2533 = pi13 & pi25;
  assign n2534 = ~n2532 ^ ~n2533;
  assign n2535 = pi03 & pi35;
  assign n2536 = ~n2534 ^ n2535;
  assign n2537 = ~n2531 ^ n2536;
  assign n2538 = n2393 & ~n2394;
  assign n2539 = ~n2391 & ~n2392;
  assign n2540 = ~n2538 & ~n2539;
  assign n2541 = ~n2537 ^ n2540;
  assign n2542 = ~n2525 ^ ~n2541;
  assign n2543 = ~n2522 ^ ~n2542;
  assign n2544 = ~n2353 & n2361;
  assign n2545 = n2356 & ~n2360;
  assign n2546 = ~n2544 & ~n2545;
  assign n2547 = n2408 & ~n2413;
  assign n2548 = ~n2402 & ~n2407;
  assign n2549 = ~n2547 & ~n2548;
  assign n2550 = n2400 & ~n2401;
  assign n2551 = ~n2398 & ~n2399;
  assign n2552 = ~n2550 & ~n2551;
  assign n2553 = n2388 & ~n2389;
  assign n2554 = ~n2386 & ~n2387;
  assign n2555 = ~n2553 & ~n2554;
  assign n2556 = ~n2552 ^ ~n2555;
  assign n2557 = pi01 & pi37;
  assign n2558 = pi18 & pi20;
  assign n2559 = ~n2557 ^ n2558;
  assign n2560 = ~n2556 ^ n2559;
  assign n2561 = ~n2549 ^ n2560;
  assign n2562 = ~n2546 ^ n2561;
  assign n2563 = ~n2543 ^ ~n2562;
  assign n2564 = ~n2502 ^ ~n2563;
  assign n2565 = ~n2499 ^ n2564;
  assign n2566 = ~n2454 ^ n2565;
  assign po039 = ~n2451 ^ n2566;
  assign n2568 = n2564 & ~n2498;
  assign n2569 = ~n2451 & ~n2568;
  assign n2570 = n2454 & ~n2457;
  assign n2571 = ~n2564 & n2498;
  assign n2572 = ~n2570 & ~n2571;
  assign n2573 = ~n2454 & n2457;
  assign n2574 = ~n2572 & ~n2573;
  assign n2575 = n2569 & n2574;
  assign n2576 = ~n2573 & ~n2568;
  assign n2577 = n2572 & ~n2576;
  assign n2578 = n2451 & n2577;
  assign n2579 = n2573 & n2568;
  assign n2580 = n2570 & n2571;
  assign n2581 = ~n2579 & ~n2580;
  assign n2582 = ~n2578 & n2581;
  assign n2583 = ~n2575 & n2582;
  assign n2584 = n2502 & n2563;
  assign n2585 = n2543 & n2562;
  assign n2586 = ~n2584 & ~n2585;
  assign n2587 = n2494 & ~n2497;
  assign n2588 = n2490 & n2493;
  assign n2589 = ~n2587 & ~n2588;
  assign n2590 = n2518 & n2521;
  assign n2591 = ~n2512 & ~n2517;
  assign n2592 = ~n2590 & ~n2591;
  assign n2593 = pi19 & pi20;
  assign n2594 = pi18 & pi21;
  assign n2595 = ~n2593 ^ ~n2594;
  assign n2596 = pi08 & pi31;
  assign n2597 = ~n2595 ^ n2596;
  assign n2598 = pi17 & pi22;
  assign n2599 = pi12 & pi27;
  assign n2600 = ~n2598 ^ ~n2599;
  assign n2601 = pi04 & pi35;
  assign n2602 = ~n2600 ^ n2601;
  assign n2603 = ~n2597 ^ ~n2602;
  assign n2604 = pi11 & pi28;
  assign n2605 = pi10 & pi29;
  assign n2606 = ~n2604 ^ ~n2605;
  assign n2607 = pi05 & pi34;
  assign n2608 = ~n2606 ^ n2607;
  assign n2609 = ~n2603 ^ n2608;
  assign n2610 = ~n2592 ^ n2609;
  assign n2611 = n2468 & ~n2469;
  assign n2612 = ~n2466 & ~n2467;
  assign n2613 = ~n2611 & ~n2612;
  assign n2614 = n2474 & ~n2475;
  assign n2615 = ~n2472 & ~n2473;
  assign n2616 = ~n2614 & ~n2615;
  assign n2617 = ~n2613 ^ ~n2616;
  assign n2618 = n2515 & ~n2516;
  assign n2619 = ~n2513 & ~n2514;
  assign n2620 = ~n2618 & ~n2619;
  assign n2621 = ~n2617 ^ n2620;
  assign n2622 = ~n2610 ^ ~n2621;
  assign n2623 = ~n2589 ^ n2622;
  assign n2624 = n2478 & ~n2489;
  assign n2625 = ~n2460 & ~n2477;
  assign n2626 = ~n2624 & ~n2625;
  assign n2627 = ~n2546 & n2561;
  assign n2628 = ~n2549 & n2560;
  assign n2629 = ~n2627 & ~n2628;
  assign n2630 = pi13 & pi26;
  assign n2631 = pi03 & pi36;
  assign n2632 = ~n2630 ^ ~n2631;
  assign n2633 = pi02 & pi37;
  assign n2634 = ~n2632 ^ n2633;
  assign n2635 = pi16 & pi23;
  assign n2636 = pi15 & pi24;
  assign n2637 = ~n2635 ^ ~n2636;
  assign n2638 = ~n2637 ^ n1357;
  assign n2639 = ~n2634 ^ ~n2638;
  assign n2640 = pi09 & pi30;
  assign n2641 = pi07 & pi32;
  assign n2642 = ~n2640 ^ ~n2641;
  assign n2643 = pi06 & pi33;
  assign n2644 = ~n2642 ^ n2643;
  assign n2645 = ~n2639 ^ n2644;
  assign n2646 = ~n2629 ^ n2645;
  assign n2647 = ~n2626 ^ ~n2646;
  assign n2648 = ~n2623 ^ n2647;
  assign n2649 = ~n2586 ^ ~n2648;
  assign n2650 = n2522 & n2542;
  assign n2651 = ~n2525 & ~n2541;
  assign n2652 = ~n2650 & ~n2651;
  assign n2653 = n2537 & ~n2540;
  assign n2654 = ~n2531 & n2536;
  assign n2655 = ~n2653 & ~n2654;
  assign n2656 = ~n2528 & ~n2530;
  assign n2657 = n2527 & ~n2656;
  assign n2658 = n2463 & ~n2464;
  assign n2659 = ~n2461 & ~n2462;
  assign n2660 = ~n2658 & ~n2659;
  assign n2661 = ~n2657 ^ ~n2660;
  assign n2662 = n2534 & ~n2535;
  assign n2663 = ~n2532 & ~n2533;
  assign n2664 = ~n2662 & ~n2663;
  assign n2665 = ~n2661 ^ ~n2664;
  assign n2666 = ~n2655 ^ ~n2665;
  assign n2667 = n2471 & ~n2476;
  assign n2668 = ~n2465 & ~n2470;
  assign n2669 = ~n2667 & ~n2668;
  assign n2670 = ~n2666 ^ n2669;
  assign n2671 = n2556 & ~n2559;
  assign n2672 = n2552 & n2555;
  assign n2673 = ~n2671 & ~n2672;
  assign n2674 = pi20 & pi37;
  assign n2675 = n761 & n2674;
  assign n2676 = ~n2675 & pi20;
  assign n2677 = pi00 & pi39;
  assign n2678 = pi01 & pi38;
  assign n2679 = ~n2677 ^ n2678;
  assign n2680 = ~n2676 ^ ~n2679;
  assign n2681 = ~n2673 ^ ~n2680;
  assign n2682 = n2485 & n2488;
  assign n2683 = n2481 & n2484;
  assign n2684 = ~n2682 & ~n2683;
  assign n2685 = ~n2681 ^ ~n2684;
  assign n2686 = ~n2670 ^ n2685;
  assign n2687 = ~n2652 ^ ~n2686;
  assign n2688 = ~n2649 ^ n2687;
  assign po040 = ~n2583 ^ ~n2688;
  assign n2690 = ~n2573 & ~n2688;
  assign n2691 = ~n2690 & ~n2571;
  assign n2692 = ~n2569 & n2691;
  assign n2693 = ~n2688 & ~n2568;
  assign n2694 = ~n2570 & ~n2693;
  assign n2695 = n2451 & n2694;
  assign n2696 = ~n2574 & n2688;
  assign n2697 = ~n2695 & ~n2696;
  assign n2698 = ~n2692 & n2697;
  assign n2699 = n2649 & ~n2687;
  assign n2700 = ~n2586 & ~n2648;
  assign n2701 = ~n2699 & ~n2700;
  assign n2702 = n2623 & ~n2647;
  assign n2703 = ~n2589 & n2622;
  assign n2704 = ~n2702 & ~n2703;
  assign n2705 = n2626 & n2646;
  assign n2706 = ~n2629 & n2645;
  assign n2707 = ~n2705 & ~n2706;
  assign n2708 = n2610 & n2621;
  assign n2709 = n2592 & ~n2609;
  assign n2710 = ~n2708 & ~n2709;
  assign n2711 = n2639 & ~n2644;
  assign n2712 = ~n2634 & ~n2638;
  assign n2713 = ~n2711 & ~n2712;
  assign n2714 = n2603 & ~n2608;
  assign n2715 = ~n2597 & ~n2602;
  assign n2716 = ~n2714 & ~n2715;
  assign n2717 = ~n2713 ^ ~n2716;
  assign n2718 = n2632 & ~n2633;
  assign n2719 = ~n2630 & ~n2631;
  assign n2720 = ~n2718 & ~n2719;
  assign n2721 = n2606 & ~n2607;
  assign n2722 = ~n2604 & ~n2605;
  assign n2723 = ~n2721 & ~n2722;
  assign n2724 = ~n2720 ^ ~n2723;
  assign n2725 = n2600 & ~n2601;
  assign n2726 = ~n2598 & ~n2599;
  assign n2727 = ~n2725 & ~n2726;
  assign n2728 = ~n2724 ^ ~n2727;
  assign n2729 = ~n2717 ^ ~n2728;
  assign n2730 = ~n2710 ^ ~n2729;
  assign n2731 = ~n2707 ^ ~n2730;
  assign n2732 = n2652 & n2686;
  assign n2733 = ~n2670 & n2685;
  assign n2734 = ~n2732 & ~n2733;
  assign n2735 = n2666 & ~n2669;
  assign n2736 = n2655 & n2665;
  assign n2737 = ~n2735 & ~n2736;
  assign n2738 = n2617 & ~n2620;
  assign n2739 = ~n2613 & ~n2616;
  assign n2740 = ~n2738 & ~n2739;
  assign n2741 = n2595 & ~n2596;
  assign n2742 = ~n2593 & ~n2594;
  assign n2743 = ~n2741 & ~n2742;
  assign n2744 = pi20 & pi38;
  assign n2745 = ~n2744 ^ ~pi39;
  assign n2746 = n2745 & pi01;
  assign n2747 = pi19 & pi21;
  assign n2748 = ~n2746 ^ n2747;
  assign n2749 = ~n2743 ^ ~n2748;
  assign n2750 = ~n2740 ^ n2749;
  assign n2751 = n2661 & n2664;
  assign n2752 = n2657 & n2660;
  assign n2753 = ~n2751 & ~n2752;
  assign n2754 = ~n2750 ^ n2753;
  assign n2755 = ~n2737 ^ n2754;
  assign n2756 = pi11 & pi29;
  assign n2757 = pi10 & pi30;
  assign n2758 = ~n2756 ^ ~n2757;
  assign n2759 = pi06 & pi34;
  assign n2760 = ~n2758 ^ n2759;
  assign n2761 = pi13 & pi27;
  assign n2762 = ~n1461 ^ ~n2761;
  assign n2763 = pi03 & pi37;
  assign n2764 = ~n2762 ^ n2763;
  assign n2765 = ~n2760 ^ ~n2764;
  assign n2766 = pi16 & pi24;
  assign n2767 = ~n2017 ^ ~n2766;
  assign n2768 = pi15 & pi25;
  assign n2769 = ~n2767 ^ n2768;
  assign n2770 = ~n2765 ^ n2769;
  assign n2771 = ~n2755 ^ ~n2770;
  assign n2772 = n2681 & n2684;
  assign n2773 = n2673 & n2680;
  assign n2774 = ~n2772 & ~n2773;
  assign n2775 = pi09 & pi31;
  assign n2776 = pi08 & pi32;
  assign n2777 = ~n2775 ^ ~n2776;
  assign n2778 = pi07 & pi33;
  assign n2779 = ~n2777 ^ n2778;
  assign n2780 = pi12 & pi28;
  assign n2781 = pi05 & pi35;
  assign n2782 = ~n2780 ^ ~n2781;
  assign n2783 = pi04 & pi36;
  assign n2784 = ~n2782 ^ n2783;
  assign n2785 = ~n2779 ^ ~n2784;
  assign n2786 = pi18 & pi22;
  assign n2787 = pi02 & pi38;
  assign n2788 = ~n2786 ^ ~n2787;
  assign n2789 = pi00 & pi40;
  assign n2790 = ~n2788 ^ n2789;
  assign n2791 = ~n2785 ^ n2790;
  assign n2792 = ~n2774 ^ ~n2791;
  assign n2793 = n2680 & n2677;
  assign n2794 = n2675 & ~pi38;
  assign n2795 = ~n2793 & ~n2794;
  assign n2796 = n2642 & ~n2643;
  assign n2797 = ~n2640 & ~n2641;
  assign n2798 = ~n2796 & ~n2797;
  assign n2799 = n2637 & ~n1357;
  assign n2800 = ~n2635 & ~n2636;
  assign n2801 = ~n2799 & ~n2800;
  assign n2802 = ~n2798 ^ ~n2801;
  assign n2803 = ~n2795 ^ ~n2802;
  assign n2804 = ~n2792 ^ n2803;
  assign n2805 = ~n2771 ^ ~n2804;
  assign n2806 = ~n2734 ^ n2805;
  assign n2807 = ~n2731 ^ n2806;
  assign n2808 = ~n2704 ^ n2807;
  assign n2809 = ~n2701 ^ n2808;
  assign po041 = ~n2698 ^ n2809;
  assign n2811 = ~n2698 & ~n2701;
  assign n2812 = ~n2731 & ~n2806;
  assign n2813 = n2811 & n2812;
  assign n2814 = n2731 & n2806;
  assign n2815 = n2701 & n2814;
  assign n2816 = ~n2813 & ~n2815;
  assign n2817 = ~n2816 & ~n2704;
  assign n2818 = ~n2811 & ~n2812;
  assign n2819 = n2698 & n2701;
  assign n2820 = n2704 & ~n2814;
  assign n2821 = ~n2819 & n2820;
  assign n2822 = ~n2818 & n2821;
  assign n2823 = ~n2820 & ~n2812;
  assign n2824 = n2823 & n2701;
  assign n2825 = ~n2704 & n2814;
  assign n2826 = ~n2824 & ~n2825;
  assign n2827 = n2698 & ~n2826;
  assign n2828 = ~n2822 & ~n2827;
  assign n2829 = ~n2817 & n2828;
  assign n2830 = n2707 & n2730;
  assign n2831 = ~n2710 & ~n2729;
  assign n2832 = ~n2830 & ~n2831;
  assign n2833 = n2795 & n2802;
  assign n2834 = ~n2798 & ~n2801;
  assign n2835 = ~n2833 & ~n2834;
  assign n2836 = n2724 & n2727;
  assign n2837 = n2720 & n2723;
  assign n2838 = ~n2836 & ~n2837;
  assign n2839 = ~n2835 ^ n2838;
  assign n2840 = n2765 & ~n2769;
  assign n2841 = ~n2760 & ~n2764;
  assign n2842 = ~n2840 & ~n2841;
  assign n2843 = ~n2839 ^ ~n2842;
  assign n2844 = n2717 & n2728;
  assign n2845 = ~n2713 & ~n2716;
  assign n2846 = ~n2844 & ~n2845;
  assign n2847 = ~n2843 ^ ~n2846;
  assign n2848 = n2782 & ~n2783;
  assign n2849 = ~n2780 & ~n2781;
  assign n2850 = ~n2848 & ~n2849;
  assign n2851 = pi15 & pi26;
  assign n2852 = pi13 & pi28;
  assign n2853 = ~n2851 ^ ~n2852;
  assign n2854 = pi03 & pi38;
  assign n2855 = ~n2853 ^ n2854;
  assign n2856 = ~n2850 ^ n2855;
  assign n2857 = n2747 & pi01;
  assign n2858 = ~n2857 ^ pi02;
  assign n2859 = ~n2858 & pi39;
  assign n2860 = pi00 & pi41;
  assign n2861 = ~n2859 ^ n2860;
  assign n2862 = ~n2856 ^ n2861;
  assign n2863 = ~n2847 ^ n2862;
  assign n2864 = ~n2832 ^ n2863;
  assign n2865 = n2750 & ~n2753;
  assign n2866 = n2740 & ~n2749;
  assign n2867 = ~n2865 & ~n2866;
  assign n2868 = ~n2747 ^ ~pi39;
  assign n2869 = n2868 & n2744;
  assign n2870 = ~n2743 & ~n2869;
  assign n2871 = ~n2868 & ~n2744;
  assign n2872 = ~n2871 & pi01;
  assign n2873 = ~n2870 & n2872;
  assign n2874 = n2747 & ~pi01;
  assign n2875 = n2743 & n2874;
  assign n2876 = ~n2873 & ~n2875;
  assign n2877 = pi11 & pi30;
  assign n2878 = pi06 & pi35;
  assign n2879 = ~n2877 ^ ~n2878;
  assign n2880 = pi05 & pi36;
  assign n2881 = ~n2879 ^ n2880;
  assign n2882 = ~n2876 ^ ~n2881;
  assign n2883 = pi20 & pi21;
  assign n2884 = pi19 & pi22;
  assign n2885 = ~n2883 ^ ~n2884;
  assign n2886 = pi08 & pi33;
  assign n2887 = ~n2885 ^ n2886;
  assign n2888 = ~n2882 ^ n2887;
  assign n2889 = pi18 & pi23;
  assign n2890 = pi17 & pi24;
  assign n2891 = ~n2889 ^ ~n2890;
  assign n2892 = pi16 & pi25;
  assign n2893 = ~n2891 ^ n2892;
  assign n2894 = pi10 & pi31;
  assign n2895 = pi09 & pi32;
  assign n2896 = ~n2894 ^ ~n2895;
  assign n2897 = pi07 & pi34;
  assign n2898 = ~n2896 ^ n2897;
  assign n2899 = ~n2893 ^ ~n2898;
  assign n2900 = pi14 & pi27;
  assign n2901 = pi12 & pi29;
  assign n2902 = ~n2900 ^ ~n2901;
  assign n2903 = pi04 & pi37;
  assign n2904 = ~n2902 ^ n2903;
  assign n2905 = ~n2899 ^ ~n2904;
  assign n2906 = ~n2888 ^ n2905;
  assign n2907 = ~n2867 ^ ~n2906;
  assign n2908 = ~n2864 ^ n2907;
  assign n2909 = ~n2734 & n2805;
  assign n2910 = ~n2771 & ~n2804;
  assign n2911 = ~n2909 & ~n2910;
  assign n2912 = ~n2908 ^ ~n2911;
  assign n2913 = n2755 & n2770;
  assign n2914 = ~n2737 & n2754;
  assign n2915 = ~n2913 & ~n2914;
  assign n2916 = n2792 & ~n2803;
  assign n2917 = n2774 & n2791;
  assign n2918 = ~n2916 & ~n2917;
  assign n2919 = n2785 & ~n2790;
  assign n2920 = ~n2779 & ~n2784;
  assign n2921 = ~n2919 & ~n2920;
  assign n2922 = n2758 & ~n2759;
  assign n2923 = ~n2756 & ~n2757;
  assign n2924 = ~n2922 & ~n2923;
  assign n2925 = n2777 & ~n2778;
  assign n2926 = ~n2775 & ~n2776;
  assign n2927 = ~n2925 & ~n2926;
  assign n2928 = ~n2924 ^ ~n2927;
  assign n2929 = pi01 & pi40;
  assign n2930 = ~n2929 ^ pi21;
  assign n2931 = ~n2928 ^ n2930;
  assign n2932 = ~n2921 ^ n2931;
  assign n2933 = n2788 & ~n2789;
  assign n2934 = ~n2786 & ~n2787;
  assign n2935 = ~n2933 & ~n2934;
  assign n2936 = n2762 & ~n2763;
  assign n2937 = ~n1461 & ~n2761;
  assign n2938 = ~n2936 & ~n2937;
  assign n2939 = ~n2935 ^ ~n2938;
  assign n2940 = n2767 & ~n2768;
  assign n2941 = ~n2017 & ~n2766;
  assign n2942 = ~n2940 & ~n2941;
  assign n2943 = ~n2939 ^ ~n2942;
  assign n2944 = ~n2932 ^ n2943;
  assign n2945 = ~n2918 ^ ~n2944;
  assign n2946 = ~n2915 ^ ~n2945;
  assign n2947 = ~n2912 ^ ~n2946;
  assign po042 = n2829 ^ ~n2947;
  assign n2949 = ~n2947 & ~n2825;
  assign n2950 = n2704 & n2812;
  assign n2951 = ~n2949 & ~n2950;
  assign n2952 = ~n2811 & n2951;
  assign n2953 = ~n2947 & ~n2823;
  assign n2954 = n2819 & ~n2953;
  assign n2955 = ~n2952 & ~n2954;
  assign n2956 = n2947 & n2823;
  assign n2957 = n2955 & ~n2956;
  assign n2958 = n2912 & n2946;
  assign n2959 = ~n2908 & ~n2911;
  assign n2960 = ~n2958 & ~n2959;
  assign n2961 = n2864 & ~n2907;
  assign n2962 = n2832 & ~n2863;
  assign n2963 = ~n2961 & ~n2962;
  assign n2964 = n2918 & n2944;
  assign n2965 = ~n2915 & ~n2964;
  assign n2966 = ~n2918 & ~n2944;
  assign n2967 = ~n2965 & ~n2966;
  assign n2968 = n2839 & n2842;
  assign n2969 = ~n2835 & n2838;
  assign n2970 = ~n2968 & ~n2969;
  assign n2971 = n2896 & ~n2897;
  assign n2972 = ~n2894 & ~n2895;
  assign n2973 = ~n2971 & ~n2972;
  assign n2974 = pi09 & pi33;
  assign n2975 = ~n2008 ^ ~n2974;
  assign n2976 = pi08 & pi34;
  assign n2977 = ~n2975 ^ n2976;
  assign n2978 = ~n2973 ^ n2977;
  assign n2979 = pi11 & pi31;
  assign n2980 = pi07 & pi35;
  assign n2981 = ~n2979 ^ ~n2980;
  assign n2982 = pi06 & pi36;
  assign n2983 = ~n2981 ^ n2982;
  assign n2984 = ~n2978 ^ ~n2983;
  assign n2985 = pi19 & pi23;
  assign n2986 = pi18 & pi24;
  assign n2987 = ~n2985 ^ ~n2986;
  assign n2988 = pi17 & pi25;
  assign n2989 = ~n2987 ^ n2988;
  assign n2990 = pi15 & pi27;
  assign n2991 = pi14 & pi28;
  assign n2992 = ~n2990 ^ ~n2991;
  assign n2993 = pi04 & pi38;
  assign n2994 = ~n2992 ^ n2993;
  assign n2995 = ~n2989 ^ ~n2994;
  assign n2996 = pi16 & pi26;
  assign n2997 = pi03 & pi39;
  assign n2998 = ~n2996 ^ ~n2997;
  assign n2999 = pi02 & pi40;
  assign n3000 = ~n2998 ^ n2999;
  assign n3001 = ~n2995 ^ ~n3000;
  assign n3002 = ~n2984 ^ ~n3001;
  assign n3003 = ~n2970 ^ n3002;
  assign n3004 = ~n2967 ^ ~n3003;
  assign n3005 = n2882 & ~n2887;
  assign n3006 = ~n2876 & ~n2881;
  assign n3007 = ~n3005 & ~n3006;
  assign n3008 = n2902 & ~n2903;
  assign n3009 = ~n2900 & ~n2901;
  assign n3010 = ~n3008 & ~n3009;
  assign n3011 = n2879 & ~n2880;
  assign n3012 = ~n2877 & ~n2878;
  assign n3013 = ~n3011 & ~n3012;
  assign n3014 = ~n3010 ^ ~n3013;
  assign n3015 = n2885 & ~n2886;
  assign n3016 = ~n2883 & ~n2884;
  assign n3017 = ~n3015 & ~n3016;
  assign n3018 = ~n3014 ^ ~n3017;
  assign n3019 = ~n3007 ^ n3018;
  assign n3020 = ~n2857 & ~pi02;
  assign n3021 = ~n3020 & n2860;
  assign n3022 = n2857 & pi02;
  assign n3023 = ~n3021 & ~n3022;
  assign n3024 = ~n3023 & pi39;
  assign n3025 = n2853 & ~n2854;
  assign n3026 = ~n2851 & ~n2852;
  assign n3027 = ~n3025 & ~n3026;
  assign n3028 = n2891 & ~n2892;
  assign n3029 = ~n2889 & ~n2890;
  assign n3030 = ~n3028 & ~n3029;
  assign n3031 = ~n3027 ^ ~n3030;
  assign n3032 = ~n3024 ^ n3031;
  assign n3033 = ~n3019 ^ ~n3032;
  assign n3034 = n2932 & ~n2943;
  assign n3035 = n2921 & ~n2931;
  assign n3036 = ~n3034 & ~n3035;
  assign n3037 = n2928 & ~n2930;
  assign n3038 = n2924 & n2927;
  assign n3039 = ~n3037 & ~n3038;
  assign n3040 = pi21 & pi40;
  assign n3041 = ~n3040 ^ ~pi41;
  assign n3042 = n3041 & pi01;
  assign n3043 = pi00 & pi42;
  assign n3044 = pi20 & pi22;
  assign n3045 = ~n3043 ^ ~n3044;
  assign n3046 = ~n3042 ^ n3045;
  assign n3047 = pi13 & pi29;
  assign n3048 = pi12 & pi30;
  assign n3049 = ~n3047 ^ ~n3048;
  assign n3050 = pi05 & pi37;
  assign n3051 = ~n3049 ^ n3050;
  assign n3052 = ~n3046 ^ ~n3051;
  assign n3053 = ~n3039 ^ n3052;
  assign n3054 = ~n3036 ^ ~n3053;
  assign n3055 = ~n3033 ^ n3054;
  assign n3056 = ~n3004 ^ n3055;
  assign n3057 = n2847 & ~n2862;
  assign n3058 = n2843 & n2846;
  assign n3059 = ~n3057 & ~n3058;
  assign n3060 = n2867 & n2906;
  assign n3061 = ~n2888 & n2905;
  assign n3062 = ~n3060 & ~n3061;
  assign n3063 = n2939 & n2942;
  assign n3064 = n2935 & n2938;
  assign n3065 = ~n3063 & ~n3064;
  assign n3066 = n2899 & n2904;
  assign n3067 = n2893 & n2898;
  assign n3068 = ~n3066 & ~n3067;
  assign n3069 = ~n3065 ^ n3068;
  assign n3070 = n2856 & ~n2861;
  assign n3071 = n2850 & ~n2855;
  assign n3072 = ~n3070 & ~n3071;
  assign n3073 = ~n3069 ^ ~n3072;
  assign n3074 = ~n3062 ^ n3073;
  assign n3075 = ~n3059 ^ n3074;
  assign n3076 = ~n3056 ^ ~n3075;
  assign n3077 = ~n2963 ^ ~n3076;
  assign n3078 = ~n2960 ^ n3077;
  assign po043 = ~n2957 ^ ~n3078;
  assign n3080 = ~n2960 & n2963;
  assign n3081 = n3056 & n3075;
  assign n3082 = ~n3080 & ~n3081;
  assign n3083 = n2960 & ~n2963;
  assign n3084 = ~n3056 & ~n3075;
  assign n3085 = ~n3083 & ~n3084;
  assign n3086 = ~n3082 & n3085;
  assign n3087 = ~n2957 & n3086;
  assign n3088 = n3083 & n3084;
  assign n3089 = ~n3087 & ~n3088;
  assign n3090 = n3082 & ~n3085;
  assign n3091 = n2957 & n3090;
  assign n3092 = n3080 & n3081;
  assign n3093 = ~n3091 & ~n3092;
  assign n3094 = n3089 & n3093;
  assign n3095 = n3004 & ~n3055;
  assign n3096 = n2967 & n3003;
  assign n3097 = ~n3095 & ~n3096;
  assign n3098 = n3062 & ~n3073;
  assign n3099 = ~n3059 & ~n3098;
  assign n3100 = ~n3062 & n3073;
  assign n3101 = ~n3099 & ~n3100;
  assign n3102 = n3019 & n3032;
  assign n3103 = n3007 & ~n3018;
  assign n3104 = ~n3102 & ~n3103;
  assign n3105 = ~n3039 & n3052;
  assign n3106 = ~n3046 & ~n3051;
  assign n3107 = ~n3105 & ~n3106;
  assign n3108 = n2981 & ~n2982;
  assign n3109 = ~n2979 & ~n2980;
  assign n3110 = ~n3108 & ~n3109;
  assign n3111 = n2987 & ~n2988;
  assign n3112 = ~n2985 & ~n2986;
  assign n3113 = ~n3111 & ~n3112;
  assign n3114 = ~n3110 ^ ~n3113;
  assign n3115 = n2992 & ~n2993;
  assign n3116 = ~n2990 & ~n2991;
  assign n3117 = ~n3115 & ~n3116;
  assign n3118 = ~n3114 ^ ~n3117;
  assign n3119 = n2998 & ~n2999;
  assign n3120 = ~n2996 & ~n2997;
  assign n3121 = ~n3119 & ~n3120;
  assign n3122 = n3049 & ~n3050;
  assign n3123 = ~n3047 & ~n3048;
  assign n3124 = ~n3122 & ~n3123;
  assign n3125 = ~n3121 ^ ~n3124;
  assign n3126 = ~n3040 & ~n3043;
  assign n3127 = ~n3044 ^ pi41;
  assign n3128 = ~n3126 & ~n3127;
  assign n3129 = n3040 & n3043;
  assign n3130 = ~n3129 & pi01;
  assign n3131 = ~n3128 & n3130;
  assign n3132 = n3043 & n3044;
  assign n3133 = ~n3132 & ~pi01;
  assign n3134 = ~n3131 & ~n3133;
  assign n3135 = ~n3125 ^ ~n3134;
  assign n3136 = ~n3118 ^ ~n3135;
  assign n3137 = ~n3107 ^ ~n3136;
  assign n3138 = ~n3024 & n3031;
  assign n3139 = ~n3027 & ~n3030;
  assign n3140 = ~n3138 & ~n3139;
  assign n3141 = n3014 & n3017;
  assign n3142 = n3010 & n3013;
  assign n3143 = ~n3141 & ~n3142;
  assign n3144 = pi12 & pi31;
  assign n3145 = pi11 & pi32;
  assign n3146 = ~n3144 ^ ~n3145;
  assign n3147 = pi06 & pi37;
  assign n3148 = ~n3146 ^ n3147;
  assign n3149 = ~n3143 ^ ~n3148;
  assign n3150 = ~n3140 ^ ~n3149;
  assign n3151 = ~n3137 ^ n3150;
  assign n3152 = ~n3104 ^ ~n3151;
  assign n3153 = n3069 & n3072;
  assign n3154 = n3065 & ~n3068;
  assign n3155 = ~n3153 & ~n3154;
  assign n3156 = pi21 & pi22;
  assign n3157 = pi20 & pi23;
  assign n3158 = ~n3156 ^ ~n3157;
  assign n3159 = pi09 & pi34;
  assign n3160 = ~n3158 ^ n3159;
  assign n3161 = pi13 & pi30;
  assign n3162 = pi05 & pi38;
  assign n3163 = ~n3161 ^ ~n3162;
  assign n3164 = pi02 & pi41;
  assign n3165 = ~n3163 ^ n3164;
  assign n3166 = ~n3160 ^ ~n3165;
  assign n3167 = pi10 & pi33;
  assign n3168 = pi08 & pi35;
  assign n3169 = ~n3167 ^ ~n3168;
  assign n3170 = pi07 & pi36;
  assign n3171 = ~n3169 ^ n3170;
  assign n3172 = ~n3166 ^ n3171;
  assign n3173 = ~n3155 ^ ~n3172;
  assign n3174 = pi15 & pi28;
  assign n3175 = pi16 & pi27;
  assign n3176 = ~n3174 ^ ~n3175;
  assign n3177 = ~n3176 ^ n1766;
  assign n3178 = pi19 & pi24;
  assign n3179 = pi18 & pi25;
  assign n3180 = ~n3178 ^ ~n3179;
  assign n3181 = pi17 & pi26;
  assign n3182 = ~n3180 ^ n3181;
  assign n3183 = ~n3177 ^ ~n3182;
  assign n3184 = pi04 & pi39;
  assign n3185 = pi03 & pi40;
  assign n3186 = ~n3184 ^ ~n3185;
  assign n3187 = pi00 & pi43;
  assign n3188 = ~n3186 ^ n3187;
  assign n3189 = ~n3183 ^ n3188;
  assign n3190 = ~n3173 ^ n3189;
  assign n3191 = ~n3152 ^ ~n3190;
  assign n3192 = ~n3101 ^ n3191;
  assign n3193 = n3036 & n3053;
  assign n3194 = n3033 & ~n3193;
  assign n3195 = ~n3036 & ~n3053;
  assign n3196 = ~n3194 & ~n3195;
  assign n3197 = ~n2970 & n3002;
  assign n3198 = n2984 & n3001;
  assign n3199 = ~n3197 & ~n3198;
  assign n3200 = ~n3001 & n2989;
  assign n3201 = n3000 & n2994;
  assign n3202 = ~n3200 & ~n3201;
  assign n3203 = n2975 & ~n2976;
  assign n3204 = ~n2008 & ~n2974;
  assign n3205 = ~n3203 & ~n3204;
  assign n3206 = pi01 & pi42;
  assign n3207 = ~n3205 ^ n3206;
  assign n3208 = pi20 & pi41;
  assign n3209 = n3208 & pi01;
  assign n3210 = ~n3209 & pi22;
  assign n3211 = ~n3207 ^ ~n3210;
  assign n3212 = ~n3202 ^ n3211;
  assign n3213 = n2978 & n2983;
  assign n3214 = ~n2973 & n2977;
  assign n3215 = ~n3213 & ~n3214;
  assign n3216 = ~n3212 ^ n3215;
  assign n3217 = ~n3199 ^ ~n3216;
  assign n3218 = ~n3196 ^ ~n3217;
  assign n3219 = ~n3192 ^ n3218;
  assign n3220 = ~n3097 ^ n3219;
  assign po044 = ~n3094 ^ n3220;
  assign n3222 = ~n3080 & ~n3220;
  assign n3223 = ~n3222 & ~n3084;
  assign n3224 = ~n3220 & ~n3081;
  assign n3225 = ~n3083 & ~n3224;
  assign n3226 = ~n3223 & ~n3225;
  assign n3227 = ~n2957 & ~n3226;
  assign n3228 = ~n3092 & ~n3220;
  assign n3229 = ~n3090 & ~n3228;
  assign n3230 = ~n3227 & ~n3229;
  assign n3231 = ~n3192 & n3218;
  assign n3232 = n3097 & ~n3231;
  assign n3233 = n3192 & ~n3218;
  assign n3234 = ~n3232 & ~n3233;
  assign n3235 = n3196 & ~n3216;
  assign n3236 = ~n3235 & ~n3199;
  assign n3237 = ~n3196 & n3216;
  assign n3238 = ~n3236 & ~n3237;
  assign n3239 = ~n3118 & ~n3135;
  assign n3240 = ~n3107 & ~n3239;
  assign n3241 = n3118 & n3135;
  assign n3242 = ~n3240 & ~n3241;
  assign n3243 = n3205 & ~n3206;
  assign n3244 = n3205 & n3208;
  assign n3245 = ~n3243 & ~n3244;
  assign n3246 = pi22 & pi42;
  assign n3247 = ~n3210 & ~n3246;
  assign n3248 = n3245 & ~n3247;
  assign n3249 = n3205 & n3206;
  assign n3250 = ~n3249 & ~pi22;
  assign n3251 = ~n3248 & ~n3250;
  assign n3252 = n3125 & n3134;
  assign n3253 = n3121 & n3124;
  assign n3254 = ~n3252 & ~n3253;
  assign n3255 = n3114 & n3117;
  assign n3256 = n3110 & n3113;
  assign n3257 = ~n3255 & ~n3256;
  assign n3258 = ~n3254 ^ ~n3257;
  assign n3259 = ~n3251 ^ n3258;
  assign n3260 = ~n3242 ^ n3259;
  assign n3261 = n3140 & n3149;
  assign n3262 = ~n3143 & ~n3148;
  assign n3263 = ~n3261 & ~n3262;
  assign n3264 = ~n1057 & ~pi02;
  assign n3265 = ~n3264 & pi42;
  assign n3266 = n1057 & pi02;
  assign n3267 = n3265 & ~n3266;
  assign n3268 = pi00 & pi44;
  assign n3269 = ~n3267 ^ ~n3268;
  assign n3270 = n3176 & ~n1766;
  assign n3271 = ~n3174 & ~n3175;
  assign n3272 = ~n3270 & ~n3271;
  assign n3273 = ~n3269 ^ ~n3272;
  assign n3274 = n3146 & ~n3147;
  assign n3275 = ~n3144 & ~n3145;
  assign n3276 = ~n3274 & ~n3275;
  assign n3277 = ~n3273 ^ ~n3276;
  assign n3278 = n3158 & ~n3159;
  assign n3279 = ~n3156 & ~n3157;
  assign n3280 = ~n3278 & ~n3279;
  assign n3281 = n3169 & ~n3170;
  assign n3282 = ~n3167 & ~n3168;
  assign n3283 = ~n3281 & ~n3282;
  assign n3284 = ~n3280 ^ ~n3283;
  assign n3285 = pi01 & pi43;
  assign n3286 = pi21 & pi23;
  assign n3287 = ~n3285 ^ ~n3286;
  assign n3288 = ~n3284 ^ ~n3287;
  assign n3289 = ~n3277 ^ ~n3288;
  assign n3290 = ~n3263 ^ ~n3289;
  assign n3291 = ~n3260 ^ n3290;
  assign n3292 = n3212 & ~n3215;
  assign n3293 = ~n3202 & n3211;
  assign n3294 = ~n3292 & ~n3293;
  assign n3295 = pi11 & pi33;
  assign n3296 = pi07 & pi37;
  assign n3297 = ~n3295 ^ ~n3296;
  assign n3298 = pi06 & pi38;
  assign n3299 = ~n3297 ^ n3298;
  assign n3300 = pi17 & pi27;
  assign n3301 = pi15 & pi29;
  assign n3302 = ~n3300 ^ ~n3301;
  assign n3303 = pi03 & pi41;
  assign n3304 = ~n3302 ^ n3303;
  assign n3305 = ~n3299 ^ ~n3304;
  assign n3306 = pi20 & pi24;
  assign n3307 = pi19 & pi25;
  assign n3308 = ~n3306 ^ ~n3307;
  assign n3309 = ~n3308 ^ n1381;
  assign n3310 = ~n3305 ^ n3309;
  assign n3311 = ~n3294 ^ ~n3310;
  assign n3312 = pi10 & pi34;
  assign n3313 = pi09 & pi35;
  assign n3314 = ~n3312 ^ ~n3313;
  assign n3315 = pi08 & pi36;
  assign n3316 = ~n3314 ^ n3315;
  assign n3317 = pi16 & pi28;
  assign n3318 = pi14 & pi30;
  assign n3319 = ~n3317 ^ ~n3318;
  assign n3320 = pi04 & pi40;
  assign n3321 = ~n3319 ^ n3320;
  assign n3322 = ~n3316 ^ ~n3321;
  assign n3323 = pi13 & pi31;
  assign n3324 = pi12 & pi32;
  assign n3325 = ~n3323 ^ ~n3324;
  assign n3326 = pi05 & pi39;
  assign n3327 = ~n3325 ^ n3326;
  assign n3328 = ~n3322 ^ n3327;
  assign n3329 = ~n3311 ^ n3328;
  assign n3330 = ~n3291 ^ ~n3329;
  assign n3331 = ~n3238 ^ n3330;
  assign n3332 = n3137 & ~n3150;
  assign n3333 = n3104 & ~n3332;
  assign n3334 = ~n3137 & n3150;
  assign n3335 = ~n3333 & ~n3334;
  assign n3336 = n3173 & ~n3189;
  assign n3337 = ~n3155 & ~n3172;
  assign n3338 = ~n3336 & ~n3337;
  assign n3339 = n3166 & ~n3171;
  assign n3340 = ~n3160 & ~n3165;
  assign n3341 = ~n3339 & ~n3340;
  assign n3342 = n3183 & ~n3188;
  assign n3343 = ~n3177 & ~n3182;
  assign n3344 = ~n3342 & ~n3343;
  assign n3345 = ~n3341 ^ ~n3344;
  assign n3346 = n3180 & ~n3181;
  assign n3347 = ~n3178 & ~n3179;
  assign n3348 = ~n3346 & ~n3347;
  assign n3349 = n3186 & ~n3187;
  assign n3350 = ~n3184 & ~n3185;
  assign n3351 = ~n3349 & ~n3350;
  assign n3352 = ~n3348 ^ ~n3351;
  assign n3353 = n3163 & ~n3164;
  assign n3354 = ~n3161 & ~n3162;
  assign n3355 = ~n3353 & ~n3354;
  assign n3356 = ~n3352 ^ ~n3355;
  assign n3357 = ~n3345 ^ ~n3356;
  assign n3358 = ~n3338 ^ ~n3357;
  assign n3359 = ~n3335 ^ ~n3358;
  assign n3360 = ~n3331 ^ n3359;
  assign n3361 = n3101 & ~n3190;
  assign n3362 = ~n3361 & ~n3152;
  assign n3363 = ~n3101 & n3190;
  assign n3364 = ~n3362 & ~n3363;
  assign n3365 = ~n3360 ^ n3364;
  assign n3366 = ~n3234 ^ n3365;
  assign po045 = n3230 ^ n3366;
  assign n3368 = n3364 & ~n3359;
  assign n3369 = ~n3368 & n3331;
  assign n3370 = ~n3364 & n3359;
  assign n3371 = ~n3369 & ~n3370;
  assign n3372 = ~n3371 & n3234;
  assign n3373 = n3370 & n3331;
  assign n3374 = ~n3372 & ~n3373;
  assign n3375 = ~n3230 & ~n3374;
  assign n3376 = n3368 & ~n3331;
  assign n3377 = ~n3234 & n3376;
  assign n3378 = ~n3375 & ~n3377;
  assign n3379 = n3234 & ~n3376;
  assign n3380 = ~n3379 & n3371;
  assign n3381 = n3230 & n3380;
  assign n3382 = n3234 & n3373;
  assign n3383 = ~n3381 & ~n3382;
  assign n3384 = n3378 & n3383;
  assign n3385 = n3291 & n3329;
  assign n3386 = n3238 & ~n3385;
  assign n3387 = ~n3291 & ~n3329;
  assign n3388 = ~n3386 & ~n3387;
  assign n3389 = ~n3338 & ~n3357;
  assign n3390 = ~n3335 & ~n3389;
  assign n3391 = n3338 & n3357;
  assign n3392 = ~n3390 & ~n3391;
  assign n3393 = n3277 & n3288;
  assign n3394 = n3263 & ~n3393;
  assign n3395 = ~n3277 & ~n3288;
  assign n3396 = ~n3394 & ~n3395;
  assign n3397 = n3273 & n3276;
  assign n3398 = n3269 & n3272;
  assign n3399 = ~n3397 & ~n3398;
  assign n3400 = n3284 & n3287;
  assign n3401 = n3280 & n3283;
  assign n3402 = ~n3400 & ~n3401;
  assign n3403 = ~n3399 ^ ~n3402;
  assign n3404 = n3352 & n3355;
  assign n3405 = n3348 & n3351;
  assign n3406 = ~n3404 & ~n3405;
  assign n3407 = ~n3403 ^ n3406;
  assign n3408 = n3305 & ~n3309;
  assign n3409 = ~n3299 & ~n3304;
  assign n3410 = ~n3408 & ~n3409;
  assign n3411 = n3322 & ~n3327;
  assign n3412 = ~n3316 & ~n3321;
  assign n3413 = ~n3411 & ~n3412;
  assign n3414 = ~n3410 ^ ~n3413;
  assign n3415 = n3325 & ~n3326;
  assign n3416 = ~n3323 & ~n3324;
  assign n3417 = ~n3415 & ~n3416;
  assign n3418 = n3319 & ~n3320;
  assign n3419 = ~n3317 & ~n3318;
  assign n3420 = ~n3418 & ~n3419;
  assign n3421 = ~n3417 ^ ~n3420;
  assign n3422 = n3297 & ~n3298;
  assign n3423 = ~n3295 & ~n3296;
  assign n3424 = ~n3422 & ~n3423;
  assign n3425 = ~n3421 ^ n3424;
  assign n3426 = ~n3414 ^ n3425;
  assign n3427 = ~n3407 ^ ~n3426;
  assign n3428 = ~n3396 ^ ~n3427;
  assign n3429 = n3345 & n3356;
  assign n3430 = ~n3341 & ~n3344;
  assign n3431 = ~n3429 & ~n3430;
  assign n3432 = pi22 & pi23;
  assign n3433 = pi21 & pi24;
  assign n3434 = ~n3432 ^ ~n3433;
  assign n3435 = pi10 & pi35;
  assign n3436 = ~n3434 ^ n3435;
  assign n3437 = pi09 & pi36;
  assign n3438 = pi08 & pi37;
  assign n3439 = ~n3437 ^ ~n3438;
  assign n3440 = pi07 & pi38;
  assign n3441 = ~n3439 ^ n3440;
  assign n3442 = ~n3436 ^ ~n3441;
  assign n3443 = pi04 & pi41;
  assign n3444 = pi02 & pi43;
  assign n3445 = ~n3443 ^ ~n3444;
  assign n3446 = pi00 & pi45;
  assign n3447 = ~n3445 ^ n3446;
  assign n3448 = ~n3442 ^ ~n3447;
  assign n3449 = ~n3431 ^ ~n3448;
  assign n3450 = n3314 & ~n3315;
  assign n3451 = ~n3312 & ~n3313;
  assign n3452 = ~n3450 & ~n3451;
  assign n3453 = pi20 & pi25;
  assign n3454 = pi19 & pi26;
  assign n3455 = ~n3453 ^ ~n3454;
  assign n3456 = pi18 & pi27;
  assign n3457 = ~n3455 ^ n3456;
  assign n3458 = ~n3452 ^ n3457;
  assign n3459 = pi14 & pi31;
  assign n3460 = pi13 & pi32;
  assign n3461 = ~n3459 ^ ~n3460;
  assign n3462 = pi05 & pi40;
  assign n3463 = ~n3461 ^ n3462;
  assign n3464 = ~n3458 ^ n3463;
  assign n3465 = ~n3449 ^ n3464;
  assign n3466 = ~n3428 ^ n3465;
  assign n3467 = ~n3392 ^ ~n3466;
  assign n3468 = ~n3290 & ~n3259;
  assign n3469 = ~n3468 & n3242;
  assign n3470 = n3290 & n3259;
  assign n3471 = ~n3469 & ~n3470;
  assign n3472 = n3311 & ~n3328;
  assign n3473 = ~n3294 & ~n3310;
  assign n3474 = ~n3472 & ~n3473;
  assign n3475 = n3254 & n3257;
  assign n3476 = n3251 & ~n3475;
  assign n3477 = ~n3254 & ~n3257;
  assign n3478 = ~n3476 & ~n3477;
  assign n3479 = ~n3266 & ~n3268;
  assign n3480 = n3265 & ~n3479;
  assign n3481 = n3308 & ~n1381;
  assign n3482 = ~n3306 & ~n3307;
  assign n3483 = ~n3481 & ~n3482;
  assign n3484 = ~n3480 ^ ~n3483;
  assign n3485 = n3302 & ~n3303;
  assign n3486 = ~n3300 & ~n3301;
  assign n3487 = ~n3485 & ~n3486;
  assign n3488 = ~n3484 ^ n3487;
  assign n3489 = pi12 & pi33;
  assign n3490 = pi11 & pi34;
  assign n3491 = ~n3489 ^ ~n3490;
  assign n3492 = pi06 & pi39;
  assign n3493 = ~n3491 ^ n3492;
  assign n3494 = pi16 & pi29;
  assign n3495 = pi17 & pi28;
  assign n3496 = ~n3494 ^ ~n3495;
  assign n3497 = pi15 & pi30;
  assign n3498 = ~n3496 ^ n3497;
  assign n3499 = ~n3493 ^ ~n3498;
  assign n3500 = pi21 & pi43;
  assign n3501 = n3500 & pi01;
  assign n3502 = ~n3501 & pi23;
  assign n3503 = pi03 & pi42;
  assign n3504 = pi01 & pi44;
  assign n3505 = ~n3503 ^ n3504;
  assign n3506 = ~n3502 ^ ~n3505;
  assign n3507 = ~n3499 ^ n3506;
  assign n3508 = ~n3488 ^ n3507;
  assign n3509 = ~n3478 ^ ~n3508;
  assign n3510 = ~n3474 ^ n3509;
  assign n3511 = ~n3471 ^ ~n3510;
  assign n3512 = ~n3467 ^ n3511;
  assign n3513 = ~n3388 ^ ~n3512;
  assign po046 = ~n3384 ^ n3513;
  assign n3515 = ~n3377 & n3513;
  assign n3516 = n3374 & ~n3515;
  assign n3517 = ~n3230 & ~n3516;
  assign n3518 = ~n3380 & n3513;
  assign n3519 = ~n3518 & ~n3382;
  assign n3520 = ~n3517 & n3519;
  assign n3521 = ~n3467 & n3511;
  assign n3522 = n3388 & ~n3521;
  assign n3523 = n3467 & ~n3511;
  assign n3524 = ~n3522 & ~n3523;
  assign n3525 = n3392 & n3466;
  assign n3526 = ~n3428 & n3465;
  assign n3527 = ~n3525 & ~n3526;
  assign n3528 = n3474 & ~n3509;
  assign n3529 = ~n3471 & ~n3528;
  assign n3530 = ~n3474 & n3509;
  assign n3531 = ~n3529 & ~n3530;
  assign n3532 = ~n3488 & n3507;
  assign n3533 = n3478 & ~n3532;
  assign n3534 = n3488 & ~n3507;
  assign n3535 = ~n3533 & ~n3534;
  assign n3536 = n3458 & ~n3463;
  assign n3537 = n3452 & ~n3457;
  assign n3538 = ~n3536 & ~n3537;
  assign n3539 = n3442 & n3447;
  assign n3540 = n3436 & n3441;
  assign n3541 = ~n3539 & ~n3540;
  assign n3542 = ~n3538 ^ n3541;
  assign n3543 = n3499 & ~n3506;
  assign n3544 = ~n3493 & ~n3498;
  assign n3545 = ~n3543 & ~n3544;
  assign n3546 = ~n3542 ^ n3545;
  assign n3547 = n3484 & ~n3487;
  assign n3548 = ~n3480 & ~n3483;
  assign n3549 = ~n3547 & ~n3548;
  assign n3550 = n3445 & ~n3446;
  assign n3551 = ~n3443 & ~n3444;
  assign n3552 = ~n3550 & ~n3551;
  assign n3553 = n3439 & ~n3440;
  assign n3554 = ~n3437 & ~n3438;
  assign n3555 = ~n3553 & ~n3554;
  assign n3556 = ~n3552 ^ ~n3555;
  assign n3557 = n3461 & ~n3462;
  assign n3558 = ~n3459 & ~n3460;
  assign n3559 = ~n3557 & ~n3558;
  assign n3560 = ~n3556 ^ n3559;
  assign n3561 = n3434 & ~n3435;
  assign n3562 = ~n3432 & ~n3433;
  assign n3563 = ~n3561 & ~n3562;
  assign n3564 = pi23 & pi44;
  assign n3565 = ~n3564 ^ ~pi45;
  assign n3566 = n3565 & pi01;
  assign n3567 = pi22 & pi24;
  assign n3568 = ~n3566 ^ n3567;
  assign n3569 = ~n3563 ^ ~n3568;
  assign n3570 = ~n3560 ^ ~n3569;
  assign n3571 = ~n3549 ^ n3570;
  assign n3572 = ~n3546 ^ n3571;
  assign n3573 = ~n3535 ^ n3572;
  assign n3574 = n3414 & ~n3425;
  assign n3575 = ~n3410 & ~n3413;
  assign n3576 = ~n3574 & ~n3575;
  assign n3577 = pi04 & pi42;
  assign n3578 = pi03 & pi43;
  assign n3579 = ~n3577 ^ ~n3578;
  assign n3580 = pi00 & pi46;
  assign n3581 = ~n3579 ^ n3580;
  assign n3582 = pi11 & pi35;
  assign n3583 = pi10 & pi36;
  assign n3584 = ~n3582 ^ ~n3583;
  assign n3585 = pi09 & pi37;
  assign n3586 = ~n3584 ^ n3585;
  assign n3587 = ~n3581 ^ ~n3586;
  assign n3588 = pi21 & pi25;
  assign n3589 = pi20 & pi26;
  assign n3590 = ~n3588 ^ ~n3589;
  assign n3591 = pi19 & pi27;
  assign n3592 = ~n3590 ^ n3591;
  assign n3593 = ~n3587 ^ ~n3592;
  assign n3594 = ~n3576 ^ ~n3593;
  assign n3595 = pi03 & pi44;
  assign n3596 = n3595 & pi42;
  assign n3597 = n3500 & pi23;
  assign n3598 = ~n3596 & ~n3597;
  assign n3599 = ~n3564 & pi01;
  assign n3600 = ~n3598 & n3599;
  assign n3601 = ~n3500 & n3504;
  assign n3602 = pi23 & pi42;
  assign n3603 = n3602 & pi03;
  assign n3604 = ~n3601 & n3603;
  assign n3605 = ~n3600 & ~n3604;
  assign n3606 = pi18 & pi28;
  assign n3607 = pi17 & pi29;
  assign n3608 = ~n3606 ^ ~n3607;
  assign n3609 = ~n3608 ^ n1814;
  assign n3610 = pi12 & pi34;
  assign n3611 = pi08 & pi38;
  assign n3612 = ~n3610 ^ ~n3611;
  assign n3613 = pi07 & pi39;
  assign n3614 = ~n3612 ^ n3613;
  assign n3615 = ~n3609 ^ ~n3614;
  assign n3616 = ~n3605 ^ n3615;
  assign n3617 = ~n3594 ^ ~n3616;
  assign n3618 = ~n3573 ^ n3617;
  assign n3619 = ~n3531 ^ n3618;
  assign n3620 = ~n3407 & ~n3426;
  assign n3621 = n3396 & ~n3620;
  assign n3622 = n3407 & n3426;
  assign n3623 = ~n3621 & ~n3622;
  assign n3624 = n3449 & ~n3464;
  assign n3625 = n3431 & n3448;
  assign n3626 = ~n3624 & ~n3625;
  assign n3627 = n3403 & ~n3406;
  assign n3628 = ~n3399 & ~n3402;
  assign n3629 = ~n3627 & ~n3628;
  assign n3630 = n3421 & ~n3424;
  assign n3631 = ~n3417 & ~n3420;
  assign n3632 = ~n3630 & ~n3631;
  assign n3633 = pi14 & pi32;
  assign n3634 = pi13 & pi33;
  assign n3635 = ~n3633 ^ ~n3634;
  assign n3636 = pi06 & pi40;
  assign n3637 = ~n3635 ^ n3636;
  assign n3638 = pi05 & pi41;
  assign n3639 = ~n1978 ^ ~n3638;
  assign n3640 = pi02 & pi44;
  assign n3641 = ~n3639 ^ n3640;
  assign n3642 = ~n3637 ^ ~n3641;
  assign n3643 = ~n3632 ^ n3642;
  assign n3644 = n3491 & ~n3492;
  assign n3645 = ~n3489 & ~n3490;
  assign n3646 = ~n3644 & ~n3645;
  assign n3647 = n3496 & ~n3497;
  assign n3648 = ~n3494 & ~n3495;
  assign n3649 = ~n3647 & ~n3648;
  assign n3650 = ~n3646 ^ ~n3649;
  assign n3651 = n3455 & ~n3456;
  assign n3652 = ~n3453 & ~n3454;
  assign n3653 = ~n3651 & ~n3652;
  assign n3654 = ~n3650 ^ ~n3653;
  assign n3655 = ~n3643 ^ n3654;
  assign n3656 = ~n3629 ^ n3655;
  assign n3657 = ~n3626 ^ ~n3656;
  assign n3658 = ~n3623 ^ n3657;
  assign n3659 = ~n3619 ^ ~n3658;
  assign n3660 = ~n3527 ^ n3659;
  assign n3661 = ~n3524 ^ ~n3660;
  assign po047 = ~n3520 ^ ~n3661;
  assign n3663 = n3619 & ~n3658;
  assign n3664 = n3527 & ~n3663;
  assign n3665 = ~n3619 & n3658;
  assign n3666 = ~n3664 & ~n3665;
  assign n3667 = n3524 & ~n3666;
  assign n3668 = n3527 & n3665;
  assign n3669 = ~n3667 & ~n3668;
  assign n3670 = n3520 & ~n3669;
  assign n3671 = n3524 & n3668;
  assign n3672 = ~n3670 & ~n3671;
  assign n3673 = ~n3527 & n3663;
  assign n3674 = n3524 & ~n3673;
  assign n3675 = ~n3674 & n3666;
  assign n3676 = ~n3520 & n3675;
  assign n3677 = ~n3524 & n3673;
  assign n3678 = ~n3676 & ~n3677;
  assign n3679 = n3672 & n3678;
  assign n3680 = ~n3626 & ~n3656;
  assign n3681 = ~n3623 & ~n3680;
  assign n3682 = n3626 & n3656;
  assign n3683 = ~n3681 & ~n3682;
  assign n3684 = n3546 & ~n3571;
  assign n3685 = ~n3535 & ~n3684;
  assign n3686 = ~n3546 & n3571;
  assign n3687 = ~n3685 & ~n3686;
  assign n3688 = n3643 & ~n3654;
  assign n3689 = ~n3629 & ~n3688;
  assign n3690 = ~n3643 & n3654;
  assign n3691 = ~n3689 & ~n3690;
  assign n3692 = n3594 & n3616;
  assign n3693 = ~n3576 & ~n3593;
  assign n3694 = ~n3692 & ~n3693;
  assign n3695 = ~n3632 & n3642;
  assign n3696 = n3637 & n3641;
  assign n3697 = ~n3695 & ~n3696;
  assign n3698 = n3590 & ~n3591;
  assign n3699 = ~n3588 & ~n3589;
  assign n3700 = ~n3698 & ~n3699;
  assign n3701 = n3579 & ~n3580;
  assign n3702 = ~n3577 & ~n3578;
  assign n3703 = ~n3701 & ~n3702;
  assign n3704 = ~n3700 ^ ~n3703;
  assign n3705 = n3639 & ~n3640;
  assign n3706 = ~n1978 & ~n3638;
  assign n3707 = ~n3705 & ~n3706;
  assign n3708 = ~n3704 ^ ~n3707;
  assign n3709 = ~n3697 ^ ~n3708;
  assign n3710 = n3587 & n3592;
  assign n3711 = n3581 & n3586;
  assign n3712 = ~n3710 & ~n3711;
  assign n3713 = ~n3709 ^ n3712;
  assign n3714 = ~n3694 ^ ~n3713;
  assign n3715 = ~n3691 ^ n3714;
  assign n3716 = ~n3687 ^ ~n3715;
  assign n3717 = ~n3683 ^ ~n3716;
  assign n3718 = n3542 & ~n3545;
  assign n3719 = ~n3538 & n3541;
  assign n3720 = ~n3718 & ~n3719;
  assign n3721 = ~n3549 & n3570;
  assign n3722 = n3560 & n3569;
  assign n3723 = ~n3721 & ~n3722;
  assign n3724 = ~n3567 ^ pi45;
  assign n3725 = ~n3724 & n3564;
  assign n3726 = ~n3563 & ~n3725;
  assign n3727 = n3724 & ~n3564;
  assign n3728 = ~n3727 & pi01;
  assign n3729 = ~n3726 & n3728;
  assign n3730 = n3567 & ~pi01;
  assign n3731 = n3563 & n3730;
  assign n3732 = ~n3729 & ~n3731;
  assign n3733 = pi13 & pi34;
  assign n3734 = pi12 & pi35;
  assign n3735 = ~n3733 ^ ~n3734;
  assign n3736 = pi07 & pi40;
  assign n3737 = ~n3735 ^ n3736;
  assign n3738 = ~n3732 ^ ~n3737;
  assign n3739 = n3650 & n3653;
  assign n3740 = n3646 & n3649;
  assign n3741 = ~n3739 & ~n3740;
  assign n3742 = ~n3738 ^ ~n3741;
  assign n3743 = ~n3723 ^ n3742;
  assign n3744 = ~n3720 ^ ~n3743;
  assign n3745 = ~n3605 & n3615;
  assign n3746 = ~n3609 & ~n3614;
  assign n3747 = ~n3745 & ~n3746;
  assign n3748 = n3612 & ~n3613;
  assign n3749 = ~n3610 & ~n3611;
  assign n3750 = ~n3748 & ~n3749;
  assign n3751 = n3584 & ~n3585;
  assign n3752 = ~n3582 & ~n3583;
  assign n3753 = ~n3751 & ~n3752;
  assign n3754 = ~n3750 ^ ~n3753;
  assign n3755 = pi01 & pi46;
  assign n3756 = ~n3755 ^ ~pi24;
  assign n3757 = ~n3754 ^ ~n3756;
  assign n3758 = ~n3747 ^ n3757;
  assign n3759 = n3556 & ~n3559;
  assign n3760 = ~n3552 & ~n3555;
  assign n3761 = ~n3759 & ~n3760;
  assign n3762 = ~n3758 ^ ~n3761;
  assign n3763 = n3608 & ~n1814;
  assign n3764 = ~n3606 & ~n3607;
  assign n3765 = ~n3763 & ~n3764;
  assign n3766 = n3635 & ~n3636;
  assign n3767 = ~n3633 & ~n3634;
  assign n3768 = ~n3766 & ~n3767;
  assign n3769 = ~n3765 ^ ~n3768;
  assign n3770 = pi15 & pi32;
  assign n3771 = pi04 & pi43;
  assign n3772 = ~n3770 ^ ~n3771;
  assign n3773 = ~n3772 ^ n3595;
  assign n3774 = ~n3769 ^ n3773;
  assign n3775 = n1057 & pi24;
  assign n3776 = ~n3775 ^ ~pi02;
  assign n3777 = n3776 & pi45;
  assign n3778 = pi00 & pi47;
  assign n3779 = ~n3777 ^ ~n3778;
  assign n3780 = pi21 & pi26;
  assign n3781 = pi20 & pi27;
  assign n3782 = ~n3780 ^ ~n3781;
  assign n3783 = pi19 & pi28;
  assign n3784 = ~n3782 ^ n3783;
  assign n3785 = pi18 & pi29;
  assign n3786 = pi17 & pi30;
  assign n3787 = ~n3785 ^ ~n3786;
  assign n3788 = pi16 & pi31;
  assign n3789 = ~n3787 ^ n3788;
  assign n3790 = ~n3784 ^ ~n3789;
  assign n3791 = ~n3779 ^ ~n3790;
  assign n3792 = ~n3774 ^ ~n3791;
  assign n3793 = pi14 & pi33;
  assign n3794 = pi06 & pi41;
  assign n3795 = ~n3793 ^ ~n3794;
  assign n3796 = pi05 & pi42;
  assign n3797 = ~n3795 ^ n3796;
  assign n3798 = pi11 & pi36;
  assign n3799 = pi09 & pi38;
  assign n3800 = ~n3798 ^ ~n3799;
  assign n3801 = pi08 & pi39;
  assign n3802 = ~n3800 ^ n3801;
  assign n3803 = ~n3797 ^ ~n3802;
  assign n3804 = pi23 & pi24;
  assign n3805 = pi22 & pi25;
  assign n3806 = ~n3804 ^ ~n3805;
  assign n3807 = pi10 & pi37;
  assign n3808 = ~n3806 ^ n3807;
  assign n3809 = ~n3803 ^ n3808;
  assign n3810 = ~n3792 ^ ~n3809;
  assign n3811 = ~n3762 ^ ~n3810;
  assign n3812 = ~n3744 ^ ~n3811;
  assign n3813 = ~n3717 ^ ~n3812;
  assign n3814 = ~n3573 & n3617;
  assign n3815 = ~n3531 & ~n3814;
  assign n3816 = n3573 & ~n3617;
  assign n3817 = ~n3815 & ~n3816;
  assign n3818 = ~n3813 ^ n3817;
  assign po048 = ~n3679 ^ n3818;
  assign n3820 = ~n3671 & n3818;
  assign n3821 = ~n3675 & ~n3820;
  assign n3822 = ~n3520 & ~n3821;
  assign n3823 = ~n3677 & ~n3818;
  assign n3824 = n3669 & ~n3823;
  assign n3825 = ~n3822 & ~n3824;
  assign n3826 = ~n3717 & ~n3812;
  assign n3827 = ~n3826 & ~n3817;
  assign n3828 = n3717 & n3812;
  assign n3829 = ~n3827 & ~n3828;
  assign n3830 = n3687 & n3715;
  assign n3831 = n3683 & ~n3830;
  assign n3832 = ~n3687 & ~n3715;
  assign n3833 = ~n3831 & ~n3832;
  assign n3834 = ~n3694 & ~n3713;
  assign n3835 = n3691 & ~n3834;
  assign n3836 = n3694 & n3713;
  assign n3837 = ~n3835 & ~n3836;
  assign n3838 = n3738 & n3741;
  assign n3839 = n3732 & n3737;
  assign n3840 = ~n3838 & ~n3839;
  assign n3841 = pi14 & pi34;
  assign n3842 = pi13 & pi35;
  assign n3843 = ~n3841 ^ ~n3842;
  assign n3844 = pi06 & pi42;
  assign n3845 = ~n3843 ^ n3844;
  assign n3846 = pi12 & pi36;
  assign n3847 = pi08 & pi40;
  assign n3848 = ~n3846 ^ ~n3847;
  assign n3849 = pi07 & pi41;
  assign n3850 = ~n3848 ^ n3849;
  assign n3851 = ~n3845 ^ ~n3850;
  assign n3852 = pi11 & pi37;
  assign n3853 = pi10 & pi38;
  assign n3854 = ~n3852 ^ ~n3853;
  assign n3855 = pi09 & pi39;
  assign n3856 = ~n3854 ^ n3855;
  assign n3857 = ~n3851 ^ n3856;
  assign n3858 = ~n3840 ^ ~n3857;
  assign n3859 = pi19 & pi29;
  assign n3860 = pi18 & pi30;
  assign n3861 = ~n3859 ^ ~n3860;
  assign n3862 = ~n3861 ^ n2010;
  assign n3863 = pi15 & pi33;
  assign n3864 = pi05 & pi43;
  assign n3865 = ~n3863 ^ ~n3864;
  assign n3866 = pi04 & pi44;
  assign n3867 = ~n3865 ^ n3866;
  assign n3868 = ~n3862 ^ ~n3867;
  assign n3869 = pi22 & pi26;
  assign n3870 = pi21 & pi27;
  assign n3871 = ~n3869 ^ ~n3870;
  assign n3872 = pi20 & pi28;
  assign n3873 = ~n3871 ^ n3872;
  assign n3874 = ~n3868 ^ n3873;
  assign n3875 = ~n3858 ^ n3874;
  assign n3876 = n3723 & ~n3742;
  assign n3877 = n3720 & ~n3876;
  assign n3878 = ~n3723 & n3742;
  assign n3879 = ~n3877 & ~n3878;
  assign n3880 = ~n3875 ^ n3879;
  assign n3881 = ~n3837 ^ ~n3880;
  assign n3882 = n3744 & n3811;
  assign n3883 = ~n3762 & ~n3810;
  assign n3884 = ~n3882 & ~n3883;
  assign n3885 = n3754 & n3756;
  assign n3886 = n3750 & n3753;
  assign n3887 = ~n3885 & ~n3886;
  assign n3888 = ~n3778 & ~pi02;
  assign n3889 = n3775 & ~n3888;
  assign n3890 = n3778 & pi02;
  assign n3891 = ~n3889 & ~n3890;
  assign n3892 = ~n3891 & pi45;
  assign n3893 = n3787 & ~n3788;
  assign n3894 = ~n3785 & ~n3786;
  assign n3895 = ~n3893 & ~n3894;
  assign n3896 = n3772 & ~n3595;
  assign n3897 = ~n3770 & ~n3771;
  assign n3898 = ~n3896 & ~n3897;
  assign n3899 = ~n3895 ^ ~n3898;
  assign n3900 = ~n3892 ^ ~n3899;
  assign n3901 = ~n3887 ^ n3900;
  assign n3902 = n3779 & n3790;
  assign n3903 = ~n3784 & ~n3789;
  assign n3904 = ~n3902 & ~n3903;
  assign n3905 = ~n3901 ^ n3904;
  assign n3906 = n3803 & ~n3808;
  assign n3907 = ~n3797 & ~n3802;
  assign n3908 = ~n3906 & ~n3907;
  assign n3909 = n3735 & ~n3736;
  assign n3910 = ~n3733 & ~n3734;
  assign n3911 = ~n3909 & ~n3910;
  assign n3912 = pi16 & pi32;
  assign n3913 = pi03 & pi45;
  assign n3914 = ~n3912 ^ ~n3913;
  assign n3915 = pi02 & pi46;
  assign n3916 = ~n3914 ^ n3915;
  assign n3917 = ~n3911 ^ n3916;
  assign n3918 = n3806 & ~n3807;
  assign n3919 = ~n3804 & ~n3805;
  assign n3920 = ~n3918 & ~n3919;
  assign n3921 = ~n3917 ^ n3920;
  assign n3922 = ~n3908 ^ ~n3921;
  assign n3923 = n3795 & ~n3796;
  assign n3924 = ~n3793 & ~n3794;
  assign n3925 = ~n3923 & ~n3924;
  assign n3926 = n3782 & ~n3783;
  assign n3927 = ~n3780 & ~n3781;
  assign n3928 = ~n3926 & ~n3927;
  assign n3929 = ~n3925 ^ ~n3928;
  assign n3930 = n3800 & ~n3801;
  assign n3931 = ~n3798 & ~n3799;
  assign n3932 = ~n3930 & ~n3931;
  assign n3933 = ~n3929 ^ n3932;
  assign n3934 = ~n3922 ^ n3933;
  assign n3935 = ~n3905 ^ ~n3934;
  assign n3936 = ~n3810 & n3791;
  assign n3937 = n3774 & n3809;
  assign n3938 = ~n3936 & ~n3937;
  assign n3939 = ~n3935 ^ ~n3938;
  assign n3940 = ~n3884 ^ n3939;
  assign n3941 = n3709 & ~n3712;
  assign n3942 = ~n3697 & ~n3708;
  assign n3943 = ~n3941 & ~n3942;
  assign n3944 = n3758 & n3761;
  assign n3945 = ~n3747 & n3757;
  assign n3946 = ~n3944 & ~n3945;
  assign n3947 = n3704 & n3707;
  assign n3948 = n3700 & n3703;
  assign n3949 = ~n3947 & ~n3948;
  assign n3950 = n1185 & pi46;
  assign n3951 = pi01 & pi47;
  assign n3952 = pi23 & pi25;
  assign n3953 = ~n3951 ^ ~n3952;
  assign n3954 = ~n3950 ^ ~n3953;
  assign n3955 = pi00 & pi48;
  assign n3956 = ~n3954 ^ n3955;
  assign n3957 = ~n3949 ^ ~n3956;
  assign n3958 = n3769 & ~n3773;
  assign n3959 = n3765 & n3768;
  assign n3960 = ~n3958 & ~n3959;
  assign n3961 = ~n3957 ^ ~n3960;
  assign n3962 = ~n3946 ^ ~n3961;
  assign n3963 = ~n3943 ^ ~n3962;
  assign n3964 = ~n3940 ^ n3963;
  assign n3965 = ~n3881 ^ n3964;
  assign n3966 = ~n3833 ^ n3965;
  assign n3967 = ~n3829 ^ n3966;
  assign po049 = n3825 ^ n3967;
  assign n3969 = n3829 & ~n3966;
  assign n3970 = ~n3825 & ~n3969;
  assign n3971 = ~n3829 & n3966;
  assign n3972 = ~n3970 & ~n3971;
  assign n3973 = n3881 & ~n3964;
  assign n3974 = ~n3833 & ~n3973;
  assign n3975 = ~n3881 & n3964;
  assign n3976 = ~n3974 & ~n3975;
  assign n3977 = n3875 & ~n3879;
  assign n3978 = n3837 & ~n3977;
  assign n3979 = ~n3875 & n3879;
  assign n3980 = ~n3978 & ~n3979;
  assign n3981 = n3858 & ~n3874;
  assign n3982 = ~n3840 & ~n3857;
  assign n3983 = ~n3981 & ~n3982;
  assign n3984 = n3957 & n3960;
  assign n3985 = n3949 & n3956;
  assign n3986 = ~n3984 & ~n3985;
  assign n3987 = n3868 & ~n3873;
  assign n3988 = ~n3862 & ~n3867;
  assign n3989 = ~n3987 & ~n3988;
  assign n3990 = ~n3986 ^ n3989;
  assign n3991 = n3861 & ~n2010;
  assign n3992 = ~n3859 & ~n3860;
  assign n3993 = ~n3991 & ~n3992;
  assign n3994 = n3848 & ~n3849;
  assign n3995 = ~n3846 & ~n3847;
  assign n3996 = ~n3994 & ~n3995;
  assign n3997 = ~n3993 ^ ~n3996;
  assign n3998 = n3843 & ~n3844;
  assign n3999 = ~n3841 & ~n3842;
  assign n4000 = ~n3998 & ~n3999;
  assign n4001 = ~n3997 ^ n4000;
  assign n4002 = ~n3990 ^ n4001;
  assign n4003 = n3851 & ~n3856;
  assign n4004 = ~n3845 & ~n3850;
  assign n4005 = ~n4003 & ~n4004;
  assign n4006 = n3854 & ~n3855;
  assign n4007 = ~n3852 & ~n3853;
  assign n4008 = ~n4006 & ~n4007;
  assign n4009 = pi23 & pi47;
  assign n4010 = n4009 & pi01;
  assign n4011 = ~n4010 & pi25;
  assign n4012 = pi01 & pi48;
  assign n4013 = ~n4011 ^ n4012;
  assign n4014 = ~n4008 ^ n4013;
  assign n4015 = ~n4005 ^ n4014;
  assign n4016 = n3865 & ~n3866;
  assign n4017 = ~n3863 & ~n3864;
  assign n4018 = ~n4016 & ~n4017;
  assign n4019 = n3914 & ~n3915;
  assign n4020 = ~n3912 & ~n3913;
  assign n4021 = ~n4019 & ~n4020;
  assign n4022 = ~n4018 ^ ~n4021;
  assign n4023 = n3871 & ~n3872;
  assign n4024 = ~n3869 & ~n3870;
  assign n4025 = ~n4023 & ~n4024;
  assign n4026 = ~n4022 ^ ~n4025;
  assign n4027 = ~n4015 ^ ~n4026;
  assign n4028 = ~n4002 ^ ~n4027;
  assign n4029 = ~n3983 ^ ~n4028;
  assign n4030 = n3901 & ~n3904;
  assign n4031 = ~n3887 & n3900;
  assign n4032 = ~n4030 & ~n4031;
  assign n4033 = n3922 & ~n3933;
  assign n4034 = ~n3908 & ~n3921;
  assign n4035 = ~n4033 & ~n4034;
  assign n4036 = n3929 & ~n3932;
  assign n4037 = ~n3925 & ~n3928;
  assign n4038 = ~n4036 & ~n4037;
  assign n4039 = n3917 & ~n3920;
  assign n4040 = ~n3911 & n3916;
  assign n4041 = ~n4039 & ~n4040;
  assign n4042 = ~n4038 ^ ~n4041;
  assign n4043 = n3892 & n3899;
  assign n4044 = n3895 & n3898;
  assign n4045 = ~n4043 & ~n4044;
  assign n4046 = ~n4042 ^ ~n4045;
  assign n4047 = ~n4035 ^ ~n4046;
  assign n4048 = ~n4032 ^ n4047;
  assign n4049 = ~n4029 ^ ~n4048;
  assign n4050 = ~n3980 ^ n4049;
  assign n4051 = ~n3884 & n3939;
  assign n4052 = ~n4051 & n3963;
  assign n4053 = n3884 & ~n3939;
  assign n4054 = ~n4052 & ~n4053;
  assign n4055 = ~n3946 & ~n3961;
  assign n4056 = ~n3943 & ~n4055;
  assign n4057 = n3946 & n3961;
  assign n4058 = ~n4056 & ~n4057;
  assign n4059 = ~n3905 & ~n3934;
  assign n4060 = ~n4059 & ~n3938;
  assign n4061 = n3905 & n3934;
  assign n4062 = ~n4060 & ~n4061;
  assign n4063 = n3956 & n3953;
  assign n4064 = n3950 & n3955;
  assign n4065 = ~n4063 & ~n4064;
  assign n4066 = pi18 & pi31;
  assign n4067 = ~n2013 ^ ~n4066;
  assign n4068 = pi16 & pi33;
  assign n4069 = ~n4067 ^ n4068;
  assign n4070 = pi05 & pi44;
  assign n4071 = pi04 & pi45;
  assign n4072 = ~n4070 ^ ~n4071;
  assign n4073 = pi00 & pi49;
  assign n4074 = ~n4072 ^ n4073;
  assign n4075 = ~n4069 ^ ~n4074;
  assign n4076 = ~n4065 ^ n4075;
  assign n4077 = pi24 & pi25;
  assign n4078 = pi23 & pi26;
  assign n4079 = ~n4077 ^ ~n4078;
  assign n4080 = pi11 & pi38;
  assign n4081 = ~n4079 ^ n4080;
  assign n4082 = pi15 & pi34;
  assign n4083 = pi14 & pi35;
  assign n4084 = ~n4082 ^ ~n4083;
  assign n4085 = pi06 & pi43;
  assign n4086 = ~n4084 ^ n4085;
  assign n4087 = ~n4081 ^ ~n4086;
  assign n4088 = pi13 & pi36;
  assign n4089 = pi08 & pi41;
  assign n4090 = ~n4088 ^ ~n4089;
  assign n4091 = pi07 & pi42;
  assign n4092 = ~n4090 ^ n4091;
  assign n4093 = ~n4087 ^ n4092;
  assign n4094 = ~n4076 ^ ~n4093;
  assign n4095 = pi21 & pi28;
  assign n4096 = pi20 & pi29;
  assign n4097 = ~n4095 ^ ~n4096;
  assign n4098 = pi19 & pi30;
  assign n4099 = ~n4097 ^ n4098;
  assign n4100 = pi22 & pi27;
  assign n4101 = pi03 & pi46;
  assign n4102 = ~n4100 ^ ~n4101;
  assign n4103 = pi02 & pi47;
  assign n4104 = ~n4102 ^ n4103;
  assign n4105 = ~n4099 ^ ~n4104;
  assign n4106 = pi12 & pi37;
  assign n4107 = pi10 & pi39;
  assign n4108 = ~n4106 ^ ~n4107;
  assign n4109 = pi09 & pi40;
  assign n4110 = ~n4108 ^ n4109;
  assign n4111 = ~n4105 ^ n4110;
  assign n4112 = ~n4094 ^ ~n4111;
  assign n4113 = ~n4062 ^ n4112;
  assign n4114 = ~n4058 ^ ~n4113;
  assign n4115 = ~n4054 ^ ~n4114;
  assign n4116 = ~n4050 ^ ~n4115;
  assign n4117 = ~n3976 ^ n4116;
  assign po050 = n3972 ^ n4117;
  assign n4119 = n4054 & ~n4114;
  assign n4120 = ~n4050 & n4119;
  assign n4121 = n3976 & ~n4120;
  assign n4122 = n4050 & ~n4119;
  assign n4123 = ~n4054 & n4114;
  assign n4124 = ~n4122 & ~n4123;
  assign n4125 = ~n4121 & n4124;
  assign n4126 = ~n3972 & n4125;
  assign n4127 = ~n3976 & n4120;
  assign n4128 = ~n4126 & ~n4127;
  assign n4129 = ~n4124 & n3976;
  assign n4130 = n4050 & n4123;
  assign n4131 = ~n4129 & ~n4130;
  assign n4132 = n3972 & ~n4131;
  assign n4133 = n3976 & n4130;
  assign n4134 = ~n4132 & ~n4133;
  assign n4135 = n4128 & n4134;
  assign n4136 = n4029 & n4048;
  assign n4137 = n3980 & ~n4136;
  assign n4138 = ~n4029 & ~n4048;
  assign n4139 = ~n4137 & ~n4138;
  assign n4140 = ~n4062 & n4112;
  assign n4141 = ~n4058 & ~n4140;
  assign n4142 = n4062 & ~n4112;
  assign n4143 = ~n4141 & ~n4142;
  assign n4144 = n3990 & ~n4001;
  assign n4145 = n3986 & ~n3989;
  assign n4146 = ~n4144 & ~n4145;
  assign n4147 = n4015 & n4026;
  assign n4148 = ~n4005 & n4014;
  assign n4149 = ~n4147 & ~n4148;
  assign n4150 = n3997 & ~n4000;
  assign n4151 = ~n3993 & ~n3996;
  assign n4152 = ~n4150 & ~n4151;
  assign n4153 = n4022 & n4025;
  assign n4154 = n4018 & n4021;
  assign n4155 = ~n4153 & ~n4154;
  assign n4156 = ~n4152 ^ n4155;
  assign n4157 = n4084 & ~n4085;
  assign n4158 = ~n4082 & ~n4083;
  assign n4159 = ~n4157 & ~n4158;
  assign n4160 = n4102 & ~n4103;
  assign n4161 = ~n4100 & ~n4101;
  assign n4162 = ~n4160 & ~n4161;
  assign n4163 = ~n4159 ^ ~n4162;
  assign n4164 = n4072 & ~n4073;
  assign n4165 = ~n4070 & ~n4071;
  assign n4166 = ~n4164 & ~n4165;
  assign n4167 = ~n4163 ^ ~n4166;
  assign n4168 = ~n4156 ^ ~n4167;
  assign n4169 = ~n4149 ^ n4168;
  assign n4170 = ~n4146 ^ ~n4169;
  assign n4171 = n4094 & n4111;
  assign n4172 = n4076 & n4093;
  assign n4173 = ~n4171 & ~n4172;
  assign n4174 = ~n4065 & n4075;
  assign n4175 = ~n4069 & ~n4074;
  assign n4176 = ~n4174 & ~n4175;
  assign n4177 = n4105 & ~n4110;
  assign n4178 = ~n4099 & ~n4104;
  assign n4179 = ~n4177 & ~n4178;
  assign n4180 = n4108 & ~n4109;
  assign n4181 = ~n4106 & ~n4107;
  assign n4182 = ~n4180 & ~n4181;
  assign n4183 = n4079 & ~n4080;
  assign n4184 = ~n4077 & ~n4078;
  assign n4185 = ~n4183 & ~n4184;
  assign n4186 = ~n4182 ^ ~n4185;
  assign n4187 = pi01 & pi49;
  assign n4188 = pi24 & pi26;
  assign n4189 = ~n4187 ^ ~n4188;
  assign n4190 = ~n4186 ^ ~n4189;
  assign n4191 = ~n4179 ^ n4190;
  assign n4192 = ~n4176 ^ n4191;
  assign n4193 = ~n4173 ^ n4192;
  assign n4194 = n4038 & n4041;
  assign n4195 = ~n4194 & n4045;
  assign n4196 = ~n4038 & ~n4041;
  assign n4197 = ~n4195 & ~n4196;
  assign n4198 = n4087 & ~n4092;
  assign n4199 = ~n4081 & ~n4086;
  assign n4200 = ~n4198 & ~n4199;
  assign n4201 = n4097 & ~n4098;
  assign n4202 = ~n4095 & ~n4096;
  assign n4203 = ~n4201 & ~n4202;
  assign n4204 = n4090 & ~n4091;
  assign n4205 = ~n4088 & ~n4089;
  assign n4206 = ~n4204 & ~n4205;
  assign n4207 = ~n4203 ^ ~n4206;
  assign n4208 = n4067 & ~n4068;
  assign n4209 = ~n2013 & ~n4066;
  assign n4210 = ~n4208 & ~n4209;
  assign n4211 = ~n4207 ^ ~n4210;
  assign n4212 = ~n4200 ^ n4211;
  assign n4213 = ~n4197 ^ ~n4212;
  assign n4214 = ~n4193 ^ ~n4213;
  assign n4215 = ~n4170 ^ n4214;
  assign n4216 = ~n4143 ^ ~n4215;
  assign n4217 = ~n4002 & ~n4027;
  assign n4218 = n3983 & ~n4217;
  assign n4219 = n4002 & n4027;
  assign n4220 = ~n4218 & ~n4219;
  assign n4221 = n4035 & n4046;
  assign n4222 = ~n4032 & ~n4221;
  assign n4223 = ~n4035 & ~n4046;
  assign n4224 = ~n4222 & ~n4223;
  assign n4225 = n4008 & pi48;
  assign n4226 = pi25 & pi47;
  assign n4227 = n4226 & pi23;
  assign n4228 = ~n4225 & ~n4227;
  assign n4229 = pi25 & pi48;
  assign n4230 = ~n4229 & pi01;
  assign n4231 = ~n4228 & n4230;
  assign n4232 = ~n4009 & n4012;
  assign n4233 = ~n4232 & pi25;
  assign n4234 = n4008 & n4233;
  assign n4235 = ~n4231 & ~n4234;
  assign n4236 = pi23 & pi27;
  assign n4237 = pi22 & pi28;
  assign n4238 = ~n4236 ^ ~n4237;
  assign n4239 = pi18 & pi32;
  assign n4240 = ~n4238 ^ n4239;
  assign n4241 = pi16 & pi34;
  assign n4242 = pi15 & pi35;
  assign n4243 = ~n4241 ^ ~n4242;
  assign n4244 = pi05 & pi45;
  assign n4245 = ~n4243 ^ n4244;
  assign n4246 = ~n4240 ^ ~n4245;
  assign n4247 = ~n4235 ^ ~n4246;
  assign n4248 = ~n1306 & ~pi02;
  assign n4249 = ~n4248 & pi48;
  assign n4250 = n1306 & pi02;
  assign n4251 = n4249 & ~n4250;
  assign n4252 = pi00 & pi50;
  assign n4253 = ~n4251 ^ ~n4252;
  assign n4254 = pi17 & pi33;
  assign n4255 = pi04 & pi46;
  assign n4256 = ~n4254 ^ ~n4255;
  assign n4257 = pi03 & pi47;
  assign n4258 = ~n4256 ^ n4257;
  assign n4259 = pi21 & pi29;
  assign n4260 = pi20 & pi30;
  assign n4261 = ~n4259 ^ ~n4260;
  assign n4262 = pi19 & pi31;
  assign n4263 = ~n4261 ^ n4262;
  assign n4264 = ~n4258 ^ ~n4263;
  assign n4265 = ~n4253 ^ n4264;
  assign n4266 = pi14 & pi36;
  assign n4267 = pi07 & pi43;
  assign n4268 = ~n4266 ^ ~n4267;
  assign n4269 = pi06 & pi44;
  assign n4270 = ~n4268 ^ n4269;
  assign n4271 = pi12 & pi38;
  assign n4272 = pi11 & pi39;
  assign n4273 = ~n4271 ^ ~n4272;
  assign n4274 = pi10 & pi40;
  assign n4275 = ~n4273 ^ n4274;
  assign n4276 = ~n4270 ^ ~n4275;
  assign n4277 = pi13 & pi37;
  assign n4278 = pi09 & pi41;
  assign n4279 = ~n4277 ^ ~n4278;
  assign n4280 = pi08 & pi42;
  assign n4281 = ~n4279 ^ n4280;
  assign n4282 = ~n4276 ^ ~n4281;
  assign n4283 = ~n4265 ^ ~n4282;
  assign n4284 = ~n4247 ^ n4283;
  assign n4285 = ~n4224 ^ n4284;
  assign n4286 = ~n4220 ^ ~n4285;
  assign n4287 = ~n4216 ^ n4286;
  assign n4288 = ~n4139 ^ n4287;
  assign po051 = ~n4135 ^ n4288;
  assign n4290 = ~n4125 & ~n4288;
  assign n4291 = ~n4290 & ~n4133;
  assign n4292 = ~n3972 & n4291;
  assign n4293 = ~n4127 & ~n4288;
  assign n4294 = n4131 & ~n4293;
  assign n4295 = ~n4292 & ~n4294;
  assign n4296 = ~n4216 & n4286;
  assign n4297 = n4139 & ~n4296;
  assign n4298 = n4216 & ~n4286;
  assign n4299 = ~n4297 & ~n4298;
  assign n4300 = n4170 & ~n4214;
  assign n4301 = n4143 & ~n4300;
  assign n4302 = ~n4170 & n4214;
  assign n4303 = ~n4301 & ~n4302;
  assign n4304 = ~n4149 & n4168;
  assign n4305 = n4146 & ~n4304;
  assign n4306 = n4149 & ~n4168;
  assign n4307 = ~n4305 & ~n4306;
  assign n4308 = n4173 & ~n4192;
  assign n4309 = ~n4308 & n4213;
  assign n4310 = ~n4173 & n4192;
  assign n4311 = ~n4309 & ~n4310;
  assign n4312 = n4207 & n4210;
  assign n4313 = n4203 & n4206;
  assign n4314 = ~n4312 & ~n4313;
  assign n4315 = pi24 & pi49;
  assign n4316 = n4315 & pi01;
  assign n4317 = ~n4316 & pi26;
  assign n4318 = pi00 & pi51;
  assign n4319 = pi01 & pi50;
  assign n4320 = ~n4318 ^ n4319;
  assign n4321 = ~n4317 ^ ~n4320;
  assign n4322 = ~n4314 ^ ~n4321;
  assign n4323 = pi20 & pi31;
  assign n4324 = pi19 & pi32;
  assign n4325 = ~n4323 ^ ~n4324;
  assign n4326 = pi17 & pi34;
  assign n4327 = ~n4325 ^ n4326;
  assign n4328 = ~n4322 ^ ~n4327;
  assign n4329 = pi25 & pi26;
  assign n4330 = pi24 & pi27;
  assign n4331 = ~n4329 ^ ~n4330;
  assign n4332 = pi11 & pi40;
  assign n4333 = ~n4331 ^ n4332;
  assign n4334 = pi13 & pi38;
  assign n4335 = pi08 & pi43;
  assign n4336 = ~n4334 ^ ~n4335;
  assign n4337 = pi07 & pi44;
  assign n4338 = ~n4336 ^ n4337;
  assign n4339 = ~n4333 ^ ~n4338;
  assign n4340 = pi12 & pi39;
  assign n4341 = pi10 & pi41;
  assign n4342 = ~n4340 ^ ~n4341;
  assign n4343 = pi09 & pi42;
  assign n4344 = ~n4342 ^ n4343;
  assign n4345 = ~n4339 ^ n4344;
  assign n4346 = pi15 & pi36;
  assign n4347 = pi14 & pi37;
  assign n4348 = ~n4346 ^ ~n4347;
  assign n4349 = pi06 & pi45;
  assign n4350 = ~n4348 ^ n4349;
  assign n4351 = pi23 & pi28;
  assign n4352 = pi22 & pi29;
  assign n4353 = ~n4351 ^ ~n4352;
  assign n4354 = pi21 & pi30;
  assign n4355 = ~n4353 ^ n4354;
  assign n4356 = ~n4350 ^ ~n4355;
  assign n4357 = pi18 & pi33;
  assign n4358 = pi16 & pi35;
  assign n4359 = ~n4357 ^ ~n4358;
  assign n4360 = pi05 & pi46;
  assign n4361 = ~n4359 ^ n4360;
  assign n4362 = ~n4356 ^ ~n4361;
  assign n4363 = ~n4345 ^ n4362;
  assign n4364 = ~n4328 ^ ~n4363;
  assign n4365 = ~n4311 ^ ~n4364;
  assign n4366 = ~n4307 ^ n4365;
  assign n4367 = ~n4303 ^ ~n4366;
  assign n4368 = ~n4224 & n4284;
  assign n4369 = n4220 & ~n4368;
  assign n4370 = n4224 & ~n4284;
  assign n4371 = ~n4369 & ~n4370;
  assign n4372 = n4265 & n4282;
  assign n4373 = ~n4247 & ~n4372;
  assign n4374 = ~n4265 & ~n4282;
  assign n4375 = ~n4373 & ~n4374;
  assign n4376 = n4276 & n4281;
  assign n4377 = n4270 & n4275;
  assign n4378 = ~n4376 & ~n4377;
  assign n4379 = n4238 & ~n4239;
  assign n4380 = ~n4236 & ~n4237;
  assign n4381 = ~n4379 & ~n4380;
  assign n4382 = n4268 & ~n4269;
  assign n4383 = ~n4266 & ~n4267;
  assign n4384 = ~n4382 & ~n4383;
  assign n4385 = ~n4381 ^ ~n4384;
  assign n4386 = n4279 & ~n4280;
  assign n4387 = ~n4277 & ~n4278;
  assign n4388 = ~n4386 & ~n4387;
  assign n4389 = ~n4385 ^ n4388;
  assign n4390 = ~n4378 ^ n4389;
  assign n4391 = ~n4250 & ~n4252;
  assign n4392 = n4249 & ~n4391;
  assign n4393 = n4256 & ~n4257;
  assign n4394 = ~n4254 & ~n4255;
  assign n4395 = ~n4393 & ~n4394;
  assign n4396 = ~n4392 ^ ~n4395;
  assign n4397 = n4261 & ~n4262;
  assign n4398 = ~n4259 & ~n4260;
  assign n4399 = ~n4397 & ~n4398;
  assign n4400 = ~n4396 ^ ~n4399;
  assign n4401 = ~n4390 ^ ~n4400;
  assign n4402 = ~n4375 ^ n4401;
  assign n4403 = n4235 & n4246;
  assign n4404 = n4240 & n4245;
  assign n4405 = ~n4403 & ~n4404;
  assign n4406 = n4273 & ~n4274;
  assign n4407 = ~n4271 & ~n4272;
  assign n4408 = ~n4406 & ~n4407;
  assign n4409 = pi04 & pi47;
  assign n4410 = pi03 & pi48;
  assign n4411 = ~n4409 ^ ~n4410;
  assign n4412 = pi02 & pi49;
  assign n4413 = ~n4411 ^ n4412;
  assign n4414 = ~n4408 ^ n4413;
  assign n4415 = n4243 & ~n4244;
  assign n4416 = ~n4241 & ~n4242;
  assign n4417 = ~n4415 & ~n4416;
  assign n4418 = ~n4414 ^ ~n4417;
  assign n4419 = ~n4405 ^ ~n4418;
  assign n4420 = n4156 & n4167;
  assign n4421 = n4152 & ~n4155;
  assign n4422 = ~n4420 & ~n4421;
  assign n4423 = ~n4419 ^ ~n4422;
  assign n4424 = ~n4402 ^ n4423;
  assign n4425 = n4200 & ~n4211;
  assign n4426 = n4197 & ~n4425;
  assign n4427 = ~n4200 & n4211;
  assign n4428 = ~n4426 & ~n4427;
  assign n4429 = ~n4176 & n4191;
  assign n4430 = ~n4179 & n4190;
  assign n4431 = ~n4429 & ~n4430;
  assign n4432 = n4186 & n4189;
  assign n4433 = n4182 & n4185;
  assign n4434 = ~n4432 & ~n4433;
  assign n4435 = n4163 & n4166;
  assign n4436 = n4159 & n4162;
  assign n4437 = ~n4435 & ~n4436;
  assign n4438 = ~n4434 ^ ~n4437;
  assign n4439 = ~n4253 & n4264;
  assign n4440 = n4258 & n4263;
  assign n4441 = ~n4439 & ~n4440;
  assign n4442 = ~n4438 ^ ~n4441;
  assign n4443 = ~n4431 ^ n4442;
  assign n4444 = ~n4428 ^ n4443;
  assign n4445 = ~n4424 ^ ~n4444;
  assign n4446 = ~n4371 ^ n4445;
  assign n4447 = ~n4367 ^ ~n4446;
  assign n4448 = ~n4299 ^ ~n4447;
  assign po052 = n4295 ^ n4448;
  assign n4450 = ~n4299 & ~n4447;
  assign n4451 = ~n4295 & ~n4450;
  assign n4452 = n4299 & n4447;
  assign n4453 = ~n4451 & ~n4452;
  assign n4454 = ~n4446 & ~n4366;
  assign n4455 = ~n4454 & n4303;
  assign n4456 = n4446 & n4366;
  assign n4457 = ~n4455 & ~n4456;
  assign n4458 = ~n4424 & ~n4444;
  assign n4459 = n4371 & ~n4458;
  assign n4460 = n4424 & n4444;
  assign n4461 = ~n4459 & ~n4460;
  assign n4462 = ~n4311 & ~n4364;
  assign n4463 = ~n4307 & ~n4462;
  assign n4464 = n4311 & n4364;
  assign n4465 = ~n4463 & ~n4464;
  assign n4466 = ~n4405 & ~n4418;
  assign n4467 = ~n4466 & ~n4422;
  assign n4468 = n4405 & n4418;
  assign n4469 = ~n4467 & ~n4468;
  assign n4470 = n4385 & ~n4388;
  assign n4471 = ~n4381 & ~n4384;
  assign n4472 = ~n4470 & ~n4471;
  assign n4473 = pi19 & pi33;
  assign n4474 = pi03 & pi49;
  assign n4475 = ~n4473 ^ ~n4474;
  assign n4476 = pi02 & pi50;
  assign n4477 = ~n4475 ^ n4476;
  assign n4478 = ~n4472 ^ n4477;
  assign n4479 = n4396 & n4399;
  assign n4480 = n4392 & n4395;
  assign n4481 = ~n4479 & ~n4480;
  assign n4482 = ~n4478 ^ n4481;
  assign n4483 = n4414 & n4417;
  assign n4484 = n4408 & ~n4413;
  assign n4485 = ~n4483 & ~n4484;
  assign n4486 = n4339 & ~n4344;
  assign n4487 = ~n4333 & ~n4338;
  assign n4488 = ~n4486 & ~n4487;
  assign n4489 = n4331 & ~n4332;
  assign n4490 = ~n4329 & ~n4330;
  assign n4491 = ~n4489 & ~n4490;
  assign n4492 = pi26 & pi50;
  assign n4493 = ~n4492 ^ ~pi51;
  assign n4494 = n4493 & pi01;
  assign n4495 = pi25 & pi27;
  assign n4496 = ~n4494 ^ n4495;
  assign n4497 = ~n4491 ^ ~n4496;
  assign n4498 = ~n4488 ^ ~n4497;
  assign n4499 = ~n4485 ^ n4498;
  assign n4500 = ~n4482 ^ ~n4499;
  assign n4501 = ~n4469 ^ ~n4500;
  assign n4502 = n4328 & n4363;
  assign n4503 = ~n4345 & n4362;
  assign n4504 = ~n4502 & ~n4503;
  assign n4505 = n4348 & ~n4349;
  assign n4506 = ~n4346 & ~n4347;
  assign n4507 = ~n4505 & ~n4506;
  assign n4508 = n4325 & ~n4326;
  assign n4509 = ~n4323 & ~n4324;
  assign n4510 = ~n4508 & ~n4509;
  assign n4511 = ~n4507 ^ ~n4510;
  assign n4512 = n4411 & ~n4412;
  assign n4513 = ~n4409 & ~n4410;
  assign n4514 = ~n4512 & ~n4513;
  assign n4515 = ~n4511 ^ ~n4514;
  assign n4516 = n4356 & n4361;
  assign n4517 = n4350 & n4355;
  assign n4518 = ~n4516 & ~n4517;
  assign n4519 = ~n4515 ^ ~n4518;
  assign n4520 = n4353 & ~n4354;
  assign n4521 = ~n4351 & ~n4352;
  assign n4522 = ~n4520 & ~n4521;
  assign n4523 = n4336 & ~n4337;
  assign n4524 = ~n4334 & ~n4335;
  assign n4525 = ~n4523 & ~n4524;
  assign n4526 = ~n4522 ^ ~n4525;
  assign n4527 = n4359 & ~n4360;
  assign n4528 = ~n4357 & ~n4358;
  assign n4529 = ~n4527 & ~n4528;
  assign n4530 = ~n4526 ^ ~n4529;
  assign n4531 = ~n4519 ^ ~n4530;
  assign n4532 = ~n4504 ^ ~n4531;
  assign n4533 = n4322 & n4327;
  assign n4534 = n4314 & n4321;
  assign n4535 = ~n4533 & ~n4534;
  assign n4536 = n4252 & pi51;
  assign n4537 = n4315 & pi26;
  assign n4538 = ~n4536 & ~n4537;
  assign n4539 = ~n4492 & pi01;
  assign n4540 = ~n4538 & n4539;
  assign n4541 = ~n4315 & n4319;
  assign n4542 = pi26 & pi51;
  assign n4543 = n4542 & pi00;
  assign n4544 = ~n4541 & n4543;
  assign n4545 = ~n4540 & ~n4544;
  assign n4546 = n4342 & ~n4343;
  assign n4547 = ~n4340 & ~n4341;
  assign n4548 = ~n4546 & ~n4547;
  assign n4549 = pi04 & pi48;
  assign n4550 = ~n2434 ^ ~n4549;
  assign n4551 = pi00 & pi52;
  assign n4552 = ~n4550 ^ n4551;
  assign n4553 = ~n4548 ^ n4552;
  assign n4554 = ~n4545 ^ n4553;
  assign n4555 = ~n4535 ^ ~n4554;
  assign n4556 = n4438 & n4441;
  assign n4557 = ~n4434 & ~n4437;
  assign n4558 = ~n4556 & ~n4557;
  assign n4559 = ~n4555 ^ n4558;
  assign n4560 = ~n4532 ^ ~n4559;
  assign n4561 = ~n4501 ^ n4560;
  assign n4562 = ~n4465 ^ n4561;
  assign n4563 = n4431 & ~n4442;
  assign n4564 = ~n4428 & ~n4563;
  assign n4565 = ~n4431 & n4442;
  assign n4566 = ~n4564 & ~n4565;
  assign n4567 = n4390 & n4400;
  assign n4568 = n4378 & ~n4389;
  assign n4569 = ~n4567 & ~n4568;
  assign n4570 = pi12 & pi40;
  assign n4571 = pi11 & pi41;
  assign n4572 = ~n4570 ^ ~n4571;
  assign n4573 = pi10 & pi42;
  assign n4574 = ~n4572 ^ n4573;
  assign n4575 = pi15 & pi37;
  assign n4576 = pi08 & pi44;
  assign n4577 = ~n4575 ^ ~n4576;
  assign n4578 = pi07 & pi45;
  assign n4579 = ~n4577 ^ n4578;
  assign n4580 = ~n4574 ^ ~n4579;
  assign n4581 = pi16 & pi36;
  assign n4582 = pi06 & pi46;
  assign n4583 = ~n4581 ^ ~n4582;
  assign n4584 = pi05 & pi47;
  assign n4585 = ~n4583 ^ n4584;
  assign n4586 = ~n4580 ^ n4585;
  assign n4587 = pi24 & pi28;
  assign n4588 = pi23 & pi29;
  assign n4589 = ~n4587 ^ ~n4588;
  assign n4590 = pi22 & pi30;
  assign n4591 = ~n4589 ^ n4590;
  assign n4592 = pi14 & pi38;
  assign n4593 = pi13 & pi39;
  assign n4594 = ~n4592 ^ ~n4593;
  assign n4595 = pi09 & pi43;
  assign n4596 = ~n4594 ^ n4595;
  assign n4597 = ~n4591 ^ ~n4596;
  assign n4598 = pi21 & pi31;
  assign n4599 = pi20 & pi32;
  assign n4600 = ~n4598 ^ ~n4599;
  assign n4601 = pi18 & pi34;
  assign n4602 = ~n4600 ^ n4601;
  assign n4603 = ~n4597 ^ ~n4602;
  assign n4604 = ~n4586 ^ n4603;
  assign n4605 = ~n4569 ^ ~n4604;
  assign n4606 = ~n4566 ^ ~n4605;
  assign n4607 = ~n4375 & n4401;
  assign n4608 = ~n4607 & n4423;
  assign n4609 = n4375 & ~n4401;
  assign n4610 = ~n4608 & ~n4609;
  assign n4611 = ~n4606 ^ ~n4610;
  assign n4612 = ~n4562 ^ ~n4611;
  assign n4613 = ~n4461 ^ n4612;
  assign n4614 = ~n4457 ^ n4613;
  assign po053 = n4453 ^ n4614;
  assign n4616 = ~n4457 & n4562;
  assign n4617 = ~n4461 & n4611;
  assign n4618 = n4616 & ~n4617;
  assign n4619 = n4457 & ~n4562;
  assign n4620 = n4461 & ~n4611;
  assign n4621 = ~n4619 & n4620;
  assign n4622 = ~n4618 & ~n4621;
  assign n4623 = ~n4453 & ~n4622;
  assign n4624 = n4616 & n4620;
  assign n4625 = n4619 & n4617;
  assign n4626 = ~n4624 & ~n4625;
  assign n4627 = ~n4623 & n4626;
  assign n4628 = ~n4616 & n4617;
  assign n4629 = n4619 & ~n4620;
  assign n4630 = ~n4628 & ~n4629;
  assign n4631 = n4453 & ~n4630;
  assign n4632 = n4627 & ~n4631;
  assign n4633 = ~n4501 & n4560;
  assign n4634 = ~n4465 & ~n4633;
  assign n4635 = n4501 & ~n4560;
  assign n4636 = ~n4634 & ~n4635;
  assign n4637 = ~n4482 & ~n4499;
  assign n4638 = ~n4469 & ~n4637;
  assign n4639 = n4482 & n4499;
  assign n4640 = ~n4638 & ~n4639;
  assign n4641 = ~n4545 & n4553;
  assign n4642 = n4548 & ~n4552;
  assign n4643 = ~n4641 & ~n4642;
  assign n4644 = n4597 & n4602;
  assign n4645 = n4591 & n4596;
  assign n4646 = ~n4644 & ~n4645;
  assign n4647 = ~n4643 ^ n4646;
  assign n4648 = n4589 & ~n4590;
  assign n4649 = ~n4587 & ~n4588;
  assign n4650 = ~n4648 & ~n4649;
  assign n4651 = n4550 & ~n4551;
  assign n4652 = ~n2434 & ~n4549;
  assign n4653 = ~n4651 & ~n4652;
  assign n4654 = ~n4650 ^ ~n4653;
  assign n4655 = n4475 & ~n4476;
  assign n4656 = ~n4473 & ~n4474;
  assign n4657 = ~n4655 & ~n4656;
  assign n4658 = ~n4654 ^ ~n4657;
  assign n4659 = ~n4647 ^ ~n4658;
  assign n4660 = n4583 & ~n4584;
  assign n4661 = ~n4581 & ~n4582;
  assign n4662 = ~n4660 & ~n4661;
  assign n4663 = n4577 & ~n4578;
  assign n4664 = ~n4575 & ~n4576;
  assign n4665 = ~n4663 & ~n4664;
  assign n4666 = ~n4662 ^ ~n4665;
  assign n4667 = n4600 & ~n4601;
  assign n4668 = ~n4598 & ~n4599;
  assign n4669 = ~n4667 & ~n4668;
  assign n4670 = ~n4666 ^ ~n4669;
  assign n4671 = n4594 & ~n4595;
  assign n4672 = ~n4592 & ~n4593;
  assign n4673 = ~n4671 & ~n4672;
  assign n4674 = n4572 & ~n4573;
  assign n4675 = ~n4570 & ~n4571;
  assign n4676 = ~n4674 & ~n4675;
  assign n4677 = ~n4673 ^ ~n4676;
  assign n4678 = pi01 & pi52;
  assign n4679 = ~n4678 ^ ~pi27;
  assign n4680 = ~n4677 ^ ~n4679;
  assign n4681 = ~n4670 ^ ~n4680;
  assign n4682 = n4580 & ~n4585;
  assign n4683 = ~n4574 & ~n4579;
  assign n4684 = ~n4682 & ~n4683;
  assign n4685 = ~n4681 ^ ~n4684;
  assign n4686 = ~n4659 ^ n4685;
  assign n4687 = ~n4640 ^ n4686;
  assign n4688 = ~n4535 & ~n4554;
  assign n4689 = ~n4688 & ~n4558;
  assign n4690 = n4535 & n4554;
  assign n4691 = ~n4689 & ~n4690;
  assign n4692 = n4586 & ~n4603;
  assign n4693 = n4569 & ~n4692;
  assign n4694 = ~n4586 & n4603;
  assign n4695 = ~n4693 & ~n4694;
  assign n4696 = ~n4495 ^ ~pi51;
  assign n4697 = n4696 & n4492;
  assign n4698 = ~n4491 & ~n4697;
  assign n4699 = ~n4696 & ~n4492;
  assign n4700 = ~n4699 & pi01;
  assign n4701 = ~n4698 & n4700;
  assign n4702 = n4495 & ~pi01;
  assign n4703 = n4491 & n4702;
  assign n4704 = ~n4701 & ~n4703;
  assign n4705 = n4511 & n4514;
  assign n4706 = n4507 & n4510;
  assign n4707 = ~n4705 & ~n4706;
  assign n4708 = ~n4704 ^ ~n4707;
  assign n4709 = n4526 & n4529;
  assign n4710 = n4522 & n4525;
  assign n4711 = ~n4709 & ~n4710;
  assign n4712 = ~n4708 ^ ~n4711;
  assign n4713 = ~n4695 ^ n4712;
  assign n4714 = ~n4691 ^ ~n4713;
  assign n4715 = ~n4687 ^ n4714;
  assign n4716 = n4610 & ~n4605;
  assign n4717 = ~n4716 & n4566;
  assign n4718 = ~n4610 & n4605;
  assign n4719 = ~n4717 & ~n4718;
  assign n4720 = ~n4715 ^ n4719;
  assign n4721 = n4504 & n4531;
  assign n4722 = ~n4721 & ~n4559;
  assign n4723 = ~n4504 & ~n4531;
  assign n4724 = ~n4722 & ~n4723;
  assign n4725 = n4478 & ~n4481;
  assign n4726 = n4472 & ~n4477;
  assign n4727 = ~n4725 & ~n4726;
  assign n4728 = n4495 & pi01;
  assign n4729 = ~n4728 ^ ~pi02;
  assign n4730 = n4729 & pi51;
  assign n4731 = pi03 & pi50;
  assign n4732 = ~n4730 ^ ~n4731;
  assign n4733 = pi18 & pi35;
  assign n4734 = pi17 & pi36;
  assign n4735 = ~n4733 ^ ~n4734;
  assign n4736 = pi04 & pi49;
  assign n4737 = ~n4735 ^ n4736;
  assign n4738 = pi21 & pi32;
  assign n4739 = pi20 & pi33;
  assign n4740 = ~n4738 ^ ~n4739;
  assign n4741 = pi19 & pi34;
  assign n4742 = ~n4740 ^ n4741;
  assign n4743 = ~n4737 ^ ~n4742;
  assign n4744 = ~n4732 ^ ~n4743;
  assign n4745 = ~n4727 ^ n4744;
  assign n4746 = pi15 & pi38;
  assign n4747 = pi07 & pi46;
  assign n4748 = ~n4746 ^ ~n4747;
  assign n4749 = pi06 & pi47;
  assign n4750 = ~n4748 ^ n4749;
  assign n4751 = pi16 & pi37;
  assign n4752 = pi05 & pi48;
  assign n4753 = ~n4751 ^ ~n4752;
  assign n4754 = pi00 & pi53;
  assign n4755 = ~n4753 ^ n4754;
  assign n4756 = ~n4750 ^ ~n4755;
  assign n4757 = pi14 & pi39;
  assign n4758 = pi09 & pi44;
  assign n4759 = ~n4757 ^ ~n4758;
  assign n4760 = pi08 & pi45;
  assign n4761 = ~n4759 ^ n4760;
  assign n4762 = ~n4756 ^ n4761;
  assign n4763 = ~n4745 ^ n4762;
  assign n4764 = ~n4485 & n4498;
  assign n4765 = ~n4488 & ~n4497;
  assign n4766 = ~n4764 & ~n4765;
  assign n4767 = pi13 & pi40;
  assign n4768 = pi12 & pi41;
  assign n4769 = ~n4767 ^ ~n4768;
  assign n4770 = pi10 & pi43;
  assign n4771 = ~n4769 ^ n4770;
  assign n4772 = pi24 & pi29;
  assign n4773 = pi23 & pi30;
  assign n4774 = ~n4772 ^ ~n4773;
  assign n4775 = pi22 & pi31;
  assign n4776 = ~n4774 ^ n4775;
  assign n4777 = ~n4771 ^ ~n4776;
  assign n4778 = pi26 & pi27;
  assign n4779 = pi25 & pi28;
  assign n4780 = ~n4778 ^ ~n4779;
  assign n4781 = pi11 & pi42;
  assign n4782 = ~n4780 ^ n4781;
  assign n4783 = ~n4777 ^ n4782;
  assign n4784 = ~n4766 ^ n4783;
  assign n4785 = n4519 & n4530;
  assign n4786 = n4515 & n4518;
  assign n4787 = ~n4785 & ~n4786;
  assign n4788 = ~n4784 ^ ~n4787;
  assign n4789 = ~n4763 ^ ~n4788;
  assign n4790 = ~n4724 ^ n4789;
  assign n4791 = ~n4720 ^ ~n4790;
  assign n4792 = ~n4636 ^ ~n4791;
  assign po054 = n4632 ^ n4792;
  assign n4794 = ~n4453 & ~n4619;
  assign n4795 = ~n4617 & ~n4792;
  assign n4796 = ~n4616 & ~n4795;
  assign n4797 = ~n4794 & n4796;
  assign n4798 = ~n4618 & n4792;
  assign n4799 = ~n4453 & ~n4798;
  assign n4800 = ~n4619 & ~n4792;
  assign n4801 = ~n4800 & ~n4620;
  assign n4802 = ~n4799 & n4801;
  assign n4803 = ~n4797 & ~n4802;
  assign n4804 = n4720 & n4790;
  assign n4805 = n4636 & ~n4804;
  assign n4806 = ~n4720 & ~n4790;
  assign n4807 = ~n4805 & ~n4806;
  assign n4808 = n4687 & ~n4714;
  assign n4809 = ~n4808 & ~n4719;
  assign n4810 = ~n4687 & n4714;
  assign n4811 = ~n4809 & ~n4810;
  assign n4812 = n4659 & ~n4685;
  assign n4813 = n4640 & ~n4812;
  assign n4814 = ~n4659 & n4685;
  assign n4815 = ~n4813 & ~n4814;
  assign n4816 = ~n4695 & n4712;
  assign n4817 = ~n4691 & ~n4816;
  assign n4818 = n4695 & ~n4712;
  assign n4819 = ~n4817 & ~n4818;
  assign n4820 = n4647 & n4658;
  assign n4821 = ~n4643 & n4646;
  assign n4822 = ~n4820 & ~n4821;
  assign n4823 = n4681 & n4684;
  assign n4824 = ~n4670 & ~n4680;
  assign n4825 = ~n4823 & ~n4824;
  assign n4826 = pi27 & pi52;
  assign n4827 = n4826 & pi01;
  assign n4828 = pi01 & pi53;
  assign n4829 = pi26 & pi28;
  assign n4830 = ~n4828 ^ ~n4829;
  assign n4831 = ~n4827 ^ ~n4830;
  assign n4832 = pi00 & pi54;
  assign n4833 = ~n4831 ^ n4832;
  assign n4834 = pi22 & pi32;
  assign n4835 = pi21 & pi33;
  assign n4836 = ~n4834 ^ ~n4835;
  assign n4837 = pi19 & pi35;
  assign n4838 = ~n4836 ^ n4837;
  assign n4839 = pi25 & pi29;
  assign n4840 = pi24 & pi30;
  assign n4841 = ~n4839 ^ ~n4840;
  assign n4842 = pi23 & pi31;
  assign n4843 = ~n4841 ^ n4842;
  assign n4844 = ~n4838 ^ ~n4843;
  assign n4845 = ~n4833 ^ ~n4844;
  assign n4846 = ~n4825 ^ n4845;
  assign n4847 = ~n4822 ^ ~n4846;
  assign n4848 = ~n4819 ^ ~n4847;
  assign n4849 = ~n4815 ^ n4848;
  assign n4850 = ~n4763 & ~n4788;
  assign n4851 = ~n4724 & ~n4850;
  assign n4852 = n4763 & n4788;
  assign n4853 = ~n4851 & ~n4852;
  assign n4854 = n4745 & ~n4762;
  assign n4855 = n4727 & ~n4744;
  assign n4856 = ~n4854 & ~n4855;
  assign n4857 = n4666 & n4669;
  assign n4858 = n4662 & n4665;
  assign n4859 = ~n4857 & ~n4858;
  assign n4860 = n4677 & n4679;
  assign n4861 = n4673 & n4676;
  assign n4862 = ~n4860 & ~n4861;
  assign n4863 = ~n4859 ^ ~n4862;
  assign n4864 = n4654 & n4657;
  assign n4865 = n4650 & n4653;
  assign n4866 = ~n4864 & ~n4865;
  assign n4867 = ~n4863 ^ n4866;
  assign n4868 = n4756 & ~n4761;
  assign n4869 = ~n4750 & ~n4755;
  assign n4870 = ~n4868 & ~n4869;
  assign n4871 = n4735 & ~n4736;
  assign n4872 = ~n4733 & ~n4734;
  assign n4873 = ~n4871 & ~n4872;
  assign n4874 = n4774 & ~n4775;
  assign n4875 = ~n4772 & ~n4773;
  assign n4876 = ~n4874 & ~n4875;
  assign n4877 = ~n4873 ^ ~n4876;
  assign n4878 = n4740 & ~n4741;
  assign n4879 = ~n4738 & ~n4739;
  assign n4880 = ~n4878 & ~n4879;
  assign n4881 = ~n4877 ^ n4880;
  assign n4882 = ~n4870 ^ ~n4881;
  assign n4883 = n4780 & ~n4781;
  assign n4884 = ~n4778 & ~n4779;
  assign n4885 = ~n4883 & ~n4884;
  assign n4886 = n4748 & ~n4749;
  assign n4887 = ~n4746 & ~n4747;
  assign n4888 = ~n4886 & ~n4887;
  assign n4889 = ~n4885 ^ ~n4888;
  assign n4890 = n4753 & ~n4754;
  assign n4891 = ~n4751 & ~n4752;
  assign n4892 = ~n4890 & ~n4891;
  assign n4893 = ~n4889 ^ ~n4892;
  assign n4894 = ~n4882 ^ n4893;
  assign n4895 = ~n4867 ^ n4894;
  assign n4896 = ~n4856 ^ n4895;
  assign n4897 = n4784 & n4787;
  assign n4898 = n4766 & ~n4783;
  assign n4899 = ~n4897 & ~n4898;
  assign n4900 = n4708 & n4711;
  assign n4901 = n4704 & n4707;
  assign n4902 = ~n4900 & ~n4901;
  assign n4903 = pi14 & pi40;
  assign n4904 = pi10 & pi44;
  assign n4905 = ~n4903 ^ ~n4904;
  assign n4906 = pi09 & pi45;
  assign n4907 = ~n4905 ^ n4906;
  assign n4908 = pi15 & pi39;
  assign n4909 = pi08 & pi46;
  assign n4910 = ~n4908 ^ ~n4909;
  assign n4911 = pi07 & pi47;
  assign n4912 = ~n4910 ^ n4911;
  assign n4913 = ~n4907 ^ ~n4912;
  assign n4914 = pi04 & pi50;
  assign n4915 = pi03 & pi51;
  assign n4916 = ~n4914 ^ ~n4915;
  assign n4917 = pi02 & pi52;
  assign n4918 = ~n4916 ^ n4917;
  assign n4919 = ~n4913 ^ n4918;
  assign n4920 = pi17 & pi37;
  assign n4921 = pi16 & pi38;
  assign n4922 = ~n4920 ^ ~n4921;
  assign n4923 = pi06 & pi48;
  assign n4924 = ~n4922 ^ n4923;
  assign n4925 = pi13 & pi41;
  assign n4926 = pi12 & pi42;
  assign n4927 = ~n4925 ^ ~n4926;
  assign n4928 = pi11 & pi43;
  assign n4929 = ~n4927 ^ n4928;
  assign n4930 = ~n4924 ^ ~n4929;
  assign n4931 = pi20 & pi34;
  assign n4932 = pi18 & pi36;
  assign n4933 = ~n4931 ^ ~n4932;
  assign n4934 = pi05 & pi49;
  assign n4935 = ~n4933 ^ n4934;
  assign n4936 = ~n4930 ^ ~n4935;
  assign n4937 = ~n4919 ^ n4936;
  assign n4938 = ~n4902 ^ n4937;
  assign n4939 = n4732 & n4743;
  assign n4940 = ~n4737 & ~n4742;
  assign n4941 = ~n4939 & ~n4940;
  assign n4942 = n4777 & ~n4782;
  assign n4943 = ~n4771 & ~n4776;
  assign n4944 = ~n4942 & ~n4943;
  assign n4945 = n4769 & ~n4770;
  assign n4946 = ~n4767 & ~n4768;
  assign n4947 = ~n4945 & ~n4946;
  assign n4948 = n4759 & ~n4760;
  assign n4949 = ~n4757 & ~n4758;
  assign n4950 = ~n4948 & ~n4949;
  assign n4951 = ~n4947 ^ ~n4950;
  assign n4952 = n4731 & pi02;
  assign n4953 = ~n4728 & ~n4952;
  assign n4954 = ~n4731 & ~pi02;
  assign n4955 = ~n4954 & pi51;
  assign n4956 = ~n4953 & n4955;
  assign n4957 = ~n4951 ^ n4956;
  assign n4958 = ~n4944 ^ ~n4957;
  assign n4959 = ~n4941 ^ ~n4958;
  assign n4960 = ~n4938 ^ ~n4959;
  assign n4961 = ~n4899 ^ ~n4960;
  assign n4962 = ~n4896 ^ n4961;
  assign n4963 = ~n4853 ^ ~n4962;
  assign n4964 = ~n4849 ^ n4963;
  assign n4965 = ~n4811 ^ n4964;
  assign n4966 = ~n4807 ^ ~n4965;
  assign po055 = ~n4803 ^ n4966;
  assign n4968 = ~n4807 & ~n4965;
  assign n4969 = n4803 & ~n4968;
  assign n4970 = n4807 & n4965;
  assign n4971 = ~n4969 & ~n4970;
  assign n4972 = n4849 & ~n4963;
  assign n4973 = n4811 & ~n4972;
  assign n4974 = ~n4849 & n4963;
  assign n4975 = ~n4973 & ~n4974;
  assign n4976 = n4819 & n4847;
  assign n4977 = n4815 & ~n4976;
  assign n4978 = ~n4819 & ~n4847;
  assign n4979 = ~n4977 & ~n4978;
  assign n4980 = n4919 & ~n4936;
  assign n4981 = ~n4902 & ~n4980;
  assign n4982 = ~n4919 & n4936;
  assign n4983 = ~n4981 & ~n4982;
  assign n4984 = n4889 & n4892;
  assign n4985 = n4885 & n4888;
  assign n4986 = ~n4984 & ~n4985;
  assign n4987 = n4927 & ~n4928;
  assign n4988 = ~n4925 & ~n4926;
  assign n4989 = ~n4987 & ~n4988;
  assign n4990 = pi26 & pi53;
  assign n4991 = n4990 & pi01;
  assign n4992 = ~n4991 & pi28;
  assign n4993 = pi01 & pi54;
  assign n4994 = ~n4992 ^ n4993;
  assign n4995 = ~n4989 ^ n4994;
  assign n4996 = ~n4986 ^ n4995;
  assign n4997 = n4951 & ~n4956;
  assign n4998 = ~n4947 & ~n4950;
  assign n4999 = ~n4997 & ~n4998;
  assign n5000 = ~n4996 ^ ~n4999;
  assign n5001 = n4831 & ~n4832;
  assign n5002 = ~n4827 & ~n4830;
  assign n5003 = ~n5001 & ~n5002;
  assign n5004 = n4910 & ~n4911;
  assign n5005 = ~n4908 & ~n4909;
  assign n5006 = ~n5004 & ~n5005;
  assign n5007 = pi18 & pi37;
  assign n5008 = ~n5007 ^ ~n2506;
  assign n5009 = pi05 & pi50;
  assign n5010 = ~n5008 ^ n5009;
  assign n5011 = ~n5006 ^ n5010;
  assign n5012 = ~n5003 ^ ~n5011;
  assign n5013 = n4916 & ~n4917;
  assign n5014 = ~n4914 & ~n4915;
  assign n5015 = ~n5013 & ~n5014;
  assign n5016 = n4933 & ~n4934;
  assign n5017 = ~n4931 & ~n4932;
  assign n5018 = ~n5016 & ~n5017;
  assign n5019 = ~n5015 ^ ~n5018;
  assign n5020 = n4905 & ~n4906;
  assign n5021 = ~n4903 & ~n4904;
  assign n5022 = ~n5020 & ~n5021;
  assign n5023 = ~n5019 ^ n5022;
  assign n5024 = ~n5012 ^ n5023;
  assign n5025 = n4833 & n4844;
  assign n5026 = n4838 & n4843;
  assign n5027 = ~n5025 & ~n5026;
  assign n5028 = ~n5024 ^ n5027;
  assign n5029 = ~n5000 ^ n5028;
  assign n5030 = ~n4983 ^ n5029;
  assign n5031 = n4859 & n4862;
  assign n5032 = ~n5031 & ~n4866;
  assign n5033 = ~n4859 & ~n4862;
  assign n5034 = ~n5032 & ~n5033;
  assign n5035 = pi22 & pi33;
  assign n5036 = pi21 & pi34;
  assign n5037 = ~n5035 ^ ~n5036;
  assign n5038 = pi20 & pi35;
  assign n5039 = ~n5037 ^ n5038;
  assign n5040 = pi25 & pi30;
  assign n5041 = pi24 & pi31;
  assign n5042 = ~n5040 ^ ~n5041;
  assign n5043 = pi23 & pi32;
  assign n5044 = ~n5042 ^ n5043;
  assign n5045 = ~n5039 ^ ~n5044;
  assign n5046 = pi04 & pi51;
  assign n5047 = pi02 & pi53;
  assign n5048 = ~n5046 ^ ~n5047;
  assign n5049 = pi00 & pi55;
  assign n5050 = ~n5048 ^ n5049;
  assign n5051 = ~n5045 ^ n5050;
  assign n5052 = pi27 & pi28;
  assign n5053 = pi26 & pi29;
  assign n5054 = ~n5052 ^ ~n5053;
  assign n5055 = pi12 & pi43;
  assign n5056 = ~n5054 ^ n5055;
  assign n5057 = pi13 & pi42;
  assign n5058 = pi11 & pi44;
  assign n5059 = ~n5057 ^ ~n5058;
  assign n5060 = pi10 & pi45;
  assign n5061 = ~n5059 ^ n5060;
  assign n5062 = ~n5056 ^ ~n5061;
  assign n5063 = pi16 & pi39;
  assign n5064 = pi08 & pi47;
  assign n5065 = ~n5063 ^ ~n5064;
  assign n5066 = pi07 & pi48;
  assign n5067 = ~n5065 ^ n5066;
  assign n5068 = ~n5062 ^ ~n5067;
  assign n5069 = ~n5051 ^ n5068;
  assign n5070 = ~n5034 ^ n5069;
  assign n5071 = n4836 & ~n4837;
  assign n5072 = ~n4834 & ~n4835;
  assign n5073 = ~n5071 & ~n5072;
  assign n5074 = n4922 & ~n4923;
  assign n5075 = ~n4920 & ~n4921;
  assign n5076 = ~n5074 & ~n5075;
  assign n5077 = ~n5073 ^ ~n5076;
  assign n5078 = n4841 & ~n4842;
  assign n5079 = ~n4839 & ~n4840;
  assign n5080 = ~n5078 & ~n5079;
  assign n5081 = ~n5077 ^ ~n5080;
  assign n5082 = n4930 & n4935;
  assign n5083 = n4924 & n4929;
  assign n5084 = ~n5082 & ~n5083;
  assign n5085 = ~n5081 ^ ~n5084;
  assign n5086 = n4913 & ~n4918;
  assign n5087 = ~n4907 & ~n4912;
  assign n5088 = ~n5086 & ~n5087;
  assign n5089 = ~n5085 ^ n5088;
  assign n5090 = ~n5070 ^ ~n5089;
  assign n5091 = ~n4825 & n4845;
  assign n5092 = ~n4822 & ~n5091;
  assign n5093 = n4825 & ~n4845;
  assign n5094 = ~n5092 & ~n5093;
  assign n5095 = ~n5090 ^ n5094;
  assign n5096 = ~n5030 ^ n5095;
  assign n5097 = ~n4979 ^ n5096;
  assign n5098 = n4896 & ~n4961;
  assign n5099 = n4853 & ~n5098;
  assign n5100 = ~n4896 & n4961;
  assign n5101 = ~n5099 & ~n5100;
  assign n5102 = n4938 & n4959;
  assign n5103 = n4899 & ~n5102;
  assign n5104 = ~n4938 & ~n4959;
  assign n5105 = ~n5103 & ~n5104;
  assign n5106 = n4882 & ~n4893;
  assign n5107 = n4870 & n4881;
  assign n5108 = ~n5106 & ~n5107;
  assign n5109 = n4877 & ~n4880;
  assign n5110 = ~n4873 & ~n4876;
  assign n5111 = ~n5109 & ~n5110;
  assign n5112 = pi17 & pi38;
  assign n5113 = pi06 & pi49;
  assign n5114 = ~n5112 ^ ~n5113;
  assign n5115 = pi03 & pi52;
  assign n5116 = ~n5114 ^ n5115;
  assign n5117 = pi15 & pi40;
  assign n5118 = pi14 & pi41;
  assign n5119 = ~n5117 ^ ~n5118;
  assign n5120 = pi09 & pi46;
  assign n5121 = ~n5119 ^ n5120;
  assign n5122 = ~n5116 ^ ~n5121;
  assign n5123 = ~n5111 ^ n5122;
  assign n5124 = ~n5108 ^ n5123;
  assign n5125 = n4959 & ~n4957;
  assign n5126 = ~n4941 & ~n4944;
  assign n5127 = ~n5125 & ~n5126;
  assign n5128 = ~n5124 ^ n5127;
  assign n5129 = ~n5105 ^ n5128;
  assign n5130 = n4867 & ~n4894;
  assign n5131 = ~n4856 & ~n5130;
  assign n5132 = ~n4867 & n4894;
  assign n5133 = ~n5131 & ~n5132;
  assign n5134 = ~n5129 ^ ~n5133;
  assign n5135 = ~n5101 ^ n5134;
  assign n5136 = ~n5097 ^ ~n5135;
  assign n5137 = ~n4975 ^ n5136;
  assign po056 = n4971 ^ n5137;
  assign n5139 = ~n4975 & n5136;
  assign n5140 = ~n4971 & ~n5139;
  assign n5141 = n4975 & ~n5136;
  assign n5142 = ~n5140 & ~n5141;
  assign n5143 = ~n5101 & n5134;
  assign n5144 = ~n5097 & ~n5143;
  assign n5145 = n5101 & ~n5134;
  assign n5146 = ~n5144 & ~n5145;
  assign n5147 = n5030 & ~n5095;
  assign n5148 = ~n4979 & ~n5147;
  assign n5149 = ~n5030 & n5095;
  assign n5150 = ~n5148 & ~n5149;
  assign n5151 = ~n5105 & n5128;
  assign n5152 = ~n5151 & ~n5133;
  assign n5153 = n5105 & ~n5128;
  assign n5154 = ~n5152 & ~n5153;
  assign n5155 = n5108 & ~n5123;
  assign n5156 = ~n5155 & n5127;
  assign n5157 = ~n5108 & n5123;
  assign n5158 = ~n5156 & ~n5157;
  assign n5159 = n5114 & ~n5115;
  assign n5160 = ~n5112 & ~n5113;
  assign n5161 = ~n5159 & ~n5160;
  assign n5162 = n5037 & ~n5038;
  assign n5163 = ~n5035 & ~n5036;
  assign n5164 = ~n5162 & ~n5163;
  assign n5165 = ~n5161 ^ ~n5164;
  assign n5166 = n5042 & ~n5043;
  assign n5167 = ~n5040 & ~n5041;
  assign n5168 = ~n5166 & ~n5167;
  assign n5169 = ~n5165 ^ n5168;
  assign n5170 = n5059 & ~n5060;
  assign n5171 = ~n5057 & ~n5058;
  assign n5172 = ~n5170 & ~n5171;
  assign n5173 = n5054 & ~n5055;
  assign n5174 = ~n5052 & ~n5053;
  assign n5175 = ~n5173 & ~n5174;
  assign n5176 = ~n5172 ^ ~n5175;
  assign n5177 = pi01 & pi55;
  assign n5178 = pi27 & pi29;
  assign n5179 = ~n5177 ^ ~n5178;
  assign n5180 = ~n5176 ^ ~n5179;
  assign n5181 = ~n5169 ^ n5180;
  assign n5182 = n5062 & n5067;
  assign n5183 = n5056 & n5061;
  assign n5184 = ~n5182 & ~n5183;
  assign n5185 = ~n5181 ^ ~n5184;
  assign n5186 = ~n1558 & ~pi02;
  assign n5187 = ~n5186 & pi54;
  assign n5188 = n1558 & pi02;
  assign n5189 = n5187 & ~n5188;
  assign n5190 = pi00 & pi56;
  assign n5191 = ~n5189 ^ ~n5190;
  assign n5192 = pi19 & pi37;
  assign n5193 = pi04 & pi52;
  assign n5194 = ~n5192 ^ ~n5193;
  assign n5195 = pi03 & pi53;
  assign n5196 = ~n5194 ^ n5195;
  assign n5197 = ~n5191 ^ n5196;
  assign n5198 = n5065 & ~n5066;
  assign n5199 = ~n5063 & ~n5064;
  assign n5200 = ~n5198 & ~n5199;
  assign n5201 = ~n5197 ^ ~n5200;
  assign n5202 = pi14 & pi42;
  assign n5203 = pi10 & pi46;
  assign n5204 = ~n5202 ^ ~n5203;
  assign n5205 = pi09 & pi47;
  assign n5206 = ~n5204 ^ n5205;
  assign n5207 = pi26 & pi30;
  assign n5208 = pi25 & pi31;
  assign n5209 = ~n5207 ^ ~n5208;
  assign n5210 = pi24 & pi32;
  assign n5211 = ~n5209 ^ n5210;
  assign n5212 = ~n5206 ^ ~n5211;
  assign n5213 = pi23 & pi33;
  assign n5214 = pi22 & pi34;
  assign n5215 = ~n5213 ^ ~n5214;
  assign n5216 = pi20 & pi36;
  assign n5217 = ~n5215 ^ n5216;
  assign n5218 = ~n5212 ^ n5217;
  assign n5219 = pi13 & pi43;
  assign n5220 = pi12 & pi44;
  assign n5221 = ~n5219 ^ ~n5220;
  assign n5222 = pi11 & pi45;
  assign n5223 = ~n5221 ^ n5222;
  assign n5224 = pi16 & pi40;
  assign n5225 = pi15 & pi41;
  assign n5226 = ~n5224 ^ ~n5225;
  assign n5227 = pi08 & pi48;
  assign n5228 = ~n5226 ^ n5227;
  assign n5229 = ~n5223 ^ ~n5228;
  assign n5230 = pi17 & pi39;
  assign n5231 = pi07 & pi49;
  assign n5232 = ~n5230 ^ ~n5231;
  assign n5233 = pi06 & pi50;
  assign n5234 = ~n5232 ^ n5233;
  assign n5235 = ~n5229 ^ ~n5234;
  assign n5236 = ~n5218 ^ n5235;
  assign n5237 = ~n5201 ^ ~n5236;
  assign n5238 = ~n5185 ^ ~n5237;
  assign n5239 = ~n5158 ^ n5238;
  assign n5240 = n4996 & n4999;
  assign n5241 = ~n4986 & n4995;
  assign n5242 = ~n5240 & ~n5241;
  assign n5243 = ~n5111 & n5122;
  assign n5244 = n5116 & n5121;
  assign n5245 = ~n5243 & ~n5244;
  assign n5246 = n5008 & ~n5009;
  assign n5247 = ~n5007 & ~n2506;
  assign n5248 = ~n5246 & ~n5247;
  assign n5249 = n5048 & ~n5049;
  assign n5250 = ~n5046 & ~n5047;
  assign n5251 = ~n5249 & ~n5250;
  assign n5252 = ~n5248 ^ ~n5251;
  assign n5253 = n5119 & ~n5120;
  assign n5254 = ~n5117 & ~n5118;
  assign n5255 = ~n5253 & ~n5254;
  assign n5256 = ~n5252 ^ ~n5255;
  assign n5257 = ~n5245 ^ ~n5256;
  assign n5258 = ~n5242 ^ n5257;
  assign n5259 = n5003 & n5011;
  assign n5260 = n5006 & ~n5010;
  assign n5261 = ~n5259 & ~n5260;
  assign n5262 = n5077 & n5080;
  assign n5263 = n5073 & n5076;
  assign n5264 = ~n5262 & ~n5263;
  assign n5265 = ~n5261 ^ ~n5264;
  assign n5266 = n5045 & ~n5050;
  assign n5267 = ~n5039 & ~n5044;
  assign n5268 = ~n5266 & ~n5267;
  assign n5269 = ~n5265 ^ ~n5268;
  assign n5270 = ~n5258 ^ n5269;
  assign n5271 = n5051 & ~n5068;
  assign n5272 = n5034 & ~n5271;
  assign n5273 = ~n5051 & n5068;
  assign n5274 = ~n5272 & ~n5273;
  assign n5275 = ~n5270 ^ ~n5274;
  assign n5276 = ~n5239 ^ n5275;
  assign n5277 = ~n5154 ^ ~n5276;
  assign n5278 = ~n5000 & n5028;
  assign n5279 = n4983 & ~n5278;
  assign n5280 = n5000 & ~n5028;
  assign n5281 = ~n5279 & ~n5280;
  assign n5282 = n4989 & pi54;
  assign n5283 = pi28 & pi53;
  assign n5284 = n5283 & pi26;
  assign n5285 = ~n5282 & ~n5284;
  assign n5286 = pi28 & pi54;
  assign n5287 = ~n5286 & pi01;
  assign n5288 = ~n5285 & n5287;
  assign n5289 = ~n4990 & n4993;
  assign n5290 = ~n5289 & pi28;
  assign n5291 = n4989 & n5290;
  assign n5292 = ~n5288 & ~n5291;
  assign n5293 = pi21 & pi35;
  assign n5294 = pi18 & pi38;
  assign n5295 = ~n5293 ^ ~n5294;
  assign n5296 = pi05 & pi51;
  assign n5297 = ~n5295 ^ n5296;
  assign n5298 = ~n5292 ^ ~n5297;
  assign n5299 = n5019 & ~n5022;
  assign n5300 = ~n5015 & ~n5018;
  assign n5301 = ~n5299 & ~n5300;
  assign n5302 = ~n5298 ^ n5301;
  assign n5303 = n5085 & ~n5088;
  assign n5304 = n5081 & n5084;
  assign n5305 = ~n5303 & ~n5304;
  assign n5306 = n5024 & ~n5027;
  assign n5307 = ~n5012 & n5023;
  assign n5308 = ~n5306 & ~n5307;
  assign n5309 = ~n5305 ^ n5308;
  assign n5310 = ~n5302 ^ n5309;
  assign n5311 = ~n5281 ^ n5310;
  assign n5312 = ~n5070 & ~n5089;
  assign n5313 = ~n5312 & ~n5094;
  assign n5314 = n5070 & n5089;
  assign n5315 = ~n5313 & ~n5314;
  assign n5316 = ~n5311 ^ n5315;
  assign n5317 = ~n5277 ^ ~n5316;
  assign n5318 = ~n5150 ^ ~n5317;
  assign n5319 = ~n5146 ^ n5318;
  assign po057 = ~n5142 ^ ~n5319;
  assign n5321 = n5146 & ~n5318;
  assign n5322 = ~n5142 & ~n5321;
  assign n5323 = ~n5146 & n5318;
  assign n5324 = ~n5322 & ~n5323;
  assign n5325 = ~n5277 & ~n5316;
  assign n5326 = ~n5150 & ~n5325;
  assign n5327 = n5277 & n5316;
  assign n5328 = ~n5326 & ~n5327;
  assign n5329 = n5239 & ~n5275;
  assign n5330 = n5154 & ~n5329;
  assign n5331 = ~n5239 & n5275;
  assign n5332 = ~n5330 & ~n5331;
  assign n5333 = n5281 & ~n5310;
  assign n5334 = ~n5333 & ~n5315;
  assign n5335 = ~n5281 & n5310;
  assign n5336 = ~n5334 & ~n5335;
  assign n5337 = ~n5305 & n5308;
  assign n5338 = n5302 & ~n5337;
  assign n5339 = n5305 & ~n5308;
  assign n5340 = ~n5338 & ~n5339;
  assign n5341 = n5265 & n5268;
  assign n5342 = n5261 & n5264;
  assign n5343 = ~n5341 & ~n5342;
  assign n5344 = pi04 & pi53;
  assign n5345 = pi03 & pi54;
  assign n5346 = ~n5344 ^ ~n5345;
  assign n5347 = pi02 & pi55;
  assign n5348 = ~n5346 ^ n5347;
  assign n5349 = pi19 & pi38;
  assign n5350 = ~n2674 ^ ~n5349;
  assign n5351 = pi05 & pi52;
  assign n5352 = ~n5350 ^ n5351;
  assign n5353 = ~n5348 ^ ~n5352;
  assign n5354 = pi15 & pi42;
  assign n5355 = pi10 & pi47;
  assign n5356 = ~n5354 ^ ~n5355;
  assign n5357 = pi09 & pi48;
  assign n5358 = ~n5356 ^ n5357;
  assign n5359 = ~n5353 ^ n5358;
  assign n5360 = pi14 & pi43;
  assign n5361 = pi13 & pi44;
  assign n5362 = ~n5360 ^ ~n5361;
  assign n5363 = pi11 & pi46;
  assign n5364 = ~n5362 ^ n5363;
  assign n5365 = pi18 & pi39;
  assign n5366 = pi17 & pi40;
  assign n5367 = ~n5365 ^ ~n5366;
  assign n5368 = pi06 & pi51;
  assign n5369 = ~n5367 ^ n5368;
  assign n5370 = ~n5364 ^ ~n5369;
  assign n5371 = pi28 & pi29;
  assign n5372 = pi27 & pi30;
  assign n5373 = ~n5371 ^ ~n5372;
  assign n5374 = pi12 & pi45;
  assign n5375 = ~n5373 ^ n5374;
  assign n5376 = ~n5370 ^ ~n5375;
  assign n5377 = ~n5359 ^ n5376;
  assign n5378 = ~n5343 ^ n5377;
  assign n5379 = ~n5340 ^ n5378;
  assign n5380 = n5298 & ~n5301;
  assign n5381 = n5292 & n5297;
  assign n5382 = ~n5380 & ~n5381;
  assign n5383 = pi26 & pi31;
  assign n5384 = pi25 & pi32;
  assign n5385 = ~n5383 ^ ~n5384;
  assign n5386 = pi24 & pi33;
  assign n5387 = ~n5385 ^ n5386;
  assign n5388 = pi23 & pi34;
  assign n5389 = pi22 & pi35;
  assign n5390 = ~n5388 ^ ~n5389;
  assign n5391 = pi21 & pi36;
  assign n5392 = ~n5390 ^ n5391;
  assign n5393 = ~n5387 ^ ~n5392;
  assign n5394 = pi16 & pi41;
  assign n5395 = pi08 & pi49;
  assign n5396 = ~n5394 ^ ~n5395;
  assign n5397 = pi07 & pi50;
  assign n5398 = ~n5396 ^ n5397;
  assign n5399 = ~n5393 ^ n5398;
  assign n5400 = ~n5382 ^ ~n5399;
  assign n5401 = n5295 & ~n5296;
  assign n5402 = ~n5293 & ~n5294;
  assign n5403 = ~n5401 & ~n5402;
  assign n5404 = n5221 & ~n5222;
  assign n5405 = ~n5219 & ~n5220;
  assign n5406 = ~n5404 & ~n5405;
  assign n5407 = ~n5403 ^ ~n5406;
  assign n5408 = n5204 & ~n5205;
  assign n5409 = ~n5202 & ~n5203;
  assign n5410 = ~n5408 & ~n5409;
  assign n5411 = ~n5407 ^ ~n5410;
  assign n5412 = ~n5400 ^ n5411;
  assign n5413 = ~n5379 ^ ~n5412;
  assign n5414 = n5201 & n5236;
  assign n5415 = n5218 & ~n5235;
  assign n5416 = ~n5414 & ~n5415;
  assign n5417 = n5209 & ~n5210;
  assign n5418 = ~n5207 & ~n5208;
  assign n5419 = ~n5417 & ~n5418;
  assign n5420 = n5226 & ~n5227;
  assign n5421 = ~n5224 & ~n5225;
  assign n5422 = ~n5420 & ~n5421;
  assign n5423 = ~n5419 ^ ~n5422;
  assign n5424 = n5232 & ~n5233;
  assign n5425 = ~n5230 & ~n5231;
  assign n5426 = ~n5424 & ~n5425;
  assign n5427 = ~n5423 ^ n5426;
  assign n5428 = n5194 & ~n5195;
  assign n5429 = ~n5192 & ~n5193;
  assign n5430 = ~n5428 & ~n5429;
  assign n5431 = n5215 & ~n5216;
  assign n5432 = ~n5213 & ~n5214;
  assign n5433 = ~n5431 & ~n5432;
  assign n5434 = ~n5430 ^ ~n5433;
  assign n5435 = ~n5188 & ~n5190;
  assign n5436 = n5187 & ~n5435;
  assign n5437 = ~n5434 ^ n5436;
  assign n5438 = ~n5427 ^ ~n5437;
  assign n5439 = n5229 & n5234;
  assign n5440 = n5223 & n5228;
  assign n5441 = ~n5439 & ~n5440;
  assign n5442 = ~n5438 ^ ~n5441;
  assign n5443 = ~n5416 ^ n5442;
  assign n5444 = n5197 & n5200;
  assign n5445 = n5191 & ~n5196;
  assign n5446 = ~n5444 & ~n5445;
  assign n5447 = n5176 & n5179;
  assign n5448 = n5172 & n5175;
  assign n5449 = ~n5447 & ~n5448;
  assign n5450 = ~n5446 ^ ~n5449;
  assign n5451 = n5212 & ~n5217;
  assign n5452 = ~n5206 & ~n5211;
  assign n5453 = ~n5451 & ~n5452;
  assign n5454 = ~n5450 ^ n5453;
  assign n5455 = ~n5443 ^ ~n5454;
  assign n5456 = ~n5413 ^ n5455;
  assign n5457 = ~n5336 ^ ~n5456;
  assign n5458 = ~n5332 ^ ~n5457;
  assign n5459 = ~n5258 & n5269;
  assign n5460 = ~n5459 & n5274;
  assign n5461 = n5258 & ~n5269;
  assign n5462 = ~n5460 & ~n5461;
  assign n5463 = n5245 & n5256;
  assign n5464 = n5242 & ~n5463;
  assign n5465 = ~n5245 & ~n5256;
  assign n5466 = ~n5464 & ~n5465;
  assign n5467 = n5181 & n5184;
  assign n5468 = ~n5169 & n5180;
  assign n5469 = ~n5467 & ~n5468;
  assign n5470 = n5165 & ~n5168;
  assign n5471 = ~n5161 & ~n5164;
  assign n5472 = ~n5470 & ~n5471;
  assign n5473 = n5252 & n5255;
  assign n5474 = n5248 & n5251;
  assign n5475 = ~n5473 & ~n5474;
  assign n5476 = ~n5472 ^ n5475;
  assign n5477 = pi27 & pi55;
  assign n5478 = n5477 & pi01;
  assign n5479 = ~n5478 & pi29;
  assign n5480 = pi00 & pi57;
  assign n5481 = pi01 & pi56;
  assign n5482 = ~n5480 ^ n5481;
  assign n5483 = ~n5479 ^ n5482;
  assign n5484 = ~n5476 ^ n5483;
  assign n5485 = ~n5469 ^ ~n5484;
  assign n5486 = ~n5466 ^ n5485;
  assign n5487 = ~n5462 ^ ~n5486;
  assign n5488 = n5185 & n5237;
  assign n5489 = ~n5158 & ~n5488;
  assign n5490 = ~n5185 & ~n5237;
  assign n5491 = ~n5489 & ~n5490;
  assign n5492 = ~n5487 ^ n5491;
  assign n5493 = ~n5458 ^ n5492;
  assign n5494 = ~n5328 ^ ~n5493;
  assign po058 = ~n5324 ^ n5494;
  assign n5496 = ~n5457 & ~n5492;
  assign n5497 = ~n5324 & ~n5496;
  assign n5498 = ~n5328 & ~n5332;
  assign n5499 = n5457 & n5492;
  assign n5500 = ~n5498 & n5499;
  assign n5501 = n5328 & n5332;
  assign n5502 = ~n5500 & ~n5501;
  assign n5503 = n5497 & ~n5502;
  assign n5504 = ~n5501 & n5496;
  assign n5505 = n5498 & ~n5499;
  assign n5506 = ~n5504 & ~n5505;
  assign n5507 = n5324 & ~n5506;
  assign n5508 = n5501 & n5499;
  assign n5509 = n5496 & ~n5332;
  assign n5510 = ~n5328 & n5509;
  assign n5511 = ~n5508 & ~n5510;
  assign n5512 = ~n5507 & n5511;
  assign n5513 = ~n5503 & n5512;
  assign n5514 = n5462 & n5486;
  assign n5515 = ~n5514 & n5491;
  assign n5516 = ~n5462 & ~n5486;
  assign n5517 = ~n5515 & ~n5516;
  assign n5518 = n5450 & ~n5453;
  assign n5519 = ~n5446 & ~n5449;
  assign n5520 = ~n5518 & ~n5519;
  assign n5521 = pi18 & pi40;
  assign n5522 = pi08 & pi50;
  assign n5523 = ~n5521 ^ ~n5522;
  assign n5524 = pi07 & pi51;
  assign n5525 = ~n5523 ^ n5524;
  assign n5526 = pi27 & pi31;
  assign n5527 = pi26 & pi32;
  assign n5528 = ~n5526 ^ ~n5527;
  assign n5529 = pi25 & pi33;
  assign n5530 = ~n5528 ^ n5529;
  assign n5531 = ~n5525 ^ ~n5530;
  assign n5532 = pi24 & pi34;
  assign n5533 = pi23 & pi35;
  assign n5534 = ~n5532 ^ ~n5533;
  assign n5535 = pi22 & pi36;
  assign n5536 = ~n5534 ^ n5535;
  assign n5537 = ~n5531 ^ ~n5536;
  assign n5538 = ~n5520 ^ ~n5537;
  assign n5539 = pi17 & pi41;
  assign n5540 = pi16 & pi42;
  assign n5541 = ~n5539 ^ ~n5540;
  assign n5542 = pi09 & pi49;
  assign n5543 = ~n5541 ^ n5542;
  assign n5544 = pi21 & pi37;
  assign n5545 = ~n2744 ^ ~n5544;
  assign n5546 = pi05 & pi53;
  assign n5547 = ~n5545 ^ n5546;
  assign n5548 = ~n5543 ^ ~n5547;
  assign n5549 = pi04 & pi54;
  assign n5550 = pi02 & pi56;
  assign n5551 = ~n5549 ^ ~n5550;
  assign n5552 = pi00 & pi58;
  assign n5553 = ~n5551 ^ n5552;
  assign n5554 = ~n5548 ^ n5553;
  assign n5555 = ~n5538 ^ ~n5554;
  assign n5556 = n5484 & n5472;
  assign n5557 = ~n5475 & n5483;
  assign n5558 = ~n5556 & ~n5557;
  assign n5559 = n1641 & n5477;
  assign n5560 = ~n5559 & ~n5481;
  assign n5561 = n5480 & ~pi29;
  assign n5562 = ~n5561 & pi56;
  assign n5563 = ~n5560 & ~n5562;
  assign n5564 = ~n5477 & n5481;
  assign n5565 = pi29 & pi57;
  assign n5566 = n5565 & pi00;
  assign n5567 = ~n5564 & n5566;
  assign n5568 = ~n5563 & ~n5567;
  assign n5569 = n5396 & ~n5397;
  assign n5570 = ~n5394 & ~n5395;
  assign n5571 = ~n5569 & ~n5570;
  assign n5572 = n5367 & ~n5368;
  assign n5573 = ~n5365 & ~n5366;
  assign n5574 = ~n5572 & ~n5573;
  assign n5575 = ~n5571 ^ ~n5574;
  assign n5576 = ~n5568 ^ n5575;
  assign n5577 = pi19 & pi39;
  assign n5578 = pi06 & pi52;
  assign n5579 = ~n5577 ^ ~n5578;
  assign n5580 = pi03 & pi55;
  assign n5581 = ~n5579 ^ n5580;
  assign n5582 = pi15 & pi43;
  assign n5583 = pi11 & pi47;
  assign n5584 = ~n5582 ^ ~n5583;
  assign n5585 = pi10 & pi48;
  assign n5586 = ~n5584 ^ n5585;
  assign n5587 = ~n5581 ^ ~n5586;
  assign n5588 = pi14 & pi44;
  assign n5589 = pi13 & pi45;
  assign n5590 = ~n5588 ^ ~n5589;
  assign n5591 = pi12 & pi46;
  assign n5592 = ~n5590 ^ n5591;
  assign n5593 = ~n5587 ^ ~n5592;
  assign n5594 = ~n5576 ^ n5593;
  assign n5595 = ~n5558 ^ n5594;
  assign n5596 = ~n5555 ^ ~n5595;
  assign n5597 = ~n5469 & ~n5484;
  assign n5598 = ~n5466 & ~n5597;
  assign n5599 = n5469 & n5484;
  assign n5600 = ~n5598 & ~n5599;
  assign n5601 = ~n5596 ^ n5600;
  assign n5602 = n5359 & ~n5376;
  assign n5603 = ~n5343 & ~n5602;
  assign n5604 = ~n5359 & n5376;
  assign n5605 = ~n5603 & ~n5604;
  assign n5606 = n5353 & ~n5358;
  assign n5607 = ~n5348 & ~n5352;
  assign n5608 = ~n5606 & ~n5607;
  assign n5609 = n5373 & ~n5374;
  assign n5610 = ~n5371 & ~n5372;
  assign n5611 = ~n5609 & ~n5610;
  assign n5612 = pi29 & pi56;
  assign n5613 = ~n5612 ^ ~pi57;
  assign n5614 = n5613 & pi01;
  assign n5615 = pi28 & pi30;
  assign n5616 = ~n5614 ^ n5615;
  assign n5617 = ~n5611 ^ n5616;
  assign n5618 = ~n5608 ^ n5617;
  assign n5619 = n5370 & n5375;
  assign n5620 = n5364 & n5369;
  assign n5621 = ~n5619 & ~n5620;
  assign n5622 = ~n5618 ^ ~n5621;
  assign n5623 = n5346 & ~n5347;
  assign n5624 = ~n5344 & ~n5345;
  assign n5625 = ~n5623 & ~n5624;
  assign n5626 = n5362 & ~n5363;
  assign n5627 = ~n5360 & ~n5361;
  assign n5628 = ~n5626 & ~n5627;
  assign n5629 = ~n5625 ^ ~n5628;
  assign n5630 = n5350 & ~n5351;
  assign n5631 = ~n2674 & ~n5349;
  assign n5632 = ~n5630 & ~n5631;
  assign n5633 = ~n5629 ^ ~n5632;
  assign n5634 = n5393 & ~n5398;
  assign n5635 = ~n5387 & ~n5392;
  assign n5636 = ~n5634 & ~n5635;
  assign n5637 = ~n5633 ^ n5636;
  assign n5638 = n5390 & ~n5391;
  assign n5639 = ~n5388 & ~n5389;
  assign n5640 = ~n5638 & ~n5639;
  assign n5641 = n5385 & ~n5386;
  assign n5642 = ~n5383 & ~n5384;
  assign n5643 = ~n5641 & ~n5642;
  assign n5644 = ~n5640 ^ ~n5643;
  assign n5645 = n5356 & ~n5357;
  assign n5646 = ~n5354 & ~n5355;
  assign n5647 = ~n5645 & ~n5646;
  assign n5648 = ~n5644 ^ n5647;
  assign n5649 = ~n5637 ^ n5648;
  assign n5650 = ~n5622 ^ ~n5649;
  assign n5651 = ~n5605 ^ n5650;
  assign n5652 = ~n5601 ^ ~n5651;
  assign n5653 = ~n5517 ^ ~n5652;
  assign n5654 = n5400 & ~n5411;
  assign n5655 = ~n5382 & ~n5399;
  assign n5656 = ~n5654 & ~n5655;
  assign n5657 = n5438 & n5441;
  assign n5658 = ~n5427 & ~n5437;
  assign n5659 = ~n5657 & ~n5658;
  assign n5660 = n5434 & ~n5436;
  assign n5661 = ~n5430 & ~n5433;
  assign n5662 = ~n5660 & ~n5661;
  assign n5663 = n5423 & ~n5426;
  assign n5664 = ~n5419 & ~n5422;
  assign n5665 = ~n5663 & ~n5664;
  assign n5666 = ~n5662 ^ ~n5665;
  assign n5667 = n5407 & n5410;
  assign n5668 = n5403 & n5406;
  assign n5669 = ~n5667 & ~n5668;
  assign n5670 = ~n5666 ^ ~n5669;
  assign n5671 = ~n5659 ^ ~n5670;
  assign n5672 = ~n5656 ^ ~n5671;
  assign n5673 = n5443 & n5454;
  assign n5674 = ~n5416 & n5442;
  assign n5675 = ~n5673 & ~n5674;
  assign n5676 = ~n5672 ^ n5675;
  assign n5677 = n5340 & ~n5378;
  assign n5678 = ~n5677 & n5412;
  assign n5679 = ~n5340 & n5378;
  assign n5680 = ~n5678 & ~n5679;
  assign n5681 = ~n5676 ^ ~n5680;
  assign n5682 = ~n5653 ^ n5681;
  assign n5683 = n5413 & ~n5455;
  assign n5684 = ~n5336 & ~n5683;
  assign n5685 = ~n5413 & n5455;
  assign n5686 = ~n5684 & ~n5685;
  assign n5687 = ~n5682 ^ n5686;
  assign po059 = n5513 ^ n5687;
  assign n5689 = ~n5500 & n5687;
  assign n5690 = ~n5324 & ~n5689;
  assign n5691 = ~n5687 & ~n5496;
  assign n5692 = ~n5501 & ~n5691;
  assign n5693 = ~n5690 & n5692;
  assign n5694 = ~n5498 & ~n5687;
  assign n5695 = ~n5694 & ~n5499;
  assign n5696 = ~n5497 & n5695;
  assign n5697 = ~n5693 & ~n5696;
  assign n5698 = n5653 & ~n5681;
  assign n5699 = ~n5698 & ~n5686;
  assign n5700 = ~n5653 & n5681;
  assign n5701 = ~n5699 & ~n5700;
  assign n5702 = ~n5659 & ~n5670;
  assign n5703 = ~n5656 & ~n5702;
  assign n5704 = n5659 & n5670;
  assign n5705 = ~n5703 & ~n5704;
  assign n5706 = n5618 & n5621;
  assign n5707 = ~n5608 & n5617;
  assign n5708 = ~n5706 & ~n5707;
  assign n5709 = pi14 & pi45;
  assign n5710 = pi12 & pi47;
  assign n5711 = ~n5709 ^ ~n5710;
  assign n5712 = pi11 & pi48;
  assign n5713 = ~n5711 ^ n5712;
  assign n5714 = pi17 & pi42;
  assign n5715 = pi16 & pi43;
  assign n5716 = ~n5714 ^ ~n5715;
  assign n5717 = pi08 & pi51;
  assign n5718 = ~n5716 ^ n5717;
  assign n5719 = ~n5713 ^ ~n5718;
  assign n5720 = pi29 & pi30;
  assign n5721 = pi28 & pi31;
  assign n5722 = ~n5720 ^ ~n5721;
  assign n5723 = pi13 & pi46;
  assign n5724 = ~n5722 ^ n5723;
  assign n5725 = ~n5719 ^ ~n5724;
  assign n5726 = ~n5708 ^ ~n5725;
  assign n5727 = n5528 & ~n5529;
  assign n5728 = ~n5526 & ~n5527;
  assign n5729 = ~n5727 & ~n5728;
  assign n5730 = pi19 & pi40;
  assign n5731 = pi05 & pi54;
  assign n5732 = ~n5730 ^ ~n5731;
  assign n5733 = pi04 & pi55;
  assign n5734 = ~n5732 ^ n5733;
  assign n5735 = ~n5729 ^ n5734;
  assign n5736 = n1769 & pi28;
  assign n5737 = ~n5736 ^ ~pi02;
  assign n5738 = n5737 & pi57;
  assign n5739 = pi03 & pi56;
  assign n5740 = ~n5738 ^ ~n5739;
  assign n5741 = ~n5735 ^ ~n5740;
  assign n5742 = ~n5726 ^ n5741;
  assign n5743 = n5666 & n5669;
  assign n5744 = ~n5662 & ~n5665;
  assign n5745 = ~n5743 & ~n5744;
  assign n5746 = ~n5615 ^ ~pi57;
  assign n5747 = n5746 & n5612;
  assign n5748 = ~n5611 & ~n5747;
  assign n5749 = ~n5746 & ~n5612;
  assign n5750 = ~n5749 & pi01;
  assign n5751 = ~n5748 & n5750;
  assign n5752 = n5615 & ~pi01;
  assign n5753 = n5611 & n5752;
  assign n5754 = ~n5751 & ~n5753;
  assign n5755 = pi18 & pi41;
  assign n5756 = pi07 & pi52;
  assign n5757 = ~n5755 ^ ~n5756;
  assign n5758 = pi06 & pi53;
  assign n5759 = ~n5757 ^ n5758;
  assign n5760 = pi15 & pi44;
  assign n5761 = pi10 & pi49;
  assign n5762 = ~n5760 ^ ~n5761;
  assign n5763 = pi09 & pi50;
  assign n5764 = ~n5762 ^ n5763;
  assign n5765 = ~n5759 ^ ~n5764;
  assign n5766 = ~n5754 ^ n5765;
  assign n5767 = pi22 & pi37;
  assign n5768 = pi21 & pi38;
  assign n5769 = ~n5767 ^ ~n5768;
  assign n5770 = pi20 & pi39;
  assign n5771 = ~n5769 ^ n5770;
  assign n5772 = pi27 & pi32;
  assign n5773 = pi26 & pi33;
  assign n5774 = ~n5772 ^ ~n5773;
  assign n5775 = pi00 & pi59;
  assign n5776 = ~n5774 ^ n5775;
  assign n5777 = ~n5771 ^ ~n5776;
  assign n5778 = pi25 & pi34;
  assign n5779 = pi24 & pi35;
  assign n5780 = ~n5778 ^ ~n5779;
  assign n5781 = pi23 & pi36;
  assign n5782 = ~n5780 ^ n5781;
  assign n5783 = ~n5777 ^ ~n5782;
  assign n5784 = ~n5766 ^ n5783;
  assign n5785 = ~n5745 ^ n5784;
  assign n5786 = ~n5742 ^ ~n5785;
  assign n5787 = ~n5705 ^ n5786;
  assign n5788 = n5538 & n5554;
  assign n5789 = ~n5520 & ~n5537;
  assign n5790 = ~n5788 & ~n5789;
  assign n5791 = n5531 & n5536;
  assign n5792 = n5525 & n5530;
  assign n5793 = ~n5791 & ~n5792;
  assign n5794 = n5548 & ~n5553;
  assign n5795 = ~n5543 & ~n5547;
  assign n5796 = ~n5794 & ~n5795;
  assign n5797 = ~n5793 ^ n5796;
  assign n5798 = n5587 & n5592;
  assign n5799 = n5581 & n5586;
  assign n5800 = ~n5798 & ~n5799;
  assign n5801 = ~n5797 ^ ~n5800;
  assign n5802 = n5551 & ~n5552;
  assign n5803 = ~n5549 & ~n5550;
  assign n5804 = ~n5802 & ~n5803;
  assign n5805 = n5579 & ~n5580;
  assign n5806 = ~n5577 & ~n5578;
  assign n5807 = ~n5805 & ~n5806;
  assign n5808 = ~n5804 ^ ~n5807;
  assign n5809 = n5541 & ~n5542;
  assign n5810 = ~n5539 & ~n5540;
  assign n5811 = ~n5809 & ~n5810;
  assign n5812 = ~n5808 ^ ~n5811;
  assign n5813 = n5584 & ~n5585;
  assign n5814 = ~n5582 & ~n5583;
  assign n5815 = ~n5813 & ~n5814;
  assign n5816 = n5590 & ~n5591;
  assign n5817 = ~n5588 & ~n5589;
  assign n5818 = ~n5816 & ~n5817;
  assign n5819 = ~n5815 ^ ~n5818;
  assign n5820 = pi01 & pi58;
  assign n5821 = ~n5820 ^ ~pi30;
  assign n5822 = ~n5819 ^ ~n5821;
  assign n5823 = ~n5812 ^ ~n5822;
  assign n5824 = n5523 & ~n5524;
  assign n5825 = ~n5521 & ~n5522;
  assign n5826 = ~n5824 & ~n5825;
  assign n5827 = n5534 & ~n5535;
  assign n5828 = ~n5532 & ~n5533;
  assign n5829 = ~n5827 & ~n5828;
  assign n5830 = ~n5826 ^ ~n5829;
  assign n5831 = n5545 & ~n5546;
  assign n5832 = ~n2744 & ~n5544;
  assign n5833 = ~n5831 & ~n5832;
  assign n5834 = ~n5830 ^ ~n5833;
  assign n5835 = ~n5823 ^ ~n5834;
  assign n5836 = ~n5801 ^ ~n5835;
  assign n5837 = ~n5790 ^ n5836;
  assign n5838 = ~n5787 ^ n5837;
  assign n5839 = ~n5680 & n5675;
  assign n5840 = ~n5839 & n5672;
  assign n5841 = n5680 & ~n5675;
  assign n5842 = ~n5840 & ~n5841;
  assign n5843 = ~n5838 ^ n5842;
  assign n5844 = n5555 & n5595;
  assign n5845 = ~n5844 & ~n5600;
  assign n5846 = ~n5555 & ~n5595;
  assign n5847 = ~n5845 & ~n5846;
  assign n5848 = n5576 & ~n5593;
  assign n5849 = n5558 & ~n5848;
  assign n5850 = ~n5576 & n5593;
  assign n5851 = ~n5849 & ~n5850;
  assign n5852 = n5637 & ~n5648;
  assign n5853 = n5633 & ~n5636;
  assign n5854 = ~n5852 & ~n5853;
  assign n5855 = ~n5568 & n5575;
  assign n5856 = n5571 & n5574;
  assign n5857 = ~n5855 & ~n5856;
  assign n5858 = n5644 & ~n5647;
  assign n5859 = ~n5640 & ~n5643;
  assign n5860 = ~n5858 & ~n5859;
  assign n5861 = ~n5857 ^ n5860;
  assign n5862 = n5629 & n5632;
  assign n5863 = n5625 & n5628;
  assign n5864 = ~n5862 & ~n5863;
  assign n5865 = ~n5861 ^ n5864;
  assign n5866 = ~n5854 ^ n5865;
  assign n5867 = ~n5851 ^ ~n5866;
  assign n5868 = n5622 & n5649;
  assign n5869 = ~n5605 & ~n5868;
  assign n5870 = ~n5622 & ~n5649;
  assign n5871 = ~n5869 & ~n5870;
  assign n5872 = ~n5867 ^ ~n5871;
  assign n5873 = ~n5847 ^ ~n5872;
  assign n5874 = ~n5843 ^ ~n5873;
  assign n5875 = n5601 & n5651;
  assign n5876 = ~n5517 & ~n5875;
  assign n5877 = ~n5601 & ~n5651;
  assign n5878 = ~n5876 & ~n5877;
  assign n5879 = ~n5874 ^ n5878;
  assign n5880 = ~n5701 ^ n5879;
  assign po060 = n5697 ^ ~n5880;
  assign n5882 = n5701 & ~n5879;
  assign n5883 = ~n5697 & ~n5882;
  assign n5884 = ~n5701 & n5879;
  assign n5885 = ~n5883 & ~n5884;
  assign n5886 = ~n5843 & ~n5873;
  assign n5887 = ~n5886 & ~n5878;
  assign n5888 = n5843 & n5873;
  assign n5889 = ~n5887 & ~n5888;
  assign n5890 = n5787 & ~n5837;
  assign n5891 = ~n5890 & ~n5842;
  assign n5892 = ~n5787 & n5837;
  assign n5893 = ~n5891 & ~n5892;
  assign n5894 = ~n5867 & ~n5871;
  assign n5895 = n5847 & ~n5894;
  assign n5896 = n5867 & n5871;
  assign n5897 = ~n5895 & ~n5896;
  assign n5898 = n5854 & ~n5865;
  assign n5899 = n5851 & ~n5898;
  assign n5900 = ~n5854 & n5865;
  assign n5901 = ~n5899 & ~n5900;
  assign n5902 = n5857 & ~n5860;
  assign n5903 = ~n5902 & ~n5864;
  assign n5904 = ~n5857 & n5860;
  assign n5905 = ~n5903 & ~n5904;
  assign n5906 = pi26 & pi34;
  assign n5907 = pi25 & pi35;
  assign n5908 = ~n5906 ^ ~n5907;
  assign n5909 = pi24 & pi36;
  assign n5910 = ~n5908 ^ n5909;
  assign n5911 = pi21 & pi39;
  assign n5912 = pi22 & pi38;
  assign n5913 = ~n5911 ^ ~n5912;
  assign n5914 = pi20 & pi40;
  assign n5915 = ~n5913 ^ n5914;
  assign n5916 = ~n5910 ^ ~n5915;
  assign n5917 = pi04 & pi56;
  assign n5918 = pi03 & pi57;
  assign n5919 = ~n5917 ^ ~n5918;
  assign n5920 = pi02 & pi58;
  assign n5921 = ~n5919 ^ n5920;
  assign n5922 = ~n5916 ^ ~n5921;
  assign n5923 = n5711 & ~n5712;
  assign n5924 = ~n5709 & ~n5710;
  assign n5925 = ~n5923 & ~n5924;
  assign n5926 = pi17 & pi43;
  assign n5927 = pi16 & pi44;
  assign n5928 = ~n5926 ^ ~n5927;
  assign n5929 = pi09 & pi51;
  assign n5930 = ~n5928 ^ n5929;
  assign n5931 = pi15 & pi45;
  assign n5932 = pi11 & pi49;
  assign n5933 = ~n5931 ^ ~n5932;
  assign n5934 = pi10 & pi50;
  assign n5935 = ~n5933 ^ n5934;
  assign n5936 = ~n5930 ^ ~n5935;
  assign n5937 = ~n5925 ^ n5936;
  assign n5938 = ~n5922 ^ ~n5937;
  assign n5939 = ~n5905 ^ n5938;
  assign n5940 = n5823 & n5834;
  assign n5941 = n5812 & n5822;
  assign n5942 = ~n5940 & ~n5941;
  assign n5943 = n5819 & n5821;
  assign n5944 = n5815 & n5818;
  assign n5945 = ~n5943 & ~n5944;
  assign n5946 = n1769 & pi58;
  assign n5947 = pi01 & pi59;
  assign n5948 = pi29 & pi31;
  assign n5949 = ~n5947 ^ ~n5948;
  assign n5950 = ~n5946 ^ ~n5949;
  assign n5951 = pi00 & pi60;
  assign n5952 = ~n5950 ^ n5951;
  assign n5953 = pi28 & pi32;
  assign n5954 = pi27 & pi33;
  assign n5955 = ~n5953 ^ ~n5954;
  assign n5956 = pi23 & pi37;
  assign n5957 = ~n5955 ^ n5956;
  assign n5958 = ~n5952 ^ ~n5957;
  assign n5959 = ~n5945 ^ n5958;
  assign n5960 = pi14 & pi46;
  assign n5961 = pi13 & pi47;
  assign n5962 = ~n5960 ^ ~n5961;
  assign n5963 = pi12 & pi48;
  assign n5964 = ~n5962 ^ n5963;
  assign n5965 = pi18 & pi42;
  assign n5966 = pi08 & pi52;
  assign n5967 = ~n5965 ^ ~n5966;
  assign n5968 = pi07 & pi53;
  assign n5969 = ~n5967 ^ n5968;
  assign n5970 = ~n5964 ^ ~n5969;
  assign n5971 = pi19 & pi41;
  assign n5972 = pi06 & pi54;
  assign n5973 = ~n5971 ^ ~n5972;
  assign n5974 = pi05 & pi55;
  assign n5975 = ~n5973 ^ n5974;
  assign n5976 = ~n5970 ^ ~n5975;
  assign n5977 = ~n5959 ^ n5976;
  assign n5978 = ~n5942 ^ n5977;
  assign n5979 = ~n5939 ^ ~n5978;
  assign n5980 = ~n5901 ^ ~n5979;
  assign n5981 = n5726 & ~n5741;
  assign n5982 = n5708 & n5725;
  assign n5983 = ~n5981 & ~n5982;
  assign n5984 = ~n5754 & n5765;
  assign n5985 = ~n5759 & ~n5764;
  assign n5986 = ~n5984 & ~n5985;
  assign n5987 = n5769 & ~n5770;
  assign n5988 = ~n5767 & ~n5768;
  assign n5989 = ~n5987 & ~n5988;
  assign n5990 = n5732 & ~n5733;
  assign n5991 = ~n5730 & ~n5731;
  assign n5992 = ~n5990 & ~n5991;
  assign n5993 = ~n5989 ^ ~n5992;
  assign n5994 = n5780 & ~n5781;
  assign n5995 = ~n5778 & ~n5779;
  assign n5996 = ~n5994 & ~n5995;
  assign n5997 = ~n5993 ^ n5996;
  assign n5998 = ~n5986 ^ ~n5997;
  assign n5999 = ~n5739 & ~pi02;
  assign n6000 = n5736 & ~n5999;
  assign n6001 = n5739 & pi02;
  assign n6002 = ~n6000 & ~n6001;
  assign n6003 = ~n6002 & pi57;
  assign n6004 = n5762 & ~n5763;
  assign n6005 = ~n5760 & ~n5761;
  assign n6006 = ~n6004 & ~n6005;
  assign n6007 = n5774 & ~n5775;
  assign n6008 = ~n5772 & ~n5773;
  assign n6009 = ~n6007 & ~n6008;
  assign n6010 = ~n6006 ^ ~n6009;
  assign n6011 = ~n6003 ^ n6010;
  assign n6012 = ~n5998 ^ n6011;
  assign n6013 = ~n5983 ^ ~n6012;
  assign n6014 = n5716 & ~n5717;
  assign n6015 = ~n5714 & ~n5715;
  assign n6016 = ~n6014 & ~n6015;
  assign n6017 = n5757 & ~n5758;
  assign n6018 = ~n5755 & ~n5756;
  assign n6019 = ~n6017 & ~n6018;
  assign n6020 = ~n6016 ^ ~n6019;
  assign n6021 = n5722 & ~n5723;
  assign n6022 = ~n5720 & ~n5721;
  assign n6023 = ~n6021 & ~n6022;
  assign n6024 = ~n6020 ^ ~n6023;
  assign n6025 = n5719 & n5724;
  assign n6026 = n5713 & n5718;
  assign n6027 = ~n6025 & ~n6026;
  assign n6028 = ~n6024 ^ ~n6027;
  assign n6029 = n5777 & n5782;
  assign n6030 = n5771 & n5776;
  assign n6031 = ~n6029 & ~n6030;
  assign n6032 = ~n6028 ^ ~n6031;
  assign n6033 = ~n6013 ^ n6032;
  assign n6034 = ~n5980 ^ ~n6033;
  assign n6035 = ~n5897 ^ n6034;
  assign n6036 = n5742 & n5785;
  assign n6037 = n5705 & ~n6036;
  assign n6038 = ~n5742 & ~n5785;
  assign n6039 = ~n6037 & ~n6038;
  assign n6040 = ~n5801 & ~n5835;
  assign n6041 = ~n5790 & ~n6040;
  assign n6042 = n5801 & n5835;
  assign n6043 = ~n6041 & ~n6042;
  assign n6044 = ~n5766 & n5783;
  assign n6045 = n5745 & ~n6044;
  assign n6046 = n5766 & ~n5783;
  assign n6047 = ~n6045 & ~n6046;
  assign n6048 = n5797 & n5800;
  assign n6049 = n5793 & ~n5796;
  assign n6050 = ~n6048 & ~n6049;
  assign n6051 = n5830 & n5833;
  assign n6052 = n5826 & n5829;
  assign n6053 = ~n6051 & ~n6052;
  assign n6054 = n5808 & n5811;
  assign n6055 = n5804 & n5807;
  assign n6056 = ~n6054 & ~n6055;
  assign n6057 = ~n6053 ^ ~n6056;
  assign n6058 = n5735 & n5740;
  assign n6059 = n5729 & ~n5734;
  assign n6060 = ~n6058 & ~n6059;
  assign n6061 = ~n6057 ^ n6060;
  assign n6062 = ~n6050 ^ n6061;
  assign n6063 = ~n6047 ^ ~n6062;
  assign n6064 = ~n6043 ^ ~n6063;
  assign n6065 = ~n6039 ^ ~n6064;
  assign n6066 = ~n6035 ^ n6065;
  assign n6067 = ~n5893 ^ ~n6066;
  assign n6068 = ~n5889 ^ ~n6067;
  assign po061 = n5885 ^ ~n6068;
  assign n6070 = ~n6035 & n6065;
  assign n6071 = n5893 & n6070;
  assign n6072 = ~n5889 & ~n6071;
  assign n6073 = ~n5893 & ~n6070;
  assign n6074 = n6035 & ~n6065;
  assign n6075 = ~n6073 & ~n6074;
  assign n6076 = ~n6072 & n6075;
  assign n6077 = n5885 & n6076;
  assign n6078 = ~n5893 & n6074;
  assign n6079 = ~n5889 & n6078;
  assign n6080 = ~n6077 & ~n6079;
  assign n6081 = n5889 & ~n6078;
  assign n6082 = ~n6081 & ~n6075;
  assign n6083 = ~n5885 & n6082;
  assign n6084 = n5889 & n6071;
  assign n6085 = ~n6083 & ~n6084;
  assign n6086 = n6080 & n6085;
  assign n6087 = ~n5980 & ~n6033;
  assign n6088 = n5897 & ~n6087;
  assign n6089 = n5980 & n6033;
  assign n6090 = ~n6088 & ~n6089;
  assign n6091 = n5939 & n5978;
  assign n6092 = n5901 & ~n6091;
  assign n6093 = ~n5939 & ~n5978;
  assign n6094 = ~n6092 & ~n6093;
  assign n6095 = n5998 & ~n6011;
  assign n6096 = ~n5986 & ~n5997;
  assign n6097 = ~n6095 & ~n6096;
  assign n6098 = n6028 & n6031;
  assign n6099 = n6024 & n6027;
  assign n6100 = ~n6098 & ~n6099;
  assign n6101 = pi28 & pi33;
  assign n6102 = pi27 & pi34;
  assign n6103 = ~n6101 ^ ~n6102;
  assign n6104 = pi26 & pi35;
  assign n6105 = ~n6103 ^ n6104;
  assign n6106 = pi19 & pi42;
  assign n6107 = pi08 & pi53;
  assign n6108 = ~n6106 ^ ~n6107;
  assign n6109 = pi07 & pi54;
  assign n6110 = ~n6108 ^ n6109;
  assign n6111 = ~n6105 ^ ~n6110;
  assign n6112 = pi18 & pi43;
  assign n6113 = pi17 & pi44;
  assign n6114 = ~n6112 ^ ~n6113;
  assign n6115 = pi09 & pi52;
  assign n6116 = ~n6114 ^ n6115;
  assign n6117 = ~n6111 ^ ~n6116;
  assign n6118 = ~n6100 ^ ~n6117;
  assign n6119 = ~n6097 ^ ~n6118;
  assign n6120 = ~n5922 & ~n5937;
  assign n6121 = n5905 & ~n6120;
  assign n6122 = n5922 & n5937;
  assign n6123 = ~n6121 & ~n6122;
  assign n6124 = n5993 & ~n5996;
  assign n6125 = ~n5989 & ~n5992;
  assign n6126 = ~n6124 & ~n6125;
  assign n6127 = n5962 & ~n5963;
  assign n6128 = ~n5960 & ~n5961;
  assign n6129 = ~n6127 & ~n6128;
  assign n6130 = pi29 & pi59;
  assign n6131 = n6130 & pi01;
  assign n6132 = ~n6131 & pi31;
  assign n6133 = pi01 & pi60;
  assign n6134 = ~n6132 ^ n6133;
  assign n6135 = ~n6129 ^ n6134;
  assign n6136 = ~n6126 ^ ~n6135;
  assign n6137 = ~n5925 & n5936;
  assign n6138 = n5930 & n5935;
  assign n6139 = ~n6137 & ~n6138;
  assign n6140 = ~n6136 ^ ~n6139;
  assign n6141 = n6020 & n6023;
  assign n6142 = n6016 & n6019;
  assign n6143 = ~n6141 & ~n6142;
  assign n6144 = pi23 & pi38;
  assign n6145 = pi04 & pi57;
  assign n6146 = ~n6144 ^ ~n6145;
  assign n6147 = pi03 & pi58;
  assign n6148 = ~n6146 ^ n6147;
  assign n6149 = ~n6143 ^ ~n6148;
  assign n6150 = ~n6003 & n6010;
  assign n6151 = ~n6006 & ~n6009;
  assign n6152 = ~n6150 & ~n6151;
  assign n6153 = ~n6149 ^ ~n6152;
  assign n6154 = ~n6140 ^ ~n6153;
  assign n6155 = ~n6123 ^ n6154;
  assign n6156 = ~n6119 ^ ~n6155;
  assign n6157 = ~n6094 ^ n6156;
  assign n6158 = ~n6090 ^ n6157;
  assign n6159 = n6043 & n6063;
  assign n6160 = ~n6039 & ~n6159;
  assign n6161 = ~n6043 & ~n6063;
  assign n6162 = ~n6160 & ~n6161;
  assign n6163 = n6013 & ~n6032;
  assign n6164 = ~n5983 & ~n6012;
  assign n6165 = ~n6163 & ~n6164;
  assign n6166 = n6050 & ~n6061;
  assign n6167 = ~n6047 & ~n6166;
  assign n6168 = ~n6050 & n6061;
  assign n6169 = ~n6167 & ~n6168;
  assign n6170 = n6057 & ~n6060;
  assign n6171 = ~n6053 & ~n6056;
  assign n6172 = ~n6170 & ~n6171;
  assign n6173 = pi14 & pi47;
  assign n6174 = pi12 & pi49;
  assign n6175 = ~n6173 ^ ~n6174;
  assign n6176 = pi11 & pi50;
  assign n6177 = ~n6175 ^ n6176;
  assign n6178 = pi16 & pi45;
  assign n6179 = pi15 & pi46;
  assign n6180 = ~n6178 ^ ~n6179;
  assign n6181 = pi10 & pi51;
  assign n6182 = ~n6180 ^ n6181;
  assign n6183 = ~n6177 ^ ~n6182;
  assign n6184 = pi30 & pi31;
  assign n6185 = pi29 & pi32;
  assign n6186 = ~n6184 ^ ~n6185;
  assign n6187 = pi13 & pi48;
  assign n6188 = ~n6186 ^ n6187;
  assign n6189 = ~n6183 ^ n6188;
  assign n6190 = pi05 & pi56;
  assign n6191 = pi02 & pi59;
  assign n6192 = ~n6190 ^ ~n6191;
  assign n6193 = pi00 & pi61;
  assign n6194 = ~n6192 ^ n6193;
  assign n6195 = pi25 & pi36;
  assign n6196 = pi24 & pi37;
  assign n6197 = ~n6195 ^ ~n6196;
  assign n6198 = pi22 & pi39;
  assign n6199 = ~n6197 ^ n6198;
  assign n6200 = ~n6194 ^ ~n6199;
  assign n6201 = ~n3040 ^ ~n3208;
  assign n6202 = pi06 & pi55;
  assign n6203 = ~n6201 ^ n6202;
  assign n6204 = ~n6200 ^ ~n6203;
  assign n6205 = ~n6189 ^ n6204;
  assign n6206 = ~n6172 ^ ~n6205;
  assign n6207 = ~n6169 ^ ~n6206;
  assign n6208 = ~n6165 ^ ~n6207;
  assign n6209 = ~n5959 & n5976;
  assign n6210 = ~n5942 & ~n6209;
  assign n6211 = n5959 & ~n5976;
  assign n6212 = ~n6210 & ~n6211;
  assign n6213 = n5913 & ~n5914;
  assign n6214 = ~n5911 & ~n5912;
  assign n6215 = ~n6213 & ~n6214;
  assign n6216 = n5955 & ~n5956;
  assign n6217 = ~n5953 & ~n5954;
  assign n6218 = ~n6216 & ~n6217;
  assign n6219 = ~n6215 ^ ~n6218;
  assign n6220 = n5908 & ~n5909;
  assign n6221 = ~n5906 & ~n5907;
  assign n6222 = ~n6220 & ~n6221;
  assign n6223 = ~n6219 ^ ~n6222;
  assign n6224 = n5973 & ~n5974;
  assign n6225 = ~n5971 & ~n5972;
  assign n6226 = ~n6224 & ~n6225;
  assign n6227 = n5919 & ~n5920;
  assign n6228 = ~n5917 & ~n5918;
  assign n6229 = ~n6227 & ~n6228;
  assign n6230 = ~n6226 ^ ~n6229;
  assign n6231 = n5933 & ~n5934;
  assign n6232 = ~n5931 & ~n5932;
  assign n6233 = ~n6231 & ~n6232;
  assign n6234 = ~n6230 ^ ~n6233;
  assign n6235 = ~n6223 ^ ~n6234;
  assign n6236 = n5916 & n5921;
  assign n6237 = n5910 & n5915;
  assign n6238 = ~n6236 & ~n6237;
  assign n6239 = ~n6235 ^ ~n6238;
  assign n6240 = ~n6212 ^ n6239;
  assign n6241 = ~n5959 & ~n5957;
  assign n6242 = ~n5945 & ~n5952;
  assign n6243 = ~n6241 & ~n6242;
  assign n6244 = n5970 & n5975;
  assign n6245 = n5964 & n5969;
  assign n6246 = ~n6244 & ~n6245;
  assign n6247 = ~n6243 ^ n6246;
  assign n6248 = n5952 & n5949;
  assign n6249 = n5946 & n5951;
  assign n6250 = ~n6248 & ~n6249;
  assign n6251 = n5928 & ~n5929;
  assign n6252 = ~n5926 & ~n5927;
  assign n6253 = ~n6251 & ~n6252;
  assign n6254 = n5967 & ~n5968;
  assign n6255 = ~n5965 & ~n5966;
  assign n6256 = ~n6254 & ~n6255;
  assign n6257 = ~n6253 ^ ~n6256;
  assign n6258 = ~n6250 ^ n6257;
  assign n6259 = ~n6247 ^ n6258;
  assign n6260 = ~n6240 ^ ~n6259;
  assign n6261 = ~n6208 ^ n6260;
  assign n6262 = ~n6162 ^ n6261;
  assign n6263 = ~n6158 ^ n6262;
  assign po062 = ~n6086 ^ n6263;
  assign n6265 = ~n6079 & n6263;
  assign n6266 = ~n6076 & ~n6265;
  assign n6267 = n5885 & ~n6266;
  assign n6268 = ~n6082 & n6263;
  assign n6269 = ~n6268 & ~n6084;
  assign n6270 = ~n6267 & n6269;
  assign n6271 = n6208 & ~n6260;
  assign n6272 = n6162 & ~n6271;
  assign n6273 = ~n6208 & n6260;
  assign n6274 = ~n6272 & ~n6273;
  assign n6275 = n6119 & n6155;
  assign n6276 = n6094 & ~n6275;
  assign n6277 = ~n6119 & ~n6155;
  assign n6278 = ~n6276 & ~n6277;
  assign n6279 = ~n6140 & ~n6153;
  assign n6280 = n6123 & ~n6279;
  assign n6281 = n6140 & n6153;
  assign n6282 = ~n6280 & ~n6281;
  assign n6283 = ~n1844 & ~pi02;
  assign n6284 = ~n6283 & pi60;
  assign n6285 = n1844 & pi02;
  assign n6286 = n6284 & ~n6285;
  assign n6287 = pi00 & pi62;
  assign n6288 = ~n6286 ^ ~n6287;
  assign n6289 = pi17 & pi45;
  assign n6290 = pi10 & pi52;
  assign n6291 = ~n6289 ^ ~n6290;
  assign n6292 = pi09 & pi53;
  assign n6293 = ~n6291 ^ n6292;
  assign n6294 = ~n6288 ^ n6293;
  assign n6295 = pi26 & pi36;
  assign n6296 = pi25 & pi37;
  assign n6297 = ~n6295 ^ ~n6296;
  assign n6298 = pi21 & pi41;
  assign n6299 = ~n6297 ^ n6298;
  assign n6300 = ~n6294 ^ ~n6299;
  assign n6301 = pi19 & pi43;
  assign n6302 = pi18 & pi44;
  assign n6303 = ~n6301 ^ ~n6302;
  assign n6304 = pi08 & pi54;
  assign n6305 = ~n6303 ^ n6304;
  assign n6306 = pi24 & pi38;
  assign n6307 = pi23 & pi39;
  assign n6308 = ~n6306 ^ ~n6307;
  assign n6309 = pi22 & pi40;
  assign n6310 = ~n6308 ^ n6309;
  assign n6311 = ~n6305 ^ ~n6310;
  assign n6312 = pi29 & pi33;
  assign n6313 = pi28 & pi34;
  assign n6314 = ~n6312 ^ ~n6313;
  assign n6315 = pi27 & pi35;
  assign n6316 = ~n6314 ^ n6315;
  assign n6317 = ~n6311 ^ ~n6316;
  assign n6318 = ~n6300 ^ ~n6317;
  assign n6319 = pi14 & pi48;
  assign n6320 = pi13 & pi49;
  assign n6321 = ~n6319 ^ ~n6320;
  assign n6322 = pi12 & pi50;
  assign n6323 = ~n6321 ^ n6322;
  assign n6324 = pi16 & pi46;
  assign n6325 = pi15 & pi47;
  assign n6326 = ~n6324 ^ ~n6325;
  assign n6327 = pi11 & pi51;
  assign n6328 = ~n6326 ^ n6327;
  assign n6329 = ~n6323 ^ ~n6328;
  assign n6330 = pi20 & pi42;
  assign n6331 = pi07 & pi55;
  assign n6332 = ~n6330 ^ ~n6331;
  assign n6333 = pi06 & pi56;
  assign n6334 = ~n6332 ^ n6333;
  assign n6335 = ~n6329 ^ ~n6334;
  assign n6336 = ~n6318 ^ n6335;
  assign n6337 = ~n6282 ^ n6336;
  assign n6338 = ~n6212 & n6239;
  assign n6339 = ~n6338 & n6259;
  assign n6340 = n6212 & ~n6239;
  assign n6341 = ~n6339 & ~n6340;
  assign n6342 = ~n6337 ^ ~n6341;
  assign n6343 = n6149 & n6152;
  assign n6344 = ~n6143 & ~n6148;
  assign n6345 = ~n6343 & ~n6344;
  assign n6346 = n6114 & ~n6115;
  assign n6347 = ~n6112 & ~n6113;
  assign n6348 = ~n6346 & ~n6347;
  assign n6349 = pi05 & pi57;
  assign n6350 = pi04 & pi58;
  assign n6351 = ~n6349 ^ ~n6350;
  assign n6352 = pi03 & pi59;
  assign n6353 = ~n6351 ^ n6352;
  assign n6354 = ~n6348 ^ n6353;
  assign n6355 = n6180 & ~n6181;
  assign n6356 = ~n6178 & ~n6179;
  assign n6357 = ~n6355 & ~n6356;
  assign n6358 = ~n6354 ^ n6357;
  assign n6359 = ~n6345 ^ ~n6358;
  assign n6360 = n6111 & n6116;
  assign n6361 = n6105 & n6110;
  assign n6362 = ~n6360 & ~n6361;
  assign n6363 = ~n6359 ^ ~n6362;
  assign n6364 = n6129 & pi60;
  assign n6365 = pi31 & pi59;
  assign n6366 = n6365 & pi29;
  assign n6367 = ~n6364 & ~n6366;
  assign n6368 = pi31 & pi60;
  assign n6369 = ~n6368 & pi01;
  assign n6370 = ~n6367 & n6369;
  assign n6371 = ~n6130 & n6133;
  assign n6372 = ~n6371 & pi31;
  assign n6373 = n6129 & n6372;
  assign n6374 = ~n6370 & ~n6373;
  assign n6375 = ~n6250 & n6257;
  assign n6376 = n6253 & n6256;
  assign n6377 = ~n6375 & ~n6376;
  assign n6378 = ~n6374 ^ ~n6377;
  assign n6379 = n6219 & n6222;
  assign n6380 = n6215 & n6218;
  assign n6381 = ~n6379 & ~n6380;
  assign n6382 = ~n6378 ^ n6381;
  assign n6383 = ~n6363 ^ ~n6382;
  assign n6384 = n6189 & ~n6204;
  assign n6385 = n6172 & ~n6384;
  assign n6386 = ~n6189 & n6204;
  assign n6387 = ~n6385 & ~n6386;
  assign n6388 = ~n6383 ^ ~n6387;
  assign n6389 = ~n6342 ^ ~n6388;
  assign n6390 = ~n6278 ^ n6389;
  assign n6391 = n6169 & n6206;
  assign n6392 = n6165 & ~n6391;
  assign n6393 = ~n6169 & ~n6206;
  assign n6394 = ~n6392 & ~n6393;
  assign n6395 = n6100 & n6117;
  assign n6396 = ~n6097 & ~n6395;
  assign n6397 = ~n6100 & ~n6117;
  assign n6398 = ~n6396 & ~n6397;
  assign n6399 = n6230 & n6233;
  assign n6400 = n6226 & n6229;
  assign n6401 = ~n6399 & ~n6400;
  assign n6402 = n6200 & n6203;
  assign n6403 = n6194 & n6199;
  assign n6404 = ~n6402 & ~n6403;
  assign n6405 = ~n6401 ^ n6404;
  assign n6406 = n6183 & ~n6188;
  assign n6407 = ~n6177 & ~n6182;
  assign n6408 = ~n6406 & ~n6407;
  assign n6409 = ~n6405 ^ n6408;
  assign n6410 = n6186 & ~n6187;
  assign n6411 = ~n6184 & ~n6185;
  assign n6412 = ~n6410 & ~n6411;
  assign n6413 = n6175 & ~n6176;
  assign n6414 = ~n6173 & ~n6174;
  assign n6415 = ~n6413 & ~n6414;
  assign n6416 = ~n6412 ^ ~n6415;
  assign n6417 = pi01 & pi61;
  assign n6418 = pi30 & pi32;
  assign n6419 = ~n6417 ^ ~n6418;
  assign n6420 = ~n6416 ^ ~n6419;
  assign n6421 = n6192 & ~n6193;
  assign n6422 = ~n6190 & ~n6191;
  assign n6423 = ~n6421 & ~n6422;
  assign n6424 = n6108 & ~n6109;
  assign n6425 = ~n6106 & ~n6107;
  assign n6426 = ~n6424 & ~n6425;
  assign n6427 = ~n6423 ^ ~n6426;
  assign n6428 = n6201 & ~n6202;
  assign n6429 = ~n3040 & ~n3208;
  assign n6430 = ~n6428 & ~n6429;
  assign n6431 = ~n6427 ^ n6430;
  assign n6432 = ~n6420 ^ n6431;
  assign n6433 = n6103 & ~n6104;
  assign n6434 = ~n6101 & ~n6102;
  assign n6435 = ~n6433 & ~n6434;
  assign n6436 = n6197 & ~n6198;
  assign n6437 = ~n6195 & ~n6196;
  assign n6438 = ~n6436 & ~n6437;
  assign n6439 = ~n6435 ^ ~n6438;
  assign n6440 = n6146 & ~n6147;
  assign n6441 = ~n6144 & ~n6145;
  assign n6442 = ~n6440 & ~n6441;
  assign n6443 = ~n6439 ^ ~n6442;
  assign n6444 = ~n6432 ^ n6443;
  assign n6445 = ~n6409 ^ n6444;
  assign n6446 = ~n6398 ^ ~n6445;
  assign n6447 = n6247 & ~n6258;
  assign n6448 = n6243 & ~n6246;
  assign n6449 = ~n6447 & ~n6448;
  assign n6450 = n6136 & n6139;
  assign n6451 = n6126 & n6135;
  assign n6452 = ~n6450 & ~n6451;
  assign n6453 = n6235 & n6238;
  assign n6454 = n6223 & n6234;
  assign n6455 = ~n6453 & ~n6454;
  assign n6456 = ~n6452 ^ ~n6455;
  assign n6457 = ~n6449 ^ ~n6456;
  assign n6458 = ~n6446 ^ n6457;
  assign n6459 = ~n6394 ^ n6458;
  assign n6460 = ~n6390 ^ ~n6459;
  assign n6461 = ~n6274 ^ n6460;
  assign n6462 = ~n6090 & n6157;
  assign n6463 = ~n6462 & n6262;
  assign n6464 = n6090 & ~n6157;
  assign n6465 = ~n6463 & ~n6464;
  assign n6466 = ~n6461 ^ ~n6465;
  assign po063 = n6270 ^ n6466;
  assign n6468 = n6461 & n6465;
  assign n6469 = n6270 & ~n6468;
  assign n6470 = ~n6461 & ~n6465;
  assign n6471 = ~n6469 & ~n6470;
  assign n6472 = ~n6390 & ~n6459;
  assign n6473 = n6274 & ~n6472;
  assign n6474 = n6390 & n6459;
  assign n6475 = ~n6473 & ~n6474;
  assign n6476 = n6342 & n6388;
  assign n6477 = n6278 & ~n6476;
  assign n6478 = ~n6342 & ~n6388;
  assign n6479 = ~n6477 & ~n6478;
  assign n6480 = n6341 & n6336;
  assign n6481 = ~n6480 & n6282;
  assign n6482 = ~n6341 & ~n6336;
  assign n6483 = ~n6481 & ~n6482;
  assign n6484 = n6359 & n6362;
  assign n6485 = ~n6345 & ~n6358;
  assign n6486 = ~n6484 & ~n6485;
  assign n6487 = n6405 & ~n6408;
  assign n6488 = ~n6401 & n6404;
  assign n6489 = ~n6487 & ~n6488;
  assign n6490 = n6432 & ~n6443;
  assign n6491 = ~n6420 & n6431;
  assign n6492 = ~n6490 & ~n6491;
  assign n6493 = ~n6489 ^ n6492;
  assign n6494 = ~n6486 ^ n6493;
  assign n6495 = n6318 & ~n6335;
  assign n6496 = ~n6300 & ~n6317;
  assign n6497 = ~n6495 & ~n6496;
  assign n6498 = n6439 & n6442;
  assign n6499 = n6435 & n6438;
  assign n6500 = ~n6498 & ~n6499;
  assign n6501 = n6354 & ~n6357;
  assign n6502 = ~n6348 & n6353;
  assign n6503 = ~n6501 & ~n6502;
  assign n6504 = ~n6500 ^ n6503;
  assign n6505 = n6416 & n6419;
  assign n6506 = n6412 & n6415;
  assign n6507 = ~n6505 & ~n6506;
  assign n6508 = ~n6504 ^ n6507;
  assign n6509 = n6427 & ~n6430;
  assign n6510 = ~n6423 & ~n6426;
  assign n6511 = ~n6509 & ~n6510;
  assign n6512 = ~n6285 & ~n6287;
  assign n6513 = n6284 & ~n6512;
  assign n6514 = n6351 & ~n6352;
  assign n6515 = ~n6349 & ~n6350;
  assign n6516 = ~n6514 & ~n6515;
  assign n6517 = ~n6513 ^ ~n6516;
  assign n6518 = n6297 & ~n6298;
  assign n6519 = ~n6295 & ~n6296;
  assign n6520 = ~n6518 & ~n6519;
  assign n6521 = ~n6517 ^ ~n6520;
  assign n6522 = n6321 & ~n6322;
  assign n6523 = ~n6319 & ~n6320;
  assign n6524 = ~n6522 & ~n6523;
  assign n6525 = n6308 & ~n6309;
  assign n6526 = ~n6306 & ~n6307;
  assign n6527 = ~n6525 & ~n6526;
  assign n6528 = ~n6524 ^ ~n6527;
  assign n6529 = n6332 & ~n6333;
  assign n6530 = ~n6330 & ~n6331;
  assign n6531 = ~n6529 & ~n6530;
  assign n6532 = ~n6528 ^ n6531;
  assign n6533 = ~n6521 ^ n6532;
  assign n6534 = ~n6511 ^ n6533;
  assign n6535 = ~n6508 ^ n6534;
  assign n6536 = ~n6497 ^ ~n6535;
  assign n6537 = ~n6494 ^ n6536;
  assign n6538 = ~n6483 ^ ~n6537;
  assign n6539 = ~n6479 ^ ~n6538;
  assign n6540 = n6446 & ~n6457;
  assign n6541 = ~n6394 & ~n6540;
  assign n6542 = ~n6446 & n6457;
  assign n6543 = ~n6541 & ~n6542;
  assign n6544 = ~n6363 & ~n6382;
  assign n6545 = ~n6544 & n6387;
  assign n6546 = n6363 & n6382;
  assign n6547 = ~n6545 & ~n6546;
  assign n6548 = pi31 & pi32;
  assign n6549 = pi30 & pi33;
  assign n6550 = ~n6548 ^ ~n6549;
  assign n6551 = pi14 & pi49;
  assign n6552 = ~n6550 ^ n6551;
  assign n6553 = pi23 & pi40;
  assign n6554 = pi20 & pi43;
  assign n6555 = ~n6553 ^ ~n6554;
  assign n6556 = pi06 & pi57;
  assign n6557 = ~n6555 ^ n6556;
  assign n6558 = ~n6552 ^ ~n6557;
  assign n6559 = pi19 & pi44;
  assign n6560 = pi08 & pi55;
  assign n6561 = ~n6559 ^ ~n6560;
  assign n6562 = pi07 & pi56;
  assign n6563 = ~n6561 ^ n6562;
  assign n6564 = ~n6558 ^ n6563;
  assign n6565 = pi15 & pi48;
  assign n6566 = pi13 & pi50;
  assign n6567 = ~n6565 ^ ~n6566;
  assign n6568 = pi12 & pi51;
  assign n6569 = ~n6567 ^ n6568;
  assign n6570 = pi18 & pi45;
  assign n6571 = pi17 & pi46;
  assign n6572 = ~n6570 ^ ~n6571;
  assign n6573 = pi09 & pi54;
  assign n6574 = ~n6572 ^ n6573;
  assign n6575 = ~n6569 ^ ~n6574;
  assign n6576 = pi16 & pi47;
  assign n6577 = pi11 & pi52;
  assign n6578 = ~n6576 ^ ~n6577;
  assign n6579 = pi10 & pi53;
  assign n6580 = ~n6578 ^ n6579;
  assign n6581 = ~n6575 ^ ~n6580;
  assign n6582 = ~n6564 ^ n6581;
  assign n6583 = n6326 & ~n6327;
  assign n6584 = ~n6324 & ~n6325;
  assign n6585 = ~n6583 & ~n6584;
  assign n6586 = pi04 & pi59;
  assign n6587 = pi03 & pi60;
  assign n6588 = ~n6586 ^ ~n6587;
  assign n6589 = pi02 & pi61;
  assign n6590 = ~n6588 ^ n6589;
  assign n6591 = pi22 & pi41;
  assign n6592 = pi21 & pi42;
  assign n6593 = ~n6591 ^ ~n6592;
  assign n6594 = pi05 & pi58;
  assign n6595 = ~n6593 ^ n6594;
  assign n6596 = ~n6590 ^ ~n6595;
  assign n6597 = ~n6585 ^ ~n6596;
  assign n6598 = ~n6582 ^ ~n6597;
  assign n6599 = ~n6547 ^ n6598;
  assign n6600 = ~n6409 & n6444;
  assign n6601 = ~n6398 & ~n6600;
  assign n6602 = n6409 & ~n6444;
  assign n6603 = ~n6601 & ~n6602;
  assign n6604 = ~n6599 ^ ~n6603;
  assign n6605 = ~n6452 & ~n6455;
  assign n6606 = ~n6449 & ~n6605;
  assign n6607 = n6452 & n6455;
  assign n6608 = ~n6606 & ~n6607;
  assign n6609 = n6378 & ~n6381;
  assign n6610 = ~n6374 & ~n6377;
  assign n6611 = ~n6609 & ~n6610;
  assign n6612 = n6294 & n6299;
  assign n6613 = ~n6288 & n6293;
  assign n6614 = ~n6612 & ~n6613;
  assign n6615 = pi29 & pi34;
  assign n6616 = pi28 & pi35;
  assign n6617 = ~n6615 ^ ~n6616;
  assign n6618 = pi27 & pi36;
  assign n6619 = ~n6617 ^ n6618;
  assign n6620 = pi26 & pi37;
  assign n6621 = pi25 & pi38;
  assign n6622 = ~n6620 ^ ~n6621;
  assign n6623 = pi24 & pi39;
  assign n6624 = ~n6622 ^ n6623;
  assign n6625 = ~n6619 ^ ~n6624;
  assign n6626 = pi30 & pi61;
  assign n6627 = n6626 & pi01;
  assign n6628 = ~n6627 & pi32;
  assign n6629 = pi00 & pi63;
  assign n6630 = pi01 & pi62;
  assign n6631 = ~n6629 ^ n6630;
  assign n6632 = ~n6628 ^ ~n6631;
  assign n6633 = ~n6625 ^ ~n6632;
  assign n6634 = ~n6614 ^ n6633;
  assign n6635 = ~n6611 ^ ~n6634;
  assign n6636 = n6303 & ~n6304;
  assign n6637 = ~n6301 & ~n6302;
  assign n6638 = ~n6636 & ~n6637;
  assign n6639 = n6291 & ~n6292;
  assign n6640 = ~n6289 & ~n6290;
  assign n6641 = ~n6639 & ~n6640;
  assign n6642 = ~n6638 ^ ~n6641;
  assign n6643 = n6314 & ~n6315;
  assign n6644 = ~n6312 & ~n6313;
  assign n6645 = ~n6643 & ~n6644;
  assign n6646 = ~n6642 ^ ~n6645;
  assign n6647 = n6329 & n6334;
  assign n6648 = n6323 & n6328;
  assign n6649 = ~n6647 & ~n6648;
  assign n6650 = ~n6646 ^ ~n6649;
  assign n6651 = n6311 & n6316;
  assign n6652 = n6305 & n6310;
  assign n6653 = ~n6651 & ~n6652;
  assign n6654 = ~n6650 ^ ~n6653;
  assign n6655 = ~n6635 ^ n6654;
  assign n6656 = ~n6608 ^ n6655;
  assign n6657 = ~n6604 ^ ~n6656;
  assign n6658 = ~n6543 ^ ~n6657;
  assign n6659 = ~n6539 ^ n6658;
  assign n6660 = ~n6475 ^ ~n6659;
  assign po064 = n6471 ^ n6660;
  assign n6662 = n6475 & ~n6479;
  assign n6663 = n6658 & ~n6538;
  assign n6664 = ~n6662 & ~n6663;
  assign n6665 = ~n6475 & n6479;
  assign n6666 = ~n6658 & n6538;
  assign n6667 = ~n6665 & ~n6666;
  assign n6668 = n6664 & ~n6667;
  assign n6669 = ~n6471 & n6668;
  assign n6670 = n6665 & n6666;
  assign n6671 = n6662 & n6663;
  assign n6672 = ~n6670 & ~n6671;
  assign n6673 = ~n6669 & n6672;
  assign n6674 = ~n6664 & n6667;
  assign n6675 = n6471 & n6674;
  assign n6676 = n6673 & ~n6675;
  assign n6677 = ~n6604 & ~n6656;
  assign n6678 = n6543 & ~n6677;
  assign n6679 = n6604 & n6656;
  assign n6680 = ~n6678 & ~n6679;
  assign n6681 = ~n6494 & n6536;
  assign n6682 = n6483 & ~n6681;
  assign n6683 = n6494 & ~n6536;
  assign n6684 = ~n6682 & ~n6683;
  assign n6685 = ~n6489 & n6492;
  assign n6686 = n6486 & ~n6685;
  assign n6687 = n6489 & ~n6492;
  assign n6688 = ~n6686 & ~n6687;
  assign n6689 = n6504 & ~n6507;
  assign n6690 = ~n6500 & n6503;
  assign n6691 = ~n6689 & ~n6690;
  assign n6692 = n6550 & ~n6551;
  assign n6693 = ~n6548 & ~n6549;
  assign n6694 = ~n6692 & ~n6693;
  assign n6695 = pi32 & pi62;
  assign n6696 = ~n6695 & ~pi63;
  assign n6697 = ~n6696 & pi01;
  assign n6698 = pi32 & pi63;
  assign n6699 = n6698 & pi62;
  assign n6700 = n6697 & ~n6699;
  assign n6701 = ~n6694 ^ ~n6700;
  assign n6702 = pi13 & pi51;
  assign n6703 = pi12 & pi52;
  assign n6704 = ~n6702 ^ ~n6703;
  assign n6705 = pi11 & pi53;
  assign n6706 = ~n6704 ^ n6705;
  assign n6707 = pi15 & pi49;
  assign n6708 = pi10 & pi54;
  assign n6709 = ~n6707 ^ ~n6708;
  assign n6710 = pi09 & pi55;
  assign n6711 = ~n6709 ^ n6710;
  assign n6712 = ~n6706 ^ ~n6711;
  assign n6713 = ~n6701 ^ ~n6712;
  assign n6714 = ~n6691 ^ n6713;
  assign n6715 = n6585 & n6596;
  assign n6716 = ~n6590 & ~n6595;
  assign n6717 = ~n6715 & ~n6716;
  assign n6718 = ~n6714 ^ n6717;
  assign n6719 = n6578 & ~n6579;
  assign n6720 = ~n6576 & ~n6577;
  assign n6721 = ~n6719 & ~n6720;
  assign n6722 = n6567 & ~n6568;
  assign n6723 = ~n6565 & ~n6566;
  assign n6724 = ~n6722 & ~n6723;
  assign n6725 = ~n6721 ^ ~n6724;
  assign n6726 = n6622 & ~n6623;
  assign n6727 = ~n6620 & ~n6621;
  assign n6728 = ~n6726 & ~n6727;
  assign n6729 = ~n6725 ^ ~n6728;
  assign n6730 = n6558 & ~n6563;
  assign n6731 = ~n6552 & ~n6557;
  assign n6732 = ~n6730 & ~n6731;
  assign n6733 = ~n6729 ^ n6732;
  assign n6734 = n6575 & n6580;
  assign n6735 = n6569 & n6574;
  assign n6736 = ~n6734 & ~n6735;
  assign n6737 = ~n6733 ^ n6736;
  assign n6738 = ~n6718 ^ n6737;
  assign n6739 = ~n6688 ^ ~n6738;
  assign n6740 = n6497 & n6535;
  assign n6741 = ~n6508 & n6534;
  assign n6742 = ~n6740 & ~n6741;
  assign n6743 = ~n6511 & n6533;
  assign n6744 = ~n6521 & n6532;
  assign n6745 = ~n6743 & ~n6744;
  assign n6746 = n6528 & ~n6531;
  assign n6747 = ~n6524 & ~n6527;
  assign n6748 = ~n6746 & ~n6747;
  assign n6749 = n6642 & n6645;
  assign n6750 = n6638 & n6641;
  assign n6751 = ~n6749 & ~n6750;
  assign n6752 = ~n6748 ^ n6751;
  assign n6753 = n6517 & n6520;
  assign n6754 = n6513 & n6516;
  assign n6755 = ~n6753 & ~n6754;
  assign n6756 = ~n6752 ^ n6755;
  assign n6757 = ~n6745 ^ ~n6756;
  assign n6758 = n6650 & n6653;
  assign n6759 = n6646 & n6649;
  assign n6760 = ~n6758 & ~n6759;
  assign n6761 = ~n6757 ^ ~n6760;
  assign n6762 = pi32 & pi61;
  assign n6763 = n1769 & n6762;
  assign n6764 = ~n6763 & ~n6630;
  assign n6765 = n6629 & ~pi32;
  assign n6766 = ~n6765 & pi62;
  assign n6767 = ~n6764 & ~n6766;
  assign n6768 = ~n6626 & n6630;
  assign n6769 = n6698 & pi00;
  assign n6770 = ~n6768 & n6769;
  assign n6771 = ~n6767 & ~n6770;
  assign n6772 = pi19 & pi45;
  assign n6773 = pi18 & pi46;
  assign n6774 = ~n6772 ^ ~n6773;
  assign n6775 = pi05 & pi59;
  assign n6776 = ~n6774 ^ n6775;
  assign n6777 = pi04 & pi60;
  assign n6778 = pi03 & pi61;
  assign n6779 = ~n6777 ^ ~n6778;
  assign n6780 = pi02 & pi62;
  assign n6781 = ~n6779 ^ n6780;
  assign n6782 = ~n6776 ^ ~n6781;
  assign n6783 = ~n6771 ^ n6782;
  assign n6784 = pi17 & pi47;
  assign n6785 = pi07 & pi57;
  assign n6786 = ~n6784 ^ ~n6785;
  assign n6787 = pi06 & pi58;
  assign n6788 = ~n6786 ^ n6787;
  assign n6789 = pi25 & pi39;
  assign n6790 = pi24 & pi40;
  assign n6791 = ~n6789 ^ ~n6790;
  assign n6792 = pi23 & pi41;
  assign n6793 = ~n6791 ^ n6792;
  assign n6794 = ~n6788 ^ ~n6793;
  assign n6795 = ~n3246 ^ ~n3500;
  assign n6796 = pi20 & pi44;
  assign n6797 = ~n6795 ^ n6796;
  assign n6798 = ~n6794 ^ ~n6797;
  assign n6799 = pi29 & pi35;
  assign n6800 = pi28 & pi36;
  assign n6801 = ~n6799 ^ ~n6800;
  assign n6802 = pi27 & pi37;
  assign n6803 = ~n6801 ^ n6802;
  assign n6804 = pi26 & pi38;
  assign n6805 = pi16 & pi48;
  assign n6806 = ~n6804 ^ ~n6805;
  assign n6807 = pi08 & pi56;
  assign n6808 = ~n6806 ^ n6807;
  assign n6809 = ~n6803 ^ ~n6808;
  assign n6810 = pi31 & pi33;
  assign n6811 = pi30 & pi34;
  assign n6812 = ~n6810 ^ ~n6811;
  assign n6813 = pi14 & pi50;
  assign n6814 = ~n6812 ^ n6813;
  assign n6815 = ~n6809 ^ ~n6814;
  assign n6816 = ~n6798 ^ ~n6815;
  assign n6817 = ~n6783 ^ ~n6816;
  assign n6818 = ~n6761 ^ n6817;
  assign n6819 = ~n6742 ^ ~n6818;
  assign n6820 = ~n6739 ^ ~n6819;
  assign n6821 = ~n6684 ^ ~n6820;
  assign n6822 = ~n6635 & n6654;
  assign n6823 = ~n6608 & ~n6822;
  assign n6824 = n6635 & ~n6654;
  assign n6825 = ~n6823 & ~n6824;
  assign n6826 = n6614 & ~n6633;
  assign n6827 = n6611 & ~n6826;
  assign n6828 = ~n6614 & n6633;
  assign n6829 = ~n6827 & ~n6828;
  assign n6830 = n6617 & ~n6618;
  assign n6831 = ~n6615 & ~n6616;
  assign n6832 = ~n6830 & ~n6831;
  assign n6833 = n6572 & ~n6573;
  assign n6834 = ~n6570 & ~n6571;
  assign n6835 = ~n6833 & ~n6834;
  assign n6836 = ~n6832 ^ ~n6835;
  assign n6837 = n6555 & ~n6556;
  assign n6838 = ~n6553 & ~n6554;
  assign n6839 = ~n6837 & ~n6838;
  assign n6840 = ~n6836 ^ ~n6839;
  assign n6841 = n6588 & ~n6589;
  assign n6842 = ~n6586 & ~n6587;
  assign n6843 = ~n6841 & ~n6842;
  assign n6844 = n6561 & ~n6562;
  assign n6845 = ~n6559 & ~n6560;
  assign n6846 = ~n6844 & ~n6845;
  assign n6847 = ~n6843 ^ ~n6846;
  assign n6848 = n6593 & ~n6594;
  assign n6849 = ~n6591 & ~n6592;
  assign n6850 = ~n6848 & ~n6849;
  assign n6851 = ~n6847 ^ n6850;
  assign n6852 = ~n6840 ^ n6851;
  assign n6853 = n6625 & n6632;
  assign n6854 = n6619 & n6624;
  assign n6855 = ~n6853 & ~n6854;
  assign n6856 = ~n6852 ^ ~n6855;
  assign n6857 = n6582 & n6597;
  assign n6858 = n6564 & ~n6581;
  assign n6859 = ~n6857 & ~n6858;
  assign n6860 = ~n6856 ^ n6859;
  assign n6861 = ~n6829 ^ n6860;
  assign n6862 = ~n6825 ^ n6861;
  assign n6863 = n6547 & ~n6598;
  assign n6864 = ~n6863 & ~n6603;
  assign n6865 = ~n6547 & n6598;
  assign n6866 = ~n6864 & ~n6865;
  assign n6867 = ~n6862 ^ n6866;
  assign n6868 = ~n6821 ^ n6867;
  assign n6869 = ~n6680 ^ ~n6868;
  assign po065 = n6676 ^ n6869;
  assign n6871 = ~n6670 & ~n6869;
  assign n6872 = ~n6674 & ~n6871;
  assign n6873 = n6471 & ~n6872;
  assign n6874 = ~n6671 & n6869;
  assign n6875 = ~n6668 & ~n6874;
  assign n6876 = ~n6873 & ~n6875;
  assign n6877 = n6821 & ~n6867;
  assign n6878 = n6680 & ~n6877;
  assign n6879 = ~n6821 & n6867;
  assign n6880 = ~n6878 & ~n6879;
  assign n6881 = n6825 & ~n6861;
  assign n6882 = ~n6881 & n6866;
  assign n6883 = ~n6825 & n6861;
  assign n6884 = ~n6882 & ~n6883;
  assign n6885 = ~n6856 & n6859;
  assign n6886 = n6829 & ~n6885;
  assign n6887 = n6856 & ~n6859;
  assign n6888 = ~n6886 & ~n6887;
  assign n6889 = n6852 & n6855;
  assign n6890 = n6840 & ~n6851;
  assign n6891 = ~n6889 & ~n6890;
  assign n6892 = n6836 & n6839;
  assign n6893 = n6832 & n6835;
  assign n6894 = ~n6892 & ~n6893;
  assign n6895 = n6725 & n6728;
  assign n6896 = n6721 & n6724;
  assign n6897 = ~n6895 & ~n6896;
  assign n6898 = ~n6894 ^ ~n6897;
  assign n6899 = n6847 & ~n6850;
  assign n6900 = ~n6843 & ~n6846;
  assign n6901 = ~n6899 & ~n6900;
  assign n6902 = ~n6898 ^ n6901;
  assign n6903 = ~n6891 ^ ~n6902;
  assign n6904 = n6733 & ~n6736;
  assign n6905 = ~n6729 & n6732;
  assign n6906 = ~n6904 & ~n6905;
  assign n6907 = ~n6903 ^ n6906;
  assign n6908 = ~n6694 & ~n6699;
  assign n6909 = ~n6908 & n6697;
  assign n6910 = pi22 & pi43;
  assign n6911 = pi21 & pi44;
  assign n6912 = ~n6910 ^ ~n6911;
  assign n6913 = pi08 & pi57;
  assign n6914 = ~n6912 ^ n6913;
  assign n6915 = pi07 & pi58;
  assign n6916 = pi06 & pi59;
  assign n6917 = ~n6915 ^ ~n6916;
  assign n6918 = pi05 & pi60;
  assign n6919 = ~n6917 ^ n6918;
  assign n6920 = ~n6914 ^ ~n6919;
  assign n6921 = ~n6909 ^ ~n6920;
  assign n6922 = pi29 & pi36;
  assign n6923 = pi19 & pi46;
  assign n6924 = ~n6922 ^ ~n6923;
  assign n6925 = pi11 & pi54;
  assign n6926 = ~n6924 ^ n6925;
  assign n6927 = pi03 & pi62;
  assign n6928 = pi17 & pi48;
  assign n6929 = ~n6927 ^ n6928;
  assign n6930 = ~n6929 ^ pi33;
  assign n6931 = ~n6926 ^ n6930;
  assign n6932 = pi32 & pi33;
  assign n6933 = pi31 & pi34;
  assign n6934 = ~n6932 ^ ~n6933;
  assign n6935 = pi30 & pi35;
  assign n6936 = ~n6934 ^ n6935;
  assign n6937 = ~n6931 ^ ~n6936;
  assign n6938 = ~n6921 ^ n6937;
  assign n6939 = pi28 & pi37;
  assign n6940 = pi27 & pi38;
  assign n6941 = ~n6939 ^ ~n6940;
  assign n6942 = pi26 & pi39;
  assign n6943 = ~n6941 ^ n6942;
  assign n6944 = pi25 & pi40;
  assign n6945 = pi24 & pi41;
  assign n6946 = ~n6944 ^ ~n6945;
  assign n6947 = ~n6946 ^ n3602;
  assign n6948 = ~n6943 ^ ~n6947;
  assign n6949 = pi20 & pi45;
  assign n6950 = pi10 & pi55;
  assign n6951 = ~n6949 ^ ~n6950;
  assign n6952 = pi09 & pi56;
  assign n6953 = ~n6951 ^ n6952;
  assign n6954 = ~n6948 ^ n6953;
  assign n6955 = ~n6938 ^ n6954;
  assign n6956 = ~n6907 ^ ~n6955;
  assign n6957 = ~n6888 ^ ~n6956;
  assign n6958 = ~n6745 & ~n6756;
  assign n6959 = ~n6958 & ~n6760;
  assign n6960 = n6745 & n6756;
  assign n6961 = ~n6959 & ~n6960;
  assign n6962 = n6752 & ~n6755;
  assign n6963 = n6748 & ~n6751;
  assign n6964 = ~n6962 & ~n6963;
  assign n6965 = ~n6771 & n6782;
  assign n6966 = ~n6776 & ~n6781;
  assign n6967 = ~n6965 & ~n6966;
  assign n6968 = n6812 & ~n6813;
  assign n6969 = ~n6810 & ~n6811;
  assign n6970 = ~n6968 & ~n6969;
  assign n6971 = pi02 & pi63;
  assign n6972 = pi04 & pi61;
  assign n6973 = ~n6971 ^ ~n6972;
  assign n6974 = ~n6970 ^ ~n6973;
  assign n6975 = pi18 & pi47;
  assign n6976 = pi13 & pi52;
  assign n6977 = ~n6975 ^ ~n6976;
  assign n6978 = pi12 & pi53;
  assign n6979 = ~n6977 ^ n6978;
  assign n6980 = pi16 & pi49;
  assign n6981 = pi15 & pi50;
  assign n6982 = ~n6980 ^ ~n6981;
  assign n6983 = pi14 & pi51;
  assign n6984 = ~n6982 ^ n6983;
  assign n6985 = ~n6979 ^ ~n6984;
  assign n6986 = ~n6974 ^ ~n6985;
  assign n6987 = ~n6967 ^ n6986;
  assign n6988 = ~n6964 ^ n6987;
  assign n6989 = n6704 & ~n6705;
  assign n6990 = ~n6702 & ~n6703;
  assign n6991 = ~n6989 & ~n6990;
  assign n6992 = n6801 & ~n6802;
  assign n6993 = ~n6799 & ~n6800;
  assign n6994 = ~n6992 & ~n6993;
  assign n6995 = ~n6991 ^ ~n6994;
  assign n6996 = n6795 & ~n6796;
  assign n6997 = ~n3246 & ~n3500;
  assign n6998 = ~n6996 & ~n6997;
  assign n6999 = ~n6995 ^ ~n6998;
  assign n7000 = n6794 & n6797;
  assign n7001 = n6788 & n6793;
  assign n7002 = ~n7000 & ~n7001;
  assign n7003 = ~n6999 ^ ~n7002;
  assign n7004 = n6809 & n6814;
  assign n7005 = n6803 & n6808;
  assign n7006 = ~n7004 & ~n7005;
  assign n7007 = ~n7003 ^ ~n7006;
  assign n7008 = ~n6988 ^ n7007;
  assign n7009 = ~n6961 ^ ~n7008;
  assign n7010 = ~n6957 ^ n7009;
  assign n7011 = ~n6884 ^ n7010;
  assign n7012 = ~n6880 ^ ~n7011;
  assign n7013 = ~n6739 & ~n6819;
  assign n7014 = ~n6684 & ~n7013;
  assign n7015 = n6739 & n6819;
  assign n7016 = ~n7014 & ~n7015;
  assign n7017 = n6718 & ~n6737;
  assign n7018 = ~n6688 & ~n7017;
  assign n7019 = ~n6718 & n6737;
  assign n7020 = ~n7018 & ~n7019;
  assign n7021 = n6714 & ~n6717;
  assign n7022 = ~n6691 & n6713;
  assign n7023 = ~n7021 & ~n7022;
  assign n7024 = n6701 & n6712;
  assign n7025 = ~n6706 & ~n6711;
  assign n7026 = ~n7024 & ~n7025;
  assign n7027 = n6774 & ~n6775;
  assign n7028 = ~n6772 & ~n6773;
  assign n7029 = ~n7027 & ~n7028;
  assign n7030 = n6779 & ~n6780;
  assign n7031 = ~n6777 & ~n6778;
  assign n7032 = ~n7030 & ~n7031;
  assign n7033 = ~n7029 ^ ~n7032;
  assign n7034 = n6806 & ~n6807;
  assign n7035 = ~n6804 & ~n6805;
  assign n7036 = ~n7034 & ~n7035;
  assign n7037 = ~n7033 ^ ~n7036;
  assign n7038 = ~n7026 ^ n7037;
  assign n7039 = n6709 & ~n6710;
  assign n7040 = ~n6707 & ~n6708;
  assign n7041 = ~n7039 & ~n7040;
  assign n7042 = n6786 & ~n6787;
  assign n7043 = ~n6784 & ~n6785;
  assign n7044 = ~n7042 & ~n7043;
  assign n7045 = ~n7041 ^ ~n7044;
  assign n7046 = n6791 & ~n6792;
  assign n7047 = ~n6789 & ~n6790;
  assign n7048 = ~n7046 & ~n7047;
  assign n7049 = ~n7045 ^ ~n7048;
  assign n7050 = ~n7038 ^ ~n7049;
  assign n7051 = n6783 & n6816;
  assign n7052 = ~n6798 & ~n6815;
  assign n7053 = ~n7051 & ~n7052;
  assign n7054 = ~n7050 ^ n7053;
  assign n7055 = ~n7023 ^ n7054;
  assign n7056 = n6761 & ~n6817;
  assign n7057 = n6742 & ~n7056;
  assign n7058 = ~n6761 & n6817;
  assign n7059 = ~n7057 & ~n7058;
  assign n7060 = ~n7055 ^ n7059;
  assign n7061 = ~n7020 ^ ~n7060;
  assign n7062 = ~n7016 ^ n7061;
  assign n7063 = ~n7012 ^ ~n7062;
  assign po066 = n6876 ^ n7063;
  assign n7065 = ~n6880 & ~n7011;
  assign n7066 = n7016 & ~n7061;
  assign n7067 = ~n7065 & n7066;
  assign n7068 = n6880 & n7011;
  assign n7069 = ~n7016 & n7061;
  assign n7070 = n7068 & ~n7069;
  assign n7071 = ~n7067 & ~n7070;
  assign n7072 = ~n6876 & ~n7071;
  assign n7073 = n7065 & n7069;
  assign n7074 = n7068 & n7066;
  assign n7075 = ~n7073 & ~n7074;
  assign n7076 = ~n7072 & n7075;
  assign n7077 = n7065 & ~n7066;
  assign n7078 = ~n7068 & n7069;
  assign n7079 = ~n7077 & ~n7078;
  assign n7080 = n6876 & ~n7079;
  assign n7081 = n7076 & ~n7080;
  assign n7082 = ~n6957 & n7009;
  assign n7083 = ~n6884 & ~n7082;
  assign n7084 = n6957 & ~n7009;
  assign n7085 = ~n7083 & ~n7084;
  assign n7086 = ~n7055 & n7059;
  assign n7087 = n7020 & ~n7086;
  assign n7088 = n7055 & ~n7059;
  assign n7089 = ~n7087 & ~n7088;
  assign n7090 = n6907 & n6955;
  assign n7091 = ~n6888 & ~n7090;
  assign n7092 = ~n6907 & ~n6955;
  assign n7093 = ~n7091 & ~n7092;
  assign n7094 = ~n7050 & n7053;
  assign n7095 = ~n7023 & ~n7094;
  assign n7096 = n7050 & ~n7053;
  assign n7097 = ~n7095 & ~n7096;
  assign n7098 = n7038 & n7049;
  assign n7099 = ~n7026 & n7037;
  assign n7100 = ~n7098 & ~n7099;
  assign n7101 = n7003 & n7006;
  assign n7102 = n6999 & n7002;
  assign n7103 = ~n7101 & ~n7102;
  assign n7104 = n7033 & n7036;
  assign n7105 = n7029 & n7032;
  assign n7106 = ~n7104 & ~n7105;
  assign n7107 = n6995 & n6998;
  assign n7108 = n6991 & n6994;
  assign n7109 = ~n7107 & ~n7108;
  assign n7110 = ~n7106 ^ ~n7109;
  assign n7111 = n7045 & n7048;
  assign n7112 = n7041 & n7044;
  assign n7113 = ~n7111 & ~n7112;
  assign n7114 = ~n7110 ^ ~n7113;
  assign n7115 = ~n7103 ^ ~n7114;
  assign n7116 = ~n7100 ^ n7115;
  assign n7117 = pi18 & pi48;
  assign n7118 = pi15 & pi51;
  assign n7119 = ~n7117 ^ ~n7118;
  assign n7120 = pi13 & pi53;
  assign n7121 = ~n7119 ^ n7120;
  assign n7122 = pi31 & pi35;
  assign n7123 = pi30 & pi36;
  assign n7124 = ~n7122 ^ ~n7123;
  assign n7125 = pi14 & pi52;
  assign n7126 = ~n7124 ^ n7125;
  assign n7127 = ~n7121 ^ ~n7126;
  assign n7128 = pi32 & pi34;
  assign n7129 = pi17 & pi49;
  assign n7130 = ~n7128 ^ ~n7129;
  assign n7131 = pi16 & pi50;
  assign n7132 = ~n7130 ^ n7131;
  assign n7133 = ~n7127 ^ n7132;
  assign n7134 = pi19 & pi47;
  assign n7135 = pi12 & pi54;
  assign n7136 = ~n7134 ^ ~n7135;
  assign n7137 = pi11 & pi55;
  assign n7138 = ~n7136 ^ n7137;
  assign n7139 = pi29 & pi37;
  assign n7140 = pi28 & pi38;
  assign n7141 = ~n7139 ^ ~n7140;
  assign n7142 = pi27 & pi39;
  assign n7143 = ~n7141 ^ n7142;
  assign n7144 = ~n7138 ^ ~n7143;
  assign n7145 = pi05 & pi61;
  assign n7146 = pi04 & pi62;
  assign n7147 = ~n7145 ^ ~n7146;
  assign n7148 = pi03 & pi63;
  assign n7149 = ~n7147 ^ n7148;
  assign n7150 = ~n7144 ^ ~n7149;
  assign n7151 = ~n7133 ^ n7150;
  assign n7152 = pi22 & pi44;
  assign n7153 = pi21 & pi45;
  assign n7154 = ~n7152 ^ ~n7153;
  assign n7155 = pi20 & pi46;
  assign n7156 = ~n7154 ^ n7155;
  assign n7157 = pi26 & pi40;
  assign n7158 = pi25 & pi41;
  assign n7159 = ~n7157 ^ ~n7158;
  assign n7160 = pi10 & pi56;
  assign n7161 = ~n7159 ^ n7160;
  assign n7162 = ~n7156 ^ ~n7161;
  assign n7163 = pi23 & pi43;
  assign n7164 = pi24 & pi42;
  assign n7165 = ~n7163 ^ ~n7164;
  assign n7166 = pi09 & pi57;
  assign n7167 = ~n7165 ^ n7166;
  assign n7168 = ~n7162 ^ n7167;
  assign n7169 = ~n7151 ^ ~n7168;
  assign n7170 = ~n7116 ^ ~n7169;
  assign n7171 = ~n7097 ^ ~n7170;
  assign n7172 = ~n7093 ^ ~n7171;
  assign n7173 = ~n7089 ^ ~n7172;
  assign n7174 = n6961 & ~n7007;
  assign n7175 = ~n7174 & n6988;
  assign n7176 = ~n6961 & n7007;
  assign n7177 = ~n7175 & ~n7176;
  assign n7178 = ~n6967 & n6986;
  assign n7179 = n6964 & ~n7178;
  assign n7180 = n6967 & ~n6986;
  assign n7181 = ~n7179 & ~n7180;
  assign n7182 = n6938 & ~n6954;
  assign n7183 = ~n6921 & n6937;
  assign n7184 = ~n7182 & ~n7183;
  assign n7185 = n6909 & n6920;
  assign n7186 = ~n6914 & ~n6919;
  assign n7187 = ~n7185 & ~n7186;
  assign n7188 = n6948 & ~n6953;
  assign n7189 = ~n6943 & ~n6947;
  assign n7190 = ~n7188 & ~n7189;
  assign n7191 = n6951 & ~n6952;
  assign n7192 = ~n6949 & ~n6950;
  assign n7193 = ~n7191 & ~n7192;
  assign n7194 = n6977 & ~n6978;
  assign n7195 = ~n6975 & ~n6976;
  assign n7196 = ~n7194 & ~n7195;
  assign n7197 = ~n7193 ^ ~n7196;
  assign n7198 = n6946 & ~n3602;
  assign n7199 = ~n6944 & ~n6945;
  assign n7200 = ~n7198 & ~n7199;
  assign n7201 = ~n7197 ^ n7200;
  assign n7202 = ~n7190 ^ ~n7201;
  assign n7203 = ~n7187 ^ n7202;
  assign n7204 = ~n7184 ^ ~n7203;
  assign n7205 = ~n7181 ^ n7204;
  assign n7206 = n6898 & ~n6901;
  assign n7207 = n6894 & n6897;
  assign n7208 = ~n7206 & ~n7207;
  assign n7209 = n6974 & n6985;
  assign n7210 = ~n6979 & ~n6984;
  assign n7211 = ~n7209 & ~n7210;
  assign n7212 = n6970 & n6973;
  assign n7213 = pi04 & pi63;
  assign n7214 = n6589 & n7213;
  assign n7215 = ~n7212 & ~n7214;
  assign n7216 = n6941 & ~n6942;
  assign n7217 = ~n6939 & ~n6940;
  assign n7218 = ~n7216 & ~n7217;
  assign n7219 = pi08 & pi58;
  assign n7220 = pi07 & pi59;
  assign n7221 = ~n7219 ^ ~n7220;
  assign n7222 = pi06 & pi60;
  assign n7223 = ~n7221 ^ n7222;
  assign n7224 = ~n7218 ^ n7223;
  assign n7225 = ~n7215 ^ n7224;
  assign n7226 = ~n7211 ^ n7225;
  assign n7227 = ~n7208 ^ ~n7226;
  assign n7228 = n6982 & ~n6983;
  assign n7229 = ~n6980 & ~n6981;
  assign n7230 = ~n7228 & ~n7229;
  assign n7231 = n6934 & ~n6935;
  assign n7232 = ~n6932 & ~n6933;
  assign n7233 = ~n7231 & ~n7232;
  assign n7234 = ~n7230 ^ ~n7233;
  assign n7235 = n4254 & pi48;
  assign n7236 = ~n7235 & ~n6927;
  assign n7237 = ~n6928 & ~pi33;
  assign n7238 = ~n7236 & ~n7237;
  assign n7239 = ~n7234 ^ ~n7238;
  assign n7240 = n6924 & ~n6925;
  assign n7241 = ~n6922 & ~n6923;
  assign n7242 = ~n7240 & ~n7241;
  assign n7243 = n6912 & ~n6913;
  assign n7244 = ~n6910 & ~n6911;
  assign n7245 = ~n7243 & ~n7244;
  assign n7246 = ~n7242 ^ ~n7245;
  assign n7247 = n6917 & ~n6918;
  assign n7248 = ~n6915 & ~n6916;
  assign n7249 = ~n7247 & ~n7248;
  assign n7250 = ~n7246 ^ n7249;
  assign n7251 = ~n7239 ^ n7250;
  assign n7252 = n6931 & n6936;
  assign n7253 = n6926 & ~n6930;
  assign n7254 = ~n7252 & ~n7253;
  assign n7255 = ~n7251 ^ n7254;
  assign n7256 = ~n7227 ^ n7255;
  assign n7257 = ~n6891 & ~n6902;
  assign n7258 = ~n7257 & ~n6906;
  assign n7259 = n6891 & n6902;
  assign n7260 = ~n7258 & ~n7259;
  assign n7261 = ~n7256 ^ n7260;
  assign n7262 = ~n7205 ^ ~n7261;
  assign n7263 = ~n7177 ^ ~n7262;
  assign n7264 = ~n7173 ^ ~n7263;
  assign n7265 = ~n7085 ^ ~n7264;
  assign po067 = n7081 ^ n7265;
  assign n7267 = ~n7065 & ~n7265;
  assign n7268 = ~n7078 & n7267;
  assign n7269 = ~n7068 & n7265;
  assign n7270 = ~n7269 & n7066;
  assign n7271 = ~n7268 & ~n7270;
  assign n7272 = n6876 & n7271;
  assign n7273 = ~n7267 & n7069;
  assign n7274 = ~n7067 & n7269;
  assign n7275 = ~n7273 & ~n7274;
  assign n7276 = ~n7272 & n7275;
  assign n7277 = n7173 & n7263;
  assign n7278 = n7085 & ~n7277;
  assign n7279 = ~n7173 & ~n7263;
  assign n7280 = ~n7278 & ~n7279;
  assign n7281 = n7093 & n7171;
  assign n7282 = ~n7089 & ~n7281;
  assign n7283 = ~n7093 & ~n7171;
  assign n7284 = ~n7282 & ~n7283;
  assign n7285 = ~n7177 & ~n7261;
  assign n7286 = ~n7285 & n7205;
  assign n7287 = n7177 & n7261;
  assign n7288 = ~n7286 & ~n7287;
  assign n7289 = ~n7116 & ~n7169;
  assign n7290 = ~n7097 & ~n7289;
  assign n7291 = n7116 & n7169;
  assign n7292 = ~n7290 & ~n7291;
  assign n7293 = ~n7184 & ~n7203;
  assign n7294 = n7181 & ~n7293;
  assign n7295 = n7184 & n7203;
  assign n7296 = ~n7294 & ~n7295;
  assign n7297 = ~n7187 & n7202;
  assign n7298 = ~n7190 & ~n7201;
  assign n7299 = ~n7297 & ~n7298;
  assign n7300 = n7197 & ~n7200;
  assign n7301 = ~n7193 & ~n7196;
  assign n7302 = ~n7300 & ~n7301;
  assign n7303 = n7246 & ~n7249;
  assign n7304 = ~n7242 & ~n7245;
  assign n7305 = ~n7303 & ~n7304;
  assign n7306 = ~n7302 ^ ~n7305;
  assign n7307 = n7234 & n7238;
  assign n7308 = n7230 & n7233;
  assign n7309 = ~n7307 & ~n7308;
  assign n7310 = ~n7306 ^ ~n7309;
  assign n7311 = n7251 & ~n7254;
  assign n7312 = ~n7239 & n7250;
  assign n7313 = ~n7311 & ~n7312;
  assign n7314 = ~n7310 ^ n7313;
  assign n7315 = ~n7299 ^ ~n7314;
  assign n7316 = pi26 & pi41;
  assign n7317 = pi25 & pi42;
  assign n7318 = ~n7316 ^ ~n7317;
  assign n7319 = pi21 & pi46;
  assign n7320 = ~n7318 ^ n7319;
  assign n7321 = pi19 & pi48;
  assign n7322 = pi17 & pi50;
  assign n7323 = ~n7321 ^ ~n7322;
  assign n7324 = pi14 & pi53;
  assign n7325 = ~n7323 ^ n7324;
  assign n7326 = ~n7320 ^ ~n7325;
  assign n7327 = pi28 & pi39;
  assign n7328 = pi27 & pi40;
  assign n7329 = ~n7327 ^ ~n7328;
  assign n7330 = ~n7329 ^ n7213;
  assign n7331 = ~n7326 ^ n7330;
  assign n7332 = pi33 & pi34;
  assign n7333 = pi32 & pi35;
  assign n7334 = ~n7332 ^ ~n7333;
  assign n7335 = pi31 & pi36;
  assign n7336 = ~n7334 ^ n7335;
  assign n7337 = pi05 & pi62;
  assign n7338 = pi18 & pi49;
  assign n7339 = ~n7337 ^ n7338;
  assign n7340 = ~n7339 ^ pi34;
  assign n7341 = ~n7336 ^ n7340;
  assign n7342 = pi29 & pi38;
  assign n7343 = pi13 & pi54;
  assign n7344 = ~n7342 ^ ~n7343;
  assign n7345 = pi12 & pi55;
  assign n7346 = ~n7344 ^ n7345;
  assign n7347 = ~n7341 ^ ~n7346;
  assign n7348 = ~n7331 ^ n7347;
  assign n7349 = pi09 & pi58;
  assign n7350 = pi08 & pi59;
  assign n7351 = ~n7349 ^ ~n7350;
  assign n7352 = pi07 & pi60;
  assign n7353 = ~n7351 ^ n7352;
  assign n7354 = pi24 & pi43;
  assign n7355 = ~n3564 ^ ~n7354;
  assign n7356 = pi22 & pi45;
  assign n7357 = ~n7355 ^ n7356;
  assign n7358 = ~n7353 ^ ~n7357;
  assign n7359 = pi30 & pi37;
  assign n7360 = pi16 & pi51;
  assign n7361 = ~n7359 ^ ~n7360;
  assign n7362 = pi15 & pi52;
  assign n7363 = ~n7361 ^ n7362;
  assign n7364 = ~n7358 ^ n7363;
  assign n7365 = ~n7348 ^ ~n7364;
  assign n7366 = ~n7315 ^ n7365;
  assign n7367 = ~n7296 ^ ~n7366;
  assign n7368 = ~n7292 ^ n7367;
  assign n7369 = ~n7288 ^ n7368;
  assign n7370 = ~n7103 & ~n7114;
  assign n7371 = n7100 & ~n7370;
  assign n7372 = n7103 & n7114;
  assign n7373 = ~n7371 & ~n7372;
  assign n7374 = ~n7215 & n7224;
  assign n7375 = n7218 & ~n7223;
  assign n7376 = ~n7374 & ~n7375;
  assign n7377 = n7144 & n7149;
  assign n7378 = n7138 & n7143;
  assign n7379 = ~n7377 & ~n7378;
  assign n7380 = ~n7376 ^ n7379;
  assign n7381 = n7162 & ~n7167;
  assign n7382 = ~n7156 & ~n7161;
  assign n7383 = ~n7381 & ~n7382;
  assign n7384 = ~n7380 ^ n7383;
  assign n7385 = n7141 & ~n7142;
  assign n7386 = ~n7139 & ~n7140;
  assign n7387 = ~n7385 & ~n7386;
  assign n7388 = n7147 & ~n7148;
  assign n7389 = ~n7145 & ~n7146;
  assign n7390 = ~n7388 & ~n7389;
  assign n7391 = ~n7387 ^ ~n7390;
  assign n7392 = n7221 & ~n7222;
  assign n7393 = ~n7219 & ~n7220;
  assign n7394 = ~n7392 & ~n7393;
  assign n7395 = ~n7391 ^ ~n7394;
  assign n7396 = n7130 & ~n7131;
  assign n7397 = ~n7128 & ~n7129;
  assign n7398 = ~n7396 & ~n7397;
  assign n7399 = pi06 & pi61;
  assign n7400 = ~n7398 ^ ~n7399;
  assign n7401 = n7124 & ~n7125;
  assign n7402 = ~n7122 & ~n7123;
  assign n7403 = ~n7401 & ~n7402;
  assign n7404 = ~n7400 ^ ~n7403;
  assign n7405 = ~n7395 ^ ~n7404;
  assign n7406 = n7154 & ~n7155;
  assign n7407 = ~n7152 & ~n7153;
  assign n7408 = ~n7406 & ~n7407;
  assign n7409 = n7165 & ~n7166;
  assign n7410 = ~n7163 & ~n7164;
  assign n7411 = ~n7409 & ~n7410;
  assign n7412 = ~n7408 ^ ~n7411;
  assign n7413 = n7159 & ~n7160;
  assign n7414 = ~n7157 & ~n7158;
  assign n7415 = ~n7413 & ~n7414;
  assign n7416 = ~n7412 ^ ~n7415;
  assign n7417 = ~n7405 ^ ~n7416;
  assign n7418 = ~n7384 ^ ~n7417;
  assign n7419 = ~n7373 ^ ~n7418;
  assign n7420 = n7110 & n7113;
  assign n7421 = n7106 & n7109;
  assign n7422 = ~n7420 & ~n7421;
  assign n7423 = n7127 & ~n7132;
  assign n7424 = ~n7121 & ~n7126;
  assign n7425 = ~n7423 & ~n7424;
  assign n7426 = n7136 & ~n7137;
  assign n7427 = ~n7134 & ~n7135;
  assign n7428 = ~n7426 & ~n7427;
  assign n7429 = pi20 & pi47;
  assign n7430 = pi11 & pi56;
  assign n7431 = ~n7429 ^ ~n7430;
  assign n7432 = pi10 & pi57;
  assign n7433 = ~n7431 ^ n7432;
  assign n7434 = ~n7428 ^ n7433;
  assign n7435 = n7119 & ~n7120;
  assign n7436 = ~n7117 & ~n7118;
  assign n7437 = ~n7435 & ~n7436;
  assign n7438 = ~n7434 ^ ~n7437;
  assign n7439 = ~n7425 ^ n7438;
  assign n7440 = ~n7422 ^ ~n7439;
  assign n7441 = n7151 & n7168;
  assign n7442 = n7133 & ~n7150;
  assign n7443 = ~n7441 & ~n7442;
  assign n7444 = ~n7440 ^ n7443;
  assign n7445 = n7211 & ~n7225;
  assign n7446 = n7208 & ~n7445;
  assign n7447 = ~n7211 & n7225;
  assign n7448 = ~n7446 & ~n7447;
  assign n7449 = ~n7444 ^ n7448;
  assign n7450 = ~n7419 ^ ~n7449;
  assign n7451 = n7227 & ~n7255;
  assign n7452 = ~n7451 & ~n7260;
  assign n7453 = ~n7227 & n7255;
  assign n7454 = ~n7452 & ~n7453;
  assign n7455 = ~n7450 ^ ~n7454;
  assign n7456 = ~n7369 ^ ~n7455;
  assign n7457 = ~n7284 ^ ~n7456;
  assign n7458 = ~n7280 ^ ~n7457;
  assign po068 = n7276 ^ ~n7458;
  assign n7460 = n7280 & n7457;
  assign n7461 = ~n7276 & ~n7460;
  assign n7462 = ~n7280 & ~n7457;
  assign n7463 = ~n7461 & ~n7462;
  assign n7464 = n7369 & n7455;
  assign n7465 = n7284 & ~n7464;
  assign n7466 = ~n7369 & ~n7455;
  assign n7467 = ~n7465 & ~n7466;
  assign n7468 = n7288 & ~n7367;
  assign n7469 = ~n7468 & n7292;
  assign n7470 = ~n7288 & n7367;
  assign n7471 = ~n7469 & ~n7470;
  assign n7472 = ~n7315 & n7365;
  assign n7473 = n7296 & ~n7472;
  assign n7474 = n7315 & ~n7365;
  assign n7475 = ~n7473 & ~n7474;
  assign n7476 = n7380 & ~n7383;
  assign n7477 = ~n7376 & n7379;
  assign n7478 = ~n7476 & ~n7477;
  assign n7479 = n7405 & n7416;
  assign n7480 = n7395 & n7404;
  assign n7481 = ~n7479 & ~n7480;
  assign n7482 = ~n7478 ^ ~n7481;
  assign n7483 = ~n7425 & n7438;
  assign n7484 = ~n7422 & ~n7483;
  assign n7485 = n7425 & ~n7438;
  assign n7486 = ~n7484 & ~n7485;
  assign n7487 = ~n7482 ^ ~n7486;
  assign n7488 = pi33 & pi35;
  assign n7489 = pi19 & pi49;
  assign n7490 = ~n7488 ^ ~n7489;
  assign n7491 = pi18 & pi50;
  assign n7492 = ~n7490 ^ n7491;
  assign n7493 = pi17 & pi51;
  assign n7494 = pi13 & pi55;
  assign n7495 = ~n7493 ^ ~n7494;
  assign n7496 = pi12 & pi56;
  assign n7497 = ~n7495 ^ n7496;
  assign n7498 = ~n7492 ^ ~n7497;
  assign n7499 = pi32 & pi36;
  assign n7500 = pi31 & pi37;
  assign n7501 = ~n7499 ^ ~n7500;
  assign n7502 = pi30 & pi38;
  assign n7503 = ~n7501 ^ n7502;
  assign n7504 = ~n7498 ^ n7503;
  assign n7505 = pi16 & pi52;
  assign n7506 = pi15 & pi53;
  assign n7507 = ~n7505 ^ ~n7506;
  assign n7508 = pi14 & pi54;
  assign n7509 = ~n7507 ^ n7508;
  assign n7510 = pi26 & pi42;
  assign n7511 = pi25 & pi43;
  assign n7512 = ~n7510 ^ ~n7511;
  assign n7513 = pi24 & pi44;
  assign n7514 = ~n7512 ^ n7513;
  assign n7515 = ~n7509 ^ ~n7514;
  assign n7516 = pi23 & pi45;
  assign n7517 = pi22 & pi46;
  assign n7518 = ~n7516 ^ ~n7517;
  assign n7519 = pi20 & pi48;
  assign n7520 = ~n7518 ^ n7519;
  assign n7521 = ~n7515 ^ ~n7520;
  assign n7522 = ~n7504 ^ n7521;
  assign n7523 = pi29 & pi39;
  assign n7524 = pi28 & pi40;
  assign n7525 = ~n7523 ^ ~n7524;
  assign n7526 = pi27 & pi41;
  assign n7527 = ~n7525 ^ n7526;
  assign n7528 = pi21 & pi47;
  assign n7529 = pi06 & pi62;
  assign n7530 = ~n7528 ^ ~n7529;
  assign n7531 = pi05 & pi63;
  assign n7532 = ~n7530 ^ n7531;
  assign n7533 = ~n7527 ^ ~n7532;
  assign n7534 = pi11 & pi57;
  assign n7535 = pi10 & pi58;
  assign n7536 = ~n7534 ^ ~n7535;
  assign n7537 = pi09 & pi59;
  assign n7538 = ~n7536 ^ n7537;
  assign n7539 = ~n7533 ^ n7538;
  assign n7540 = ~n7522 ^ ~n7539;
  assign n7541 = ~n7487 ^ ~n7540;
  assign n7542 = ~n7440 & n7443;
  assign n7543 = ~n7542 & ~n7448;
  assign n7544 = n7440 & ~n7443;
  assign n7545 = ~n7543 & ~n7544;
  assign n7546 = ~n7541 ^ ~n7545;
  assign n7547 = ~n7475 ^ ~n7546;
  assign n7548 = ~n7419 & ~n7449;
  assign n7549 = ~n7548 & n7454;
  assign n7550 = n7419 & n7449;
  assign n7551 = ~n7549 & ~n7550;
  assign n7552 = ~n7547 ^ n7551;
  assign n7553 = n7384 & n7417;
  assign n7554 = ~n7373 & ~n7553;
  assign n7555 = ~n7384 & ~n7417;
  assign n7556 = ~n7554 & ~n7555;
  assign n7557 = n7299 & n7314;
  assign n7558 = n7310 & ~n7313;
  assign n7559 = ~n7557 & ~n7558;
  assign n7560 = n7306 & n7309;
  assign n7561 = ~n7302 & ~n7305;
  assign n7562 = ~n7560 & ~n7561;
  assign n7563 = n7351 & ~n7352;
  assign n7564 = ~n7349 & ~n7350;
  assign n7565 = ~n7563 & ~n7564;
  assign n7566 = n7355 & ~n7356;
  assign n7567 = ~n3564 & ~n7354;
  assign n7568 = ~n7566 & ~n7567;
  assign n7569 = ~n7565 ^ ~n7568;
  assign n7570 = n7431 & ~n7432;
  assign n7571 = ~n7429 & ~n7430;
  assign n7572 = ~n7570 & ~n7571;
  assign n7573 = ~n7569 ^ ~n7572;
  assign n7574 = n7361 & ~n7362;
  assign n7575 = ~n7359 & ~n7360;
  assign n7576 = ~n7574 & ~n7575;
  assign n7577 = n7334 & ~n7335;
  assign n7578 = ~n7332 & ~n7333;
  assign n7579 = ~n7577 & ~n7578;
  assign n7580 = ~n7576 ^ ~n7579;
  assign n7581 = n7329 & ~n7213;
  assign n7582 = ~n7327 & ~n7328;
  assign n7583 = ~n7581 & ~n7582;
  assign n7584 = ~n7580 ^ n7583;
  assign n7585 = ~n7573 ^ n7584;
  assign n7586 = ~n7562 ^ n7585;
  assign n7587 = n7344 & ~n7345;
  assign n7588 = ~n7342 & ~n7343;
  assign n7589 = ~n7587 & ~n7588;
  assign n7590 = n7318 & ~n7319;
  assign n7591 = ~n7316 & ~n7317;
  assign n7592 = ~n7590 & ~n7591;
  assign n7593 = ~n7589 ^ ~n7592;
  assign n7594 = n7323 & ~n7324;
  assign n7595 = ~n7321 & ~n7322;
  assign n7596 = ~n7594 & ~n7595;
  assign n7597 = ~n7593 ^ ~n7596;
  assign n7598 = n7341 & n7346;
  assign n7599 = n7336 & ~n7340;
  assign n7600 = ~n7598 & ~n7599;
  assign n7601 = ~n7597 ^ ~n7600;
  assign n7602 = n7326 & ~n7330;
  assign n7603 = ~n7320 & ~n7325;
  assign n7604 = ~n7602 & ~n7603;
  assign n7605 = ~n7601 ^ ~n7604;
  assign n7606 = ~n7586 ^ ~n7605;
  assign n7607 = ~n7559 ^ ~n7606;
  assign n7608 = n7434 & n7437;
  assign n7609 = n7428 & ~n7433;
  assign n7610 = ~n7608 & ~n7609;
  assign n7611 = n7358 & ~n7363;
  assign n7612 = ~n7353 & ~n7357;
  assign n7613 = ~n7611 & ~n7612;
  assign n7614 = ~n7610 ^ ~n7613;
  assign n7615 = n7412 & n7415;
  assign n7616 = n7408 & n7411;
  assign n7617 = ~n7615 & ~n7616;
  assign n7618 = ~n7614 ^ n7617;
  assign n7619 = n7348 & n7364;
  assign n7620 = n7331 & ~n7347;
  assign n7621 = ~n7619 & ~n7620;
  assign n7622 = ~n7618 ^ n7621;
  assign n7623 = n7391 & n7394;
  assign n7624 = n7387 & n7390;
  assign n7625 = ~n7623 & ~n7624;
  assign n7626 = n4601 & pi49;
  assign n7627 = ~n7626 & ~n7337;
  assign n7628 = ~n7338 & ~pi34;
  assign n7629 = ~n7627 & ~n7628;
  assign n7630 = pi07 & pi61;
  assign n7631 = pi08 & pi60;
  assign n7632 = ~n7630 ^ ~n7631;
  assign n7633 = ~n7629 ^ ~n7632;
  assign n7634 = ~n7625 ^ n7633;
  assign n7635 = n7400 & n7403;
  assign n7636 = n7398 & n7399;
  assign n7637 = ~n7635 & ~n7636;
  assign n7638 = ~n7634 ^ n7637;
  assign n7639 = ~n7622 ^ n7638;
  assign n7640 = ~n7607 ^ n7639;
  assign n7641 = ~n7556 ^ n7640;
  assign n7642 = ~n7552 ^ ~n7641;
  assign n7643 = ~n7471 ^ n7642;
  assign n7644 = ~n7467 ^ ~n7643;
  assign po069 = ~n7463 ^ ~n7644;
  assign n7646 = n7552 & n7641;
  assign n7647 = ~n7471 & n7646;
  assign n7648 = ~n7467 & n7647;
  assign n7649 = ~n7463 & ~n7648;
  assign n7650 = ~n7552 & ~n7641;
  assign n7651 = ~n7471 & ~n7650;
  assign n7652 = ~n7651 & ~n7646;
  assign n7653 = ~n7467 & ~n7652;
  assign n7654 = ~n7653 & ~n7647;
  assign n7655 = ~n7649 & ~n7654;
  assign n7656 = n7471 & n7650;
  assign n7657 = ~n7467 & ~n7656;
  assign n7658 = ~n7657 & n7652;
  assign n7659 = ~n7463 & n7658;
  assign n7660 = n7467 & n7656;
  assign n7661 = ~n7659 & ~n7660;
  assign n7662 = ~n7655 & n7661;
  assign n7663 = ~n7551 & ~n7546;
  assign n7664 = ~n7663 & ~n7475;
  assign n7665 = n7551 & n7546;
  assign n7666 = ~n7664 & ~n7665;
  assign n7667 = ~n7586 & ~n7605;
  assign n7668 = ~n7559 & ~n7667;
  assign n7669 = n7586 & n7605;
  assign n7670 = ~n7668 & ~n7669;
  assign n7671 = n7573 & ~n7584;
  assign n7672 = ~n7562 & ~n7671;
  assign n7673 = ~n7573 & n7584;
  assign n7674 = ~n7672 & ~n7673;
  assign n7675 = n7593 & n7596;
  assign n7676 = n7589 & n7592;
  assign n7677 = ~n7675 & ~n7676;
  assign n7678 = n7580 & ~n7583;
  assign n7679 = ~n7576 & ~n7579;
  assign n7680 = ~n7678 & ~n7679;
  assign n7681 = ~n7677 ^ n7680;
  assign n7682 = n7525 & ~n7526;
  assign n7683 = ~n7523 & ~n7524;
  assign n7684 = ~n7682 & ~n7683;
  assign n7685 = n7495 & ~n7496;
  assign n7686 = ~n7493 & ~n7494;
  assign n7687 = ~n7685 & ~n7686;
  assign n7688 = ~n7684 ^ ~n7687;
  assign n7689 = n7512 & ~n7513;
  assign n7690 = ~n7510 & ~n7511;
  assign n7691 = ~n7689 & ~n7690;
  assign n7692 = ~n7688 ^ ~n7691;
  assign n7693 = ~n7681 ^ ~n7692;
  assign n7694 = n7522 & n7539;
  assign n7695 = n7504 & ~n7521;
  assign n7696 = ~n7694 & ~n7695;
  assign n7697 = ~n7693 ^ n7696;
  assign n7698 = ~n7674 ^ n7697;
  assign n7699 = ~n7670 ^ n7698;
  assign n7700 = ~n7478 & ~n7481;
  assign n7701 = ~n7700 & ~n7486;
  assign n7702 = n7478 & n7481;
  assign n7703 = ~n7701 & ~n7702;
  assign n7704 = n7634 & ~n7637;
  assign n7705 = ~n7625 & n7633;
  assign n7706 = ~n7704 & ~n7705;
  assign n7707 = n7498 & ~n7503;
  assign n7708 = ~n7492 & ~n7497;
  assign n7709 = ~n7707 & ~n7708;
  assign n7710 = n7515 & n7520;
  assign n7711 = n7509 & n7514;
  assign n7712 = ~n7710 & ~n7711;
  assign n7713 = ~n7709 ^ n7712;
  assign n7714 = ~n7706 ^ n7713;
  assign n7715 = n7530 & ~n7531;
  assign n7716 = ~n7528 & ~n7529;
  assign n7717 = ~n7715 & ~n7716;
  assign n7718 = n7536 & ~n7537;
  assign n7719 = ~n7534 & ~n7535;
  assign n7720 = ~n7718 & ~n7719;
  assign n7721 = ~n7717 ^ ~n7720;
  assign n7722 = n7518 & ~n7519;
  assign n7723 = ~n7516 & ~n7517;
  assign n7724 = ~n7722 & ~n7723;
  assign n7725 = ~n7721 ^ ~n7724;
  assign n7726 = n7501 & ~n7502;
  assign n7727 = ~n7499 & ~n7500;
  assign n7728 = ~n7726 & ~n7727;
  assign n7729 = n7490 & ~n7491;
  assign n7730 = ~n7488 & ~n7489;
  assign n7731 = ~n7729 & ~n7730;
  assign n7732 = ~n7728 ^ ~n7731;
  assign n7733 = n7507 & ~n7508;
  assign n7734 = ~n7505 & ~n7506;
  assign n7735 = ~n7733 & ~n7734;
  assign n7736 = ~n7732 ^ n7735;
  assign n7737 = ~n7725 ^ n7736;
  assign n7738 = n7533 & ~n7538;
  assign n7739 = ~n7527 & ~n7532;
  assign n7740 = ~n7738 & ~n7739;
  assign n7741 = ~n7737 ^ ~n7740;
  assign n7742 = ~n7714 ^ n7741;
  assign n7743 = ~n7703 ^ ~n7742;
  assign n7744 = ~n7699 ^ n7743;
  assign n7745 = ~n7666 ^ n7744;
  assign n7746 = ~n7487 & ~n7540;
  assign n7747 = ~n7746 & ~n7545;
  assign n7748 = n7487 & n7540;
  assign n7749 = ~n7747 & ~n7748;
  assign n7750 = n7614 & ~n7617;
  assign n7751 = ~n7610 & ~n7613;
  assign n7752 = ~n7750 & ~n7751;
  assign n7753 = pi10 & pi59;
  assign n7754 = pi09 & pi60;
  assign n7755 = ~n7753 ^ ~n7754;
  assign n7756 = pi08 & pi61;
  assign n7757 = ~n7755 ^ n7756;
  assign n7758 = pi25 & pi44;
  assign n7759 = pi24 & pi45;
  assign n7760 = ~n7758 ^ ~n7759;
  assign n7761 = pi23 & pi46;
  assign n7762 = ~n7760 ^ n7761;
  assign n7763 = ~n7757 ^ ~n7762;
  assign n7764 = pi27 & pi42;
  assign n7765 = pi26 & pi43;
  assign n7766 = ~n7764 ^ ~n7765;
  assign n7767 = pi06 & pi63;
  assign n7768 = ~n7766 ^ n7767;
  assign n7769 = ~n7763 ^ ~n7768;
  assign n7770 = ~n7752 ^ ~n7769;
  assign n7771 = n7629 & n7632;
  assign n7772 = pi60 & pi61;
  assign n7773 = n559 & n7772;
  assign n7774 = ~n7771 & ~n7773;
  assign n7775 = pi22 & pi47;
  assign n7776 = pi21 & pi48;
  assign n7777 = ~n7775 ^ ~n7776;
  assign n7778 = pi14 & pi55;
  assign n7779 = ~n7777 ^ n7778;
  assign n7780 = pi13 & pi56;
  assign n7781 = pi12 & pi57;
  assign n7782 = ~n7780 ^ ~n7781;
  assign n7783 = pi11 & pi58;
  assign n7784 = ~n7782 ^ n7783;
  assign n7785 = ~n7779 ^ ~n7784;
  assign n7786 = ~n7774 ^ n7785;
  assign n7787 = ~n7770 ^ ~n7786;
  assign n7788 = n7601 & n7604;
  assign n7789 = ~n7597 & ~n7600;
  assign n7790 = ~n7788 & ~n7789;
  assign n7791 = n7569 & n7572;
  assign n7792 = n7565 & n7568;
  assign n7793 = ~n7791 & ~n7792;
  assign n7794 = pi30 & pi39;
  assign n7795 = pi29 & pi40;
  assign n7796 = ~n7794 ^ ~n7795;
  assign n7797 = pi28 & pi41;
  assign n7798 = ~n7796 ^ n7797;
  assign n7799 = pi19 & pi50;
  assign n7800 = pi18 & pi51;
  assign n7801 = ~n7799 ^ ~n7800;
  assign n7802 = pi17 & pi52;
  assign n7803 = ~n7801 ^ n7802;
  assign n7804 = ~n7798 ^ ~n7803;
  assign n7805 = ~n7793 ^ ~n7804;
  assign n7806 = pi20 & pi49;
  assign n7807 = pi16 & pi53;
  assign n7808 = ~n7806 ^ ~n7807;
  assign n7809 = pi15 & pi54;
  assign n7810 = ~n7808 ^ n7809;
  assign n7811 = pi33 & pi36;
  assign n7812 = pi32 & pi37;
  assign n7813 = ~n7811 ^ ~n7812;
  assign n7814 = pi31 & pi38;
  assign n7815 = ~n7813 ^ n7814;
  assign n7816 = ~n7810 ^ ~n7815;
  assign n7817 = pi07 & pi62;
  assign n7818 = ~pi34 & pi35;
  assign n7819 = ~n7817 ^ ~n7818;
  assign n7820 = ~n7816 ^ ~n7819;
  assign n7821 = ~n7805 ^ n7820;
  assign n7822 = ~n7790 ^ ~n7821;
  assign n7823 = ~n7787 ^ ~n7822;
  assign n7824 = n7622 & ~n7638;
  assign n7825 = ~n7618 & n7621;
  assign n7826 = ~n7824 & ~n7825;
  assign n7827 = ~n7823 ^ ~n7826;
  assign n7828 = ~n7749 ^ n7827;
  assign n7829 = ~n7607 & n7639;
  assign n7830 = n7556 & ~n7829;
  assign n7831 = n7607 & ~n7639;
  assign n7832 = ~n7830 & ~n7831;
  assign n7833 = ~n7828 ^ ~n7832;
  assign n7834 = ~n7745 ^ n7833;
  assign po070 = ~n7662 ^ ~n7834;
  assign n7836 = ~n7660 & ~n7834;
  assign n7837 = n7654 & ~n7836;
  assign n7838 = n7463 & ~n7837;
  assign n7839 = ~n7658 & ~n7834;
  assign n7840 = ~n7839 & ~n7648;
  assign n7841 = ~n7838 & n7840;
  assign n7842 = n7666 & ~n7744;
  assign n7843 = ~n7842 & n7833;
  assign n7844 = ~n7666 & n7744;
  assign n7845 = ~n7843 & ~n7844;
  assign n7846 = ~n7832 & n7827;
  assign n7847 = ~n7846 & n7749;
  assign n7848 = n7832 & ~n7827;
  assign n7849 = ~n7847 & ~n7848;
  assign n7850 = ~n7670 & n7698;
  assign n7851 = ~n7850 & n7743;
  assign n7852 = n7670 & ~n7698;
  assign n7853 = ~n7851 & ~n7852;
  assign n7854 = n7693 & ~n7696;
  assign n7855 = ~n7674 & ~n7854;
  assign n7856 = ~n7693 & n7696;
  assign n7857 = ~n7855 & ~n7856;
  assign n7858 = n7681 & n7692;
  assign n7859 = ~n7677 & n7680;
  assign n7860 = ~n7858 & ~n7859;
  assign n7861 = n7801 & ~n7802;
  assign n7862 = ~n7799 & ~n7800;
  assign n7863 = ~n7861 & ~n7862;
  assign n7864 = n7808 & ~n7809;
  assign n7865 = ~n7806 & ~n7807;
  assign n7866 = ~n7864 & ~n7865;
  assign n7867 = ~n7863 ^ ~n7866;
  assign n7868 = pi34 & pi36;
  assign n7869 = pi33 & pi37;
  assign n7870 = ~n7868 ^ ~n7869;
  assign n7871 = pi32 & pi38;
  assign n7872 = ~n7870 ^ n7871;
  assign n7873 = ~n7867 ^ n7872;
  assign n7874 = ~n7860 ^ n7873;
  assign n7875 = pi11 & pi59;
  assign n7876 = pi10 & pi60;
  assign n7877 = ~n7875 ^ ~n7876;
  assign n7878 = pi09 & pi61;
  assign n7879 = ~n7877 ^ n7878;
  assign n7880 = pi18 & pi52;
  assign n7881 = pi17 & pi53;
  assign n7882 = ~n7880 ^ ~n7881;
  assign n7883 = pi16 & pi54;
  assign n7884 = ~n7882 ^ n7883;
  assign n7885 = ~n7879 ^ ~n7884;
  assign n7886 = pi24 & pi46;
  assign n7887 = pi13 & pi57;
  assign n7888 = ~n7886 ^ ~n7887;
  assign n7889 = pi12 & pi58;
  assign n7890 = ~n7888 ^ n7889;
  assign n7891 = ~n7885 ^ n7890;
  assign n7892 = ~n7874 ^ ~n7891;
  assign n7893 = n7737 & n7740;
  assign n7894 = ~n7725 & n7736;
  assign n7895 = ~n7893 & ~n7894;
  assign n7896 = n7732 & ~n7735;
  assign n7897 = ~n7728 & ~n7731;
  assign n7898 = ~n7896 & ~n7897;
  assign n7899 = pi28 & pi42;
  assign n7900 = ~n4009 ^ ~n7899;
  assign n7901 = pi07 & pi63;
  assign n7902 = ~n7900 ^ n7901;
  assign n7903 = pi31 & pi39;
  assign n7904 = pi30 & pi40;
  assign n7905 = ~n7903 ^ ~n7904;
  assign n7906 = pi29 & pi41;
  assign n7907 = ~n7905 ^ n7906;
  assign n7908 = ~n7902 ^ ~n7907;
  assign n7909 = ~n7898 ^ ~n7908;
  assign n7910 = pi27 & pi43;
  assign n7911 = pi26 & pi44;
  assign n7912 = ~n7910 ^ ~n7911;
  assign n7913 = pi25 & pi45;
  assign n7914 = ~n7912 ^ n7913;
  assign n7915 = pi21 & pi49;
  assign n7916 = pi20 & pi50;
  assign n7917 = ~n7915 ^ ~n7916;
  assign n7918 = pi19 & pi51;
  assign n7919 = ~n7917 ^ n7918;
  assign n7920 = ~n7914 ^ ~n7919;
  assign n7921 = pi22 & pi48;
  assign n7922 = pi15 & pi55;
  assign n7923 = ~n7921 ^ ~n7922;
  assign n7924 = pi14 & pi56;
  assign n7925 = ~n7923 ^ n7924;
  assign n7926 = ~n7920 ^ n7925;
  assign n7927 = ~n7909 ^ ~n7926;
  assign n7928 = ~n7895 ^ ~n7927;
  assign n7929 = ~n7892 ^ ~n7928;
  assign n7930 = ~n7857 ^ n7929;
  assign n7931 = n7793 & n7804;
  assign n7932 = n7798 & n7803;
  assign n7933 = ~n7931 & ~n7932;
  assign n7934 = n7813 & ~n7814;
  assign n7935 = ~n7811 & ~n7812;
  assign n7936 = ~n7934 & ~n7935;
  assign n7937 = ~n7817 & ~pi34;
  assign n7938 = ~n7937 & pi35;
  assign n7939 = pi08 & pi62;
  assign n7940 = ~n7938 ^ ~n7939;
  assign n7941 = ~n7936 ^ n7940;
  assign n7942 = ~n7933 ^ n7941;
  assign n7943 = n7760 & ~n7761;
  assign n7944 = ~n7758 & ~n7759;
  assign n7945 = ~n7943 & ~n7944;
  assign n7946 = n7766 & ~n7767;
  assign n7947 = ~n7764 & ~n7765;
  assign n7948 = ~n7946 & ~n7947;
  assign n7949 = ~n7945 ^ ~n7948;
  assign n7950 = n7796 & ~n7797;
  assign n7951 = ~n7794 & ~n7795;
  assign n7952 = ~n7950 & ~n7951;
  assign n7953 = ~n7949 ^ ~n7952;
  assign n7954 = ~n7942 ^ n7953;
  assign n7955 = ~n7774 & n7785;
  assign n7956 = ~n7779 & ~n7784;
  assign n7957 = ~n7955 & ~n7956;
  assign n7958 = n7763 & n7768;
  assign n7959 = n7757 & n7762;
  assign n7960 = ~n7958 & ~n7959;
  assign n7961 = n7816 & n7819;
  assign n7962 = ~n7810 & ~n7815;
  assign n7963 = ~n7961 & ~n7962;
  assign n7964 = ~n7960 ^ n7963;
  assign n7965 = ~n7957 ^ n7964;
  assign n7966 = ~n7954 ^ n7965;
  assign n7967 = n7790 & n7821;
  assign n7968 = ~n7805 & n7820;
  assign n7969 = ~n7967 & ~n7968;
  assign n7970 = ~n7966 ^ ~n7969;
  assign n7971 = ~n7930 ^ ~n7970;
  assign n7972 = ~n7853 ^ ~n7971;
  assign n7973 = n7787 & n7822;
  assign n7974 = ~n7973 & ~n7826;
  assign n7975 = ~n7787 & ~n7822;
  assign n7976 = ~n7974 & ~n7975;
  assign n7977 = n7770 & n7786;
  assign n7978 = ~n7752 & ~n7769;
  assign n7979 = ~n7977 & ~n7978;
  assign n7980 = ~n7706 & n7713;
  assign n7981 = ~n7709 & n7712;
  assign n7982 = ~n7980 & ~n7981;
  assign n7983 = n7688 & n7691;
  assign n7984 = n7684 & n7687;
  assign n7985 = ~n7983 & ~n7984;
  assign n7986 = n7721 & n7724;
  assign n7987 = n7717 & n7720;
  assign n7988 = ~n7986 & ~n7987;
  assign n7989 = ~n7985 ^ ~n7988;
  assign n7990 = n7782 & ~n7783;
  assign n7991 = ~n7780 & ~n7781;
  assign n7992 = ~n7990 & ~n7991;
  assign n7993 = n7777 & ~n7778;
  assign n7994 = ~n7775 & ~n7776;
  assign n7995 = ~n7993 & ~n7994;
  assign n7996 = ~n7992 ^ ~n7995;
  assign n7997 = n7755 & ~n7756;
  assign n7998 = ~n7753 & ~n7754;
  assign n7999 = ~n7997 & ~n7998;
  assign n8000 = ~n7996 ^ ~n7999;
  assign n8001 = ~n7989 ^ n8000;
  assign n8002 = ~n7982 ^ ~n8001;
  assign n8003 = ~n7979 ^ n8002;
  assign n8004 = ~n7976 ^ ~n8003;
  assign n8005 = ~n7714 & n7741;
  assign n8006 = n7703 & ~n8005;
  assign n8007 = n7714 & ~n7741;
  assign n8008 = ~n8006 & ~n8007;
  assign n8009 = ~n8004 ^ ~n8008;
  assign n8010 = ~n7972 ^ ~n8009;
  assign n8011 = ~n7849 ^ ~n8010;
  assign n8012 = ~n7845 ^ ~n8011;
  assign po071 = ~n7841 ^ ~n8012;
  assign n8014 = ~n7845 & ~n8011;
  assign n8015 = n7841 & ~n8014;
  assign n8016 = n7845 & n8011;
  assign n8017 = ~n8015 & ~n8016;
  assign n8018 = n7972 & n8009;
  assign n8019 = n7849 & ~n8018;
  assign n8020 = ~n7972 & ~n8009;
  assign n8021 = ~n8019 & ~n8020;
  assign n8022 = ~n7930 & ~n7970;
  assign n8023 = n7853 & ~n8022;
  assign n8024 = n7930 & n7970;
  assign n8025 = ~n8023 & ~n8024;
  assign n8026 = n7892 & n7928;
  assign n8027 = ~n7857 & ~n8026;
  assign n8028 = ~n7892 & ~n7928;
  assign n8029 = ~n8027 & ~n8028;
  assign n8030 = n7966 & n7969;
  assign n8031 = n7954 & ~n7965;
  assign n8032 = ~n8030 & ~n8031;
  assign n8033 = n7874 & n7891;
  assign n8034 = ~n7860 & n7873;
  assign n8035 = ~n8033 & ~n8034;
  assign n8036 = n7942 & ~n7953;
  assign n8037 = ~n7933 & n7941;
  assign n8038 = ~n8036 & ~n8037;
  assign n8039 = n7949 & n7952;
  assign n8040 = n7945 & n7948;
  assign n8041 = ~n8039 & ~n8040;
  assign n8042 = ~n7936 & n7940;
  assign n8043 = ~n7938 & ~n7939;
  assign n8044 = ~n8042 & ~n8043;
  assign n8045 = ~n8041 ^ n8044;
  assign n8046 = n7867 & ~n7872;
  assign n8047 = n7863 & n7866;
  assign n8048 = ~n8046 & ~n8047;
  assign n8049 = ~n8045 ^ n8048;
  assign n8050 = ~n8038 ^ ~n8049;
  assign n8051 = ~n8035 ^ n8050;
  assign n8052 = ~n8032 ^ ~n8051;
  assign n8053 = ~n8029 ^ n8052;
  assign n8054 = ~n8025 ^ ~n8053;
  assign n8055 = n7976 & n8003;
  assign n8056 = ~n8055 & n8008;
  assign n8057 = ~n7976 & ~n8003;
  assign n8058 = ~n8056 & ~n8057;
  assign n8059 = ~n7982 & ~n8001;
  assign n8060 = n7979 & ~n8059;
  assign n8061 = n7982 & n8001;
  assign n8062 = ~n8060 & ~n8061;
  assign n8063 = ~n7957 & n7964;
  assign n8064 = n7960 & ~n7963;
  assign n8065 = ~n8063 & ~n8064;
  assign n8066 = n7917 & ~n7918;
  assign n8067 = ~n7915 & ~n7916;
  assign n8068 = ~n8066 & ~n8067;
  assign n8069 = pi12 & pi59;
  assign n8070 = pi13 & pi58;
  assign n8071 = ~n8069 ^ ~n8070;
  assign n8072 = ~n8068 ^ ~n8071;
  assign n8073 = pi16 & pi55;
  assign n8074 = pi15 & pi56;
  assign n8075 = ~n8073 ^ ~n8074;
  assign n8076 = pi14 & pi57;
  assign n8077 = ~n8075 ^ n8076;
  assign n8078 = pi26 & pi45;
  assign n8079 = pi25 & pi46;
  assign n8080 = ~n8078 ^ ~n8079;
  assign n8081 = pi24 & pi47;
  assign n8082 = ~n8080 ^ n8081;
  assign n8083 = ~n8077 ^ ~n8082;
  assign n8084 = ~n8072 ^ ~n8083;
  assign n8085 = ~n8065 ^ n8084;
  assign n8086 = pi32 & pi39;
  assign n8087 = pi31 & pi40;
  assign n8088 = ~n8086 ^ ~n8087;
  assign n8089 = pi30 & pi41;
  assign n8090 = ~n8088 ^ n8089;
  assign n8091 = pi29 & pi42;
  assign n8092 = pi28 & pi43;
  assign n8093 = ~n8091 ^ ~n8092;
  assign n8094 = pi27 & pi44;
  assign n8095 = ~n8093 ^ n8094;
  assign n8096 = ~n8090 ^ ~n8095;
  assign n8097 = pi23 & pi48;
  assign n8098 = pi18 & pi53;
  assign n8099 = ~n8097 ^ ~n8098;
  assign n8100 = pi17 & pi54;
  assign n8101 = ~n8099 ^ n8100;
  assign n8102 = ~n8096 ^ n8101;
  assign n8103 = ~n8085 ^ n8102;
  assign n8104 = n7989 & ~n8000;
  assign n8105 = n7985 & n7988;
  assign n8106 = ~n8104 & ~n8105;
  assign n8107 = n7882 & ~n7883;
  assign n8108 = ~n7880 & ~n7881;
  assign n8109 = ~n8107 & ~n8108;
  assign n8110 = pi11 & pi60;
  assign n8111 = pi10 & pi61;
  assign n8112 = ~n8110 ^ ~n8111;
  assign n8113 = pi08 & pi63;
  assign n8114 = ~n8112 ^ n8113;
  assign n8115 = ~n8109 ^ n8114;
  assign n8116 = n7870 & ~n7871;
  assign n8117 = ~n7868 & ~n7869;
  assign n8118 = ~n8116 & ~n8117;
  assign n8119 = ~n8115 ^ ~n8118;
  assign n8120 = pi21 & pi50;
  assign n8121 = pi20 & pi51;
  assign n8122 = ~n8120 ^ ~n8121;
  assign n8123 = pi19 & pi52;
  assign n8124 = ~n8122 ^ n8123;
  assign n8125 = pi35 & pi36;
  assign n8126 = pi34 & pi37;
  assign n8127 = ~n8125 ^ ~n8126;
  assign n8128 = pi33 & pi38;
  assign n8129 = ~n8127 ^ n8128;
  assign n8130 = ~n8124 ^ ~n8129;
  assign n8131 = pi09 & pi62;
  assign n8132 = pi22 & pi49;
  assign n8133 = ~n8131 ^ n8132;
  assign n8134 = ~n8133 ^ pi36;
  assign n8135 = ~n8130 ^ ~n8134;
  assign n8136 = ~n8119 ^ ~n8135;
  assign n8137 = ~n8106 ^ n8136;
  assign n8138 = ~n8103 ^ ~n8137;
  assign n8139 = ~n8062 ^ ~n8138;
  assign n8140 = n7898 & n7908;
  assign n8141 = ~n7902 & ~n7907;
  assign n8142 = ~n8140 & ~n8141;
  assign n8143 = n7888 & ~n7889;
  assign n8144 = ~n7886 & ~n7887;
  assign n8145 = ~n8143 & ~n8144;
  assign n8146 = n7877 & ~n7878;
  assign n8147 = ~n7875 & ~n7876;
  assign n8148 = ~n8146 & ~n8147;
  assign n8149 = ~n8145 ^ ~n8148;
  assign n8150 = n7912 & ~n7913;
  assign n8151 = ~n7910 & ~n7911;
  assign n8152 = ~n8150 & ~n8151;
  assign n8153 = ~n8149 ^ n8152;
  assign n8154 = ~n8142 ^ ~n8153;
  assign n8155 = n7923 & ~n7924;
  assign n8156 = ~n7921 & ~n7922;
  assign n8157 = ~n8155 & ~n8156;
  assign n8158 = n7905 & ~n7906;
  assign n8159 = ~n7903 & ~n7904;
  assign n8160 = ~n8158 & ~n8159;
  assign n8161 = ~n8157 ^ ~n8160;
  assign n8162 = n7900 & ~n7901;
  assign n8163 = ~n4009 & ~n7899;
  assign n8164 = ~n8162 & ~n8163;
  assign n8165 = ~n8161 ^ ~n8164;
  assign n8166 = ~n8154 ^ n8165;
  assign n8167 = n7996 & n7999;
  assign n8168 = n7992 & n7995;
  assign n8169 = ~n8167 & ~n8168;
  assign n8170 = n7920 & ~n7925;
  assign n8171 = ~n7914 & ~n7919;
  assign n8172 = ~n8170 & ~n8171;
  assign n8173 = ~n8169 ^ ~n8172;
  assign n8174 = n7885 & ~n7890;
  assign n8175 = ~n7879 & ~n7884;
  assign n8176 = ~n8174 & ~n8175;
  assign n8177 = ~n8173 ^ n8176;
  assign n8178 = ~n8166 ^ n8177;
  assign n8179 = ~n7928 & n7926;
  assign n8180 = n7895 & n7909;
  assign n8181 = ~n8179 & ~n8180;
  assign n8182 = ~n8178 ^ n8181;
  assign n8183 = ~n8139 ^ ~n8182;
  assign n8184 = ~n8058 ^ ~n8183;
  assign n8185 = ~n8054 ^ n8184;
  assign n8186 = ~n8021 ^ ~n8185;
  assign po072 = ~n8017 ^ ~n8186;
  assign n8188 = ~n8021 & n8025;
  assign n8189 = n8184 & ~n8053;
  assign n8190 = ~n8188 & ~n8189;
  assign n8191 = n8021 & ~n8025;
  assign n8192 = ~n8184 & n8053;
  assign n8193 = ~n8191 & ~n8192;
  assign n8194 = ~n8190 & n8193;
  assign n8195 = ~n8017 & n8194;
  assign n8196 = n8191 & n8192;
  assign n8197 = n8188 & n8189;
  assign n8198 = ~n8196 & ~n8197;
  assign n8199 = ~n8195 & n8198;
  assign n8200 = n8190 & ~n8193;
  assign n8201 = n8017 & n8200;
  assign n8202 = n8199 & ~n8201;
  assign n8203 = ~n8139 & ~n8182;
  assign n8204 = n8058 & ~n8203;
  assign n8205 = n8139 & n8182;
  assign n8206 = ~n8204 & ~n8205;
  assign n8207 = n8032 & n8051;
  assign n8208 = ~n8029 & ~n8207;
  assign n8209 = ~n8032 & ~n8051;
  assign n8210 = ~n8208 & ~n8209;
  assign n8211 = ~n8035 & n8050;
  assign n8212 = n8038 & n8049;
  assign n8213 = ~n8211 & ~n8212;
  assign n8214 = n8173 & ~n8176;
  assign n8215 = ~n8169 & ~n8172;
  assign n8216 = ~n8214 & ~n8215;
  assign n8217 = pi20 & pi52;
  assign n8218 = pi18 & pi54;
  assign n8219 = ~n8217 ^ ~n8218;
  assign n8220 = pi17 & pi55;
  assign n8221 = ~n8219 ^ n8220;
  assign n8222 = pi35 & pi37;
  assign n8223 = pi22 & pi50;
  assign n8224 = ~n8222 ^ ~n8223;
  assign n8225 = pi21 & pi51;
  assign n8226 = ~n8224 ^ n8225;
  assign n8227 = ~n8221 ^ ~n8226;
  assign n8228 = pi32 & pi40;
  assign n8229 = pi23 & pi49;
  assign n8230 = ~n8228 ^ ~n8229;
  assign n8231 = pi16 & pi56;
  assign n8232 = ~n8230 ^ n8231;
  assign n8233 = ~n8227 ^ n8232;
  assign n8234 = ~n8216 ^ n8233;
  assign n8235 = n8068 & n8071;
  assign n8236 = pi13 & pi59;
  assign n8237 = n7889 & n8236;
  assign n8238 = ~n8235 & ~n8237;
  assign n8239 = pi11 & pi61;
  assign n8240 = pi10 & pi62;
  assign n8241 = ~n8239 ^ ~n8240;
  assign n8242 = pi09 & pi63;
  assign n8243 = ~n8241 ^ n8242;
  assign n8244 = pi24 & pi48;
  assign n8245 = ~n4226 ^ ~n8244;
  assign n8246 = pi12 & pi60;
  assign n8247 = ~n8245 ^ n8246;
  assign n8248 = ~n8243 ^ ~n8247;
  assign n8249 = ~n8238 ^ n8248;
  assign n8250 = ~n8234 ^ ~n8249;
  assign n8251 = n8045 & ~n8048;
  assign n8252 = ~n8041 & n8044;
  assign n8253 = ~n8251 & ~n8252;
  assign n8254 = n8112 & ~n8113;
  assign n8255 = ~n8110 & ~n8111;
  assign n8256 = ~n8254 & ~n8255;
  assign n8257 = n8080 & ~n8081;
  assign n8258 = ~n8078 & ~n8079;
  assign n8259 = ~n8257 & ~n8258;
  assign n8260 = ~n8256 ^ ~n8259;
  assign n8261 = n8075 & ~n8076;
  assign n8262 = ~n8073 & ~n8074;
  assign n8263 = ~n8261 & ~n8262;
  assign n8264 = ~n8260 ^ n8263;
  assign n8265 = ~n8253 ^ ~n8264;
  assign n8266 = pi34 & pi38;
  assign n8267 = pi33 & pi39;
  assign n8268 = ~n8266 ^ ~n8267;
  assign n8269 = pi19 & pi53;
  assign n8270 = ~n8268 ^ n8269;
  assign n8271 = pi15 & pi57;
  assign n8272 = pi14 & pi58;
  assign n8273 = ~n8271 ^ ~n8272;
  assign n8274 = ~n8273 ^ n8236;
  assign n8275 = ~n8270 ^ ~n8274;
  assign n8276 = pi28 & pi44;
  assign n8277 = pi27 & pi45;
  assign n8278 = ~n8276 ^ ~n8277;
  assign n8279 = pi26 & pi46;
  assign n8280 = ~n8278 ^ n8279;
  assign n8281 = ~n8275 ^ n8280;
  assign n8282 = ~n8265 ^ ~n8281;
  assign n8283 = ~n8250 ^ ~n8282;
  assign n8284 = ~n8213 ^ ~n8283;
  assign n8285 = n8085 & ~n8102;
  assign n8286 = n8065 & ~n8084;
  assign n8287 = ~n8285 & ~n8286;
  assign n8288 = n8072 & n8083;
  assign n8289 = ~n8077 & ~n8082;
  assign n8290 = ~n8288 & ~n8289;
  assign n8291 = n8122 & ~n8123;
  assign n8292 = ~n8120 & ~n8121;
  assign n8293 = ~n8291 & ~n8292;
  assign n8294 = n8127 & ~n8128;
  assign n8295 = ~n8125 & ~n8126;
  assign n8296 = ~n8294 & ~n8295;
  assign n8297 = ~n8293 ^ ~n8296;
  assign n8298 = n5535 & pi49;
  assign n8299 = ~n8298 & ~n8131;
  assign n8300 = ~n8132 & ~pi36;
  assign n8301 = ~n8299 & ~n8300;
  assign n8302 = ~n8297 ^ ~n8301;
  assign n8303 = ~n8290 ^ n8302;
  assign n8304 = n8093 & ~n8094;
  assign n8305 = ~n8091 & ~n8092;
  assign n8306 = ~n8304 & ~n8305;
  assign n8307 = n8099 & ~n8100;
  assign n8308 = ~n8097 & ~n8098;
  assign n8309 = ~n8307 & ~n8308;
  assign n8310 = ~n8306 ^ ~n8309;
  assign n8311 = n8088 & ~n8089;
  assign n8312 = ~n8086 & ~n8087;
  assign n8313 = ~n8311 & ~n8312;
  assign n8314 = ~n8310 ^ ~n8313;
  assign n8315 = ~n8303 ^ ~n8314;
  assign n8316 = n8149 & ~n8152;
  assign n8317 = ~n8145 & ~n8148;
  assign n8318 = ~n8316 & ~n8317;
  assign n8319 = n8130 & n8134;
  assign n8320 = ~n8124 & ~n8129;
  assign n8321 = ~n8319 & ~n8320;
  assign n8322 = n8096 & ~n8101;
  assign n8323 = ~n8090 & ~n8095;
  assign n8324 = ~n8322 & ~n8323;
  assign n8325 = ~n8321 ^ ~n8324;
  assign n8326 = ~n8318 ^ ~n8325;
  assign n8327 = ~n8315 ^ ~n8326;
  assign n8328 = ~n8287 ^ n8327;
  assign n8329 = ~n8284 ^ ~n8328;
  assign n8330 = ~n8210 ^ ~n8329;
  assign n8331 = ~n8103 & ~n8137;
  assign n8332 = ~n8062 & ~n8331;
  assign n8333 = n8103 & n8137;
  assign n8334 = ~n8332 & ~n8333;
  assign n8335 = n8178 & ~n8181;
  assign n8336 = ~n8166 & n8177;
  assign n8337 = ~n8335 & ~n8336;
  assign n8338 = n8154 & ~n8165;
  assign n8339 = n8142 & n8153;
  assign n8340 = ~n8338 & ~n8339;
  assign n8341 = n8161 & n8164;
  assign n8342 = n8157 & n8160;
  assign n8343 = ~n8341 & ~n8342;
  assign n8344 = pi31 & pi41;
  assign n8345 = pi30 & pi42;
  assign n8346 = ~n8344 ^ ~n8345;
  assign n8347 = pi29 & pi43;
  assign n8348 = ~n8346 ^ n8347;
  assign n8349 = ~n8343 ^ ~n8348;
  assign n8350 = n8115 & n8118;
  assign n8351 = n8109 & ~n8114;
  assign n8352 = ~n8350 & ~n8351;
  assign n8353 = ~n8349 ^ n8352;
  assign n8354 = ~n8340 ^ ~n8353;
  assign n8355 = ~n8106 & n8136;
  assign n8356 = ~n8119 & ~n8135;
  assign n8357 = ~n8355 & ~n8356;
  assign n8358 = ~n8354 ^ ~n8357;
  assign n8359 = ~n8337 ^ n8358;
  assign n8360 = ~n8334 ^ ~n8359;
  assign n8361 = ~n8330 ^ ~n8360;
  assign n8362 = ~n8206 ^ ~n8361;
  assign po073 = ~n8202 ^ n8362;
  assign n8364 = ~n8191 & ~n8362;
  assign n8365 = ~n8364 & ~n8189;
  assign n8366 = ~n8362 & ~n8192;
  assign n8367 = ~n8188 & ~n8366;
  assign n8368 = ~n8365 & ~n8367;
  assign n8369 = n8017 & ~n8368;
  assign n8370 = ~n8196 & ~n8362;
  assign n8371 = ~n8194 & ~n8370;
  assign n8372 = ~n8369 & ~n8371;
  assign n8373 = n8330 & n8360;
  assign n8374 = n8206 & ~n8373;
  assign n8375 = ~n8330 & ~n8360;
  assign n8376 = ~n8374 & ~n8375;
  assign n8377 = n8284 & n8328;
  assign n8378 = n8210 & ~n8377;
  assign n8379 = ~n8284 & ~n8328;
  assign n8380 = ~n8378 & ~n8379;
  assign n8381 = n8213 & n8283;
  assign n8382 = ~n8250 & ~n8282;
  assign n8383 = ~n8381 & ~n8382;
  assign n8384 = ~n8328 & ~n8315;
  assign n8385 = ~n8287 & ~n8326;
  assign n8386 = ~n8384 & ~n8385;
  assign n8387 = n8265 & n8281;
  assign n8388 = ~n8253 & ~n8264;
  assign n8389 = ~n8387 & ~n8388;
  assign n8390 = n8260 & ~n8263;
  assign n8391 = ~n8256 & ~n8259;
  assign n8392 = ~n8390 & ~n8391;
  assign n8393 = pi33 & pi40;
  assign n8394 = pi32 & pi41;
  assign n8395 = ~n8393 ^ ~n8394;
  assign n8396 = pi31 & pi42;
  assign n8397 = ~n8395 ^ n8396;
  assign n8398 = ~n8392 ^ n8397;
  assign n8399 = n8310 & n8313;
  assign n8400 = n8306 & n8309;
  assign n8401 = ~n8399 & ~n8400;
  assign n8402 = ~n8398 ^ n8401;
  assign n8403 = ~n8389 ^ n8402;
  assign n8404 = n8303 & n8314;
  assign n8405 = ~n8290 & n8302;
  assign n8406 = ~n8404 & ~n8405;
  assign n8407 = ~n8403 ^ n8406;
  assign n8408 = ~n8386 ^ ~n8407;
  assign n8409 = ~n8383 ^ n8408;
  assign n8410 = ~n8380 ^ ~n8409;
  assign n8411 = ~n8337 & n8358;
  assign n8412 = ~n8334 & ~n8411;
  assign n8413 = n8337 & ~n8358;
  assign n8414 = ~n8412 & ~n8413;
  assign n8415 = n8354 & n8357;
  assign n8416 = n8340 & n8353;
  assign n8417 = ~n8415 & ~n8416;
  assign n8418 = n8349 & ~n8352;
  assign n8419 = ~n8343 & ~n8348;
  assign n8420 = ~n8418 & ~n8419;
  assign n8421 = pi30 & pi43;
  assign n8422 = pi29 & pi44;
  assign n8423 = ~n8421 ^ ~n8422;
  assign n8424 = pi28 & pi45;
  assign n8425 = ~n8423 ^ n8424;
  assign n8426 = pi12 & pi61;
  assign n8427 = ~n4229 ^ ~n8426;
  assign n8428 = pi10 & pi63;
  assign n8429 = ~n8427 ^ n8428;
  assign n8430 = ~n8425 ^ ~n8429;
  assign n8431 = pi36 & pi37;
  assign n8432 = pi35 & pi38;
  assign n8433 = ~n8431 ^ ~n8432;
  assign n8434 = pi34 & pi39;
  assign n8435 = ~n8433 ^ n8434;
  assign n8436 = ~n8430 ^ ~n8435;
  assign n8437 = ~n8420 ^ ~n8436;
  assign n8438 = n8346 & ~n8347;
  assign n8439 = ~n8344 & ~n8345;
  assign n8440 = ~n8438 & ~n8439;
  assign n8441 = n8273 & ~n8236;
  assign n8442 = ~n8271 & ~n8272;
  assign n8443 = ~n8441 & ~n8442;
  assign n8444 = ~n8440 ^ ~n8443;
  assign n8445 = n8278 & ~n8279;
  assign n8446 = ~n8276 & ~n8277;
  assign n8447 = ~n8445 & ~n8446;
  assign n8448 = ~n8444 ^ ~n8447;
  assign n8449 = ~n8437 ^ n8448;
  assign n8450 = n8318 & n8325;
  assign n8451 = ~n8321 & ~n8324;
  assign n8452 = ~n8450 & ~n8451;
  assign n8453 = pi22 & pi51;
  assign n8454 = pi21 & pi52;
  assign n8455 = ~n8453 ^ ~n8454;
  assign n8456 = pi20 & pi53;
  assign n8457 = ~n8455 ^ n8456;
  assign n8458 = pi19 & pi54;
  assign n8459 = ~n4315 ^ ~n8458;
  assign n8460 = pi18 & pi55;
  assign n8461 = ~n8459 ^ n8460;
  assign n8462 = ~n8457 ^ ~n8461;
  assign n8463 = pi11 & pi62;
  assign n8464 = pi23 & pi50;
  assign n8465 = ~n8463 ^ n8464;
  assign n8466 = ~n8465 ^ pi37;
  assign n8467 = ~n8462 ^ n8466;
  assign n8468 = ~n8452 ^ ~n8467;
  assign n8469 = n8230 & ~n8231;
  assign n8470 = ~n8228 & ~n8229;
  assign n8471 = ~n8469 & ~n8470;
  assign n8472 = pi27 & pi46;
  assign n8473 = pi26 & pi47;
  assign n8474 = ~n8472 ^ ~n8473;
  assign n8475 = pi17 & pi56;
  assign n8476 = ~n8474 ^ n8475;
  assign n8477 = ~n8471 ^ n8476;
  assign n8478 = pi16 & pi57;
  assign n8479 = pi15 & pi58;
  assign n8480 = ~n8478 ^ ~n8479;
  assign n8481 = pi14 & pi59;
  assign n8482 = ~n8480 ^ n8481;
  assign n8483 = ~n8477 ^ n8482;
  assign n8484 = ~n8468 ^ ~n8483;
  assign n8485 = ~n8449 ^ n8484;
  assign n8486 = ~n8417 ^ n8485;
  assign n8487 = n8234 & n8249;
  assign n8488 = ~n8216 & n8233;
  assign n8489 = ~n8487 & ~n8488;
  assign n8490 = n8224 & ~n8225;
  assign n8491 = ~n8222 & ~n8223;
  assign n8492 = ~n8490 & ~n8491;
  assign n8493 = pi13 & pi60;
  assign n8494 = ~n8492 ^ ~n8493;
  assign n8495 = n8268 & ~n8269;
  assign n8496 = ~n8266 & ~n8267;
  assign n8497 = ~n8495 & ~n8496;
  assign n8498 = ~n8494 ^ ~n8497;
  assign n8499 = n8227 & ~n8232;
  assign n8500 = ~n8221 & ~n8226;
  assign n8501 = ~n8499 & ~n8500;
  assign n8502 = ~n8498 ^ n8501;
  assign n8503 = n8219 & ~n8220;
  assign n8504 = ~n8217 & ~n8218;
  assign n8505 = ~n8503 & ~n8504;
  assign n8506 = n8241 & ~n8242;
  assign n8507 = ~n8239 & ~n8240;
  assign n8508 = ~n8506 & ~n8507;
  assign n8509 = ~n8505 ^ ~n8508;
  assign n8510 = n8245 & ~n8246;
  assign n8511 = ~n4226 & ~n8244;
  assign n8512 = ~n8510 & ~n8511;
  assign n8513 = ~n8509 ^ n8512;
  assign n8514 = ~n8502 ^ ~n8513;
  assign n8515 = ~n8489 ^ ~n8514;
  assign n8516 = ~n8238 & n8248;
  assign n8517 = ~n8243 & ~n8247;
  assign n8518 = ~n8516 & ~n8517;
  assign n8519 = n8297 & n8301;
  assign n8520 = n8293 & n8296;
  assign n8521 = ~n8519 & ~n8520;
  assign n8522 = ~n8518 ^ ~n8521;
  assign n8523 = n8275 & ~n8280;
  assign n8524 = ~n8270 & ~n8274;
  assign n8525 = ~n8523 & ~n8524;
  assign n8526 = ~n8522 ^ n8525;
  assign n8527 = ~n8515 ^ ~n8526;
  assign n8528 = ~n8486 ^ ~n8527;
  assign n8529 = ~n8414 ^ ~n8528;
  assign n8530 = ~n8410 ^ ~n8529;
  assign n8531 = ~n8376 ^ ~n8530;
  assign po074 = n8372 ^ n8531;
  assign n8533 = ~n8376 & ~n8529;
  assign n8534 = n8372 & ~n8533;
  assign n8535 = n8376 & n8529;
  assign n8536 = ~n8380 & ~n8409;
  assign n8537 = ~n8535 & ~n8536;
  assign n8538 = n8380 & n8409;
  assign n8539 = ~n8537 & ~n8538;
  assign n8540 = n8534 & n8539;
  assign n8541 = ~n8533 & ~n8538;
  assign n8542 = n8537 & ~n8541;
  assign n8543 = ~n8372 & n8542;
  assign n8544 = n8535 & n8536;
  assign n8545 = n8533 & n8538;
  assign n8546 = ~n8544 & ~n8545;
  assign n8547 = ~n8543 & n8546;
  assign n8548 = ~n8540 & n8547;
  assign n8549 = ~n8383 & n8408;
  assign n8550 = ~n8386 & ~n8407;
  assign n8551 = ~n8549 & ~n8550;
  assign n8552 = n8437 & ~n8448;
  assign n8553 = n8420 & n8436;
  assign n8554 = ~n8552 & ~n8553;
  assign n8555 = n8468 & n8483;
  assign n8556 = ~n8452 & ~n8467;
  assign n8557 = ~n8555 & ~n8556;
  assign n8558 = ~n8554 ^ n8557;
  assign n8559 = n8398 & ~n8401;
  assign n8560 = n8392 & ~n8397;
  assign n8561 = ~n8559 & ~n8560;
  assign n8562 = n8433 & ~n8434;
  assign n8563 = ~n8431 & ~n8432;
  assign n8564 = ~n8562 & ~n8563;
  assign n8565 = pi16 & pi58;
  assign n8566 = pi15 & pi59;
  assign n8567 = ~n8565 ^ ~n8566;
  assign n8568 = pi14 & pi60;
  assign n8569 = ~n8567 ^ n8568;
  assign n8570 = ~n8564 ^ n8569;
  assign n8571 = n8395 & ~n8396;
  assign n8572 = ~n8393 & ~n8394;
  assign n8573 = ~n8571 & ~n8572;
  assign n8574 = ~n8570 ^ n8573;
  assign n8575 = ~n8561 ^ ~n8574;
  assign n8576 = n8462 & ~n8466;
  assign n8577 = n8457 & n8461;
  assign n8578 = ~n8576 & ~n8577;
  assign n8579 = ~n8575 ^ n8578;
  assign n8580 = ~n8558 ^ n8579;
  assign n8581 = ~n8551 ^ ~n8580;
  assign n8582 = n8403 & ~n8406;
  assign n8583 = ~n8389 & n8402;
  assign n8584 = ~n8582 & ~n8583;
  assign n8585 = n8444 & n8447;
  assign n8586 = n8440 & n8443;
  assign n8587 = ~n8585 & ~n8586;
  assign n8588 = n5956 & pi50;
  assign n8589 = ~n8588 & ~n8463;
  assign n8590 = ~n8464 & ~pi37;
  assign n8591 = ~n8589 & ~n8590;
  assign n8592 = pi12 & pi62;
  assign n8593 = pi13 & pi61;
  assign n8594 = ~n8592 ^ ~n8593;
  assign n8595 = ~n8591 ^ ~n8594;
  assign n8596 = pi30 & pi44;
  assign n8597 = pi29 & pi45;
  assign n8598 = ~n8596 ^ ~n8597;
  assign n8599 = pi17 & pi57;
  assign n8600 = ~n8598 ^ n8599;
  assign n8601 = ~n8595 ^ n8600;
  assign n8602 = ~n8587 ^ n8601;
  assign n8603 = pi33 & pi41;
  assign n8604 = pi25 & pi49;
  assign n8605 = ~n8603 ^ ~n8604;
  assign n8606 = pi18 & pi56;
  assign n8607 = ~n8605 ^ n8606;
  assign n8608 = pi32 & pi42;
  assign n8609 = pi31 & pi43;
  assign n8610 = ~n8608 ^ ~n8609;
  assign n8611 = pi11 & pi63;
  assign n8612 = ~n8610 ^ n8611;
  assign n8613 = ~n8607 ^ ~n8612;
  assign n8614 = pi28 & pi46;
  assign n8615 = pi27 & pi47;
  assign n8616 = ~n8614 ^ ~n8615;
  assign n8617 = pi26 & pi48;
  assign n8618 = ~n8616 ^ n8617;
  assign n8619 = ~n8613 ^ n8618;
  assign n8620 = pi22 & pi52;
  assign n8621 = pi21 & pi53;
  assign n8622 = ~n8620 ^ ~n8621;
  assign n8623 = pi19 & pi55;
  assign n8624 = ~n8622 ^ n8623;
  assign n8625 = pi35 & pi39;
  assign n8626 = pi34 & pi40;
  assign n8627 = ~n8625 ^ ~n8626;
  assign n8628 = pi20 & pi54;
  assign n8629 = ~n8627 ^ n8628;
  assign n8630 = ~n8624 ^ ~n8629;
  assign n8631 = pi36 & pi38;
  assign n8632 = pi24 & pi50;
  assign n8633 = ~n8631 ^ ~n8632;
  assign n8634 = pi23 & pi51;
  assign n8635 = ~n8633 ^ n8634;
  assign n8636 = ~n8630 ^ n8635;
  assign n8637 = ~n8619 ^ ~n8636;
  assign n8638 = ~n8602 ^ n8637;
  assign n8639 = n8423 & ~n8424;
  assign n8640 = ~n8421 & ~n8422;
  assign n8641 = ~n8639 & ~n8640;
  assign n8642 = n8474 & ~n8475;
  assign n8643 = ~n8472 & ~n8473;
  assign n8644 = ~n8642 & ~n8643;
  assign n8645 = ~n8641 ^ ~n8644;
  assign n8646 = n8480 & ~n8481;
  assign n8647 = ~n8478 & ~n8479;
  assign n8648 = ~n8646 & ~n8647;
  assign n8649 = ~n8645 ^ ~n8648;
  assign n8650 = n8430 & n8435;
  assign n8651 = n8425 & n8429;
  assign n8652 = ~n8650 & ~n8651;
  assign n8653 = ~n8649 ^ ~n8652;
  assign n8654 = n8455 & ~n8456;
  assign n8655 = ~n8453 & ~n8454;
  assign n8656 = ~n8654 & ~n8655;
  assign n8657 = n8459 & ~n8460;
  assign n8658 = ~n4315 & ~n8458;
  assign n8659 = ~n8657 & ~n8658;
  assign n8660 = ~n8656 ^ ~n8659;
  assign n8661 = n8427 & ~n8428;
  assign n8662 = ~n4229 & ~n8426;
  assign n8663 = ~n8661 & ~n8662;
  assign n8664 = ~n8660 ^ ~n8663;
  assign n8665 = ~n8653 ^ n8664;
  assign n8666 = ~n8638 ^ ~n8665;
  assign n8667 = ~n8584 ^ n8666;
  assign n8668 = ~n8581 ^ n8667;
  assign n8669 = n8515 & n8526;
  assign n8670 = ~n8489 & ~n8514;
  assign n8671 = ~n8669 & ~n8670;
  assign n8672 = n8522 & ~n8525;
  assign n8673 = ~n8518 & ~n8521;
  assign n8674 = ~n8672 & ~n8673;
  assign n8675 = n8477 & ~n8482;
  assign n8676 = n8471 & ~n8476;
  assign n8677 = ~n8675 & ~n8676;
  assign n8678 = n8494 & n8497;
  assign n8679 = n8492 & n8493;
  assign n8680 = ~n8678 & ~n8679;
  assign n8681 = ~n8677 ^ ~n8680;
  assign n8682 = n8509 & ~n8512;
  assign n8683 = ~n8505 & ~n8508;
  assign n8684 = ~n8682 & ~n8683;
  assign n8685 = ~n8681 ^ n8684;
  assign n8686 = ~n8674 ^ ~n8685;
  assign n8687 = n8502 & n8513;
  assign n8688 = ~n8498 & n8501;
  assign n8689 = ~n8687 & ~n8688;
  assign n8690 = ~n8686 ^ ~n8689;
  assign n8691 = ~n8671 ^ n8690;
  assign n8692 = n8449 & ~n8484;
  assign n8693 = ~n8417 & ~n8692;
  assign n8694 = ~n8449 & n8484;
  assign n8695 = ~n8693 & ~n8694;
  assign n8696 = ~n8691 ^ n8695;
  assign n8697 = ~n8668 ^ n8696;
  assign n8698 = n8414 & n8528;
  assign n8699 = n8486 & n8527;
  assign n8700 = ~n8698 & ~n8699;
  assign n8701 = ~n8697 ^ ~n8700;
  assign po075 = ~n8548 ^ n8701;
  assign n8703 = ~n8701 & ~n8538;
  assign n8704 = ~n8703 & ~n8535;
  assign n8705 = ~n8534 & n8704;
  assign n8706 = ~n8533 & ~n8701;
  assign n8707 = ~n8706 & ~n8536;
  assign n8708 = ~n8372 & n8707;
  assign n8709 = ~n8539 & n8701;
  assign n8710 = ~n8708 & ~n8709;
  assign n8711 = ~n8705 & n8710;
  assign n8712 = ~n8668 & n8696;
  assign n8713 = ~n8712 & n8700;
  assign n8714 = n8668 & ~n8696;
  assign n8715 = ~n8713 & ~n8714;
  assign n8716 = n8581 & ~n8667;
  assign n8717 = ~n8551 & ~n8580;
  assign n8718 = ~n8716 & ~n8717;
  assign n8719 = ~n8584 & n8666;
  assign n8720 = ~n8638 & ~n8665;
  assign n8721 = ~n8719 & ~n8720;
  assign n8722 = n8575 & ~n8578;
  assign n8723 = n8561 & n8574;
  assign n8724 = ~n8722 & ~n8723;
  assign n8725 = n8653 & ~n8664;
  assign n8726 = ~n8649 & ~n8652;
  assign n8727 = ~n8725 & ~n8726;
  assign n8728 = ~n8724 ^ ~n8727;
  assign n8729 = pi33 & pi42;
  assign n8730 = pi32 & pi43;
  assign n8731 = ~n8729 ^ ~n8730;
  assign n8732 = pi31 & pi44;
  assign n8733 = ~n8731 ^ n8732;
  assign n8734 = pi24 & pi51;
  assign n8735 = pi22 & pi53;
  assign n8736 = ~n8734 ^ ~n8735;
  assign n8737 = pi21 & pi54;
  assign n8738 = ~n8736 ^ n8737;
  assign n8739 = ~n8733 ^ ~n8738;
  assign n8740 = pi34 & pi41;
  assign n8741 = pi25 & pi50;
  assign n8742 = ~n8740 ^ ~n8741;
  assign n8743 = pi20 & pi55;
  assign n8744 = ~n8742 ^ n8743;
  assign n8745 = ~n8739 ^ n8744;
  assign n8746 = ~n8728 ^ n8745;
  assign n8747 = ~n8721 ^ ~n8746;
  assign n8748 = n8558 & ~n8579;
  assign n8749 = n8554 & ~n8557;
  assign n8750 = ~n8748 & ~n8749;
  assign n8751 = ~n8747 ^ n8750;
  assign n8752 = n8691 & ~n8695;
  assign n8753 = ~n8671 & n8690;
  assign n8754 = ~n8752 & ~n8753;
  assign n8755 = n8686 & n8689;
  assign n8756 = ~n8674 & ~n8685;
  assign n8757 = ~n8755 & ~n8756;
  assign n8758 = n8613 & ~n8618;
  assign n8759 = ~n8607 & ~n8612;
  assign n8760 = ~n8758 & ~n8759;
  assign n8761 = n8598 & ~n8599;
  assign n8762 = ~n8596 & ~n8597;
  assign n8763 = ~n8761 & ~n8762;
  assign n8764 = n8616 & ~n8617;
  assign n8765 = ~n8614 & ~n8615;
  assign n8766 = ~n8764 & ~n8765;
  assign n8767 = ~n8763 ^ ~n8766;
  assign n8768 = n8567 & ~n8568;
  assign n8769 = ~n8565 & ~n8566;
  assign n8770 = ~n8768 & ~n8769;
  assign n8771 = ~n8767 ^ n8770;
  assign n8772 = ~n8760 ^ ~n8771;
  assign n8773 = n8630 & ~n8635;
  assign n8774 = ~n8624 & ~n8629;
  assign n8775 = ~n8773 & ~n8774;
  assign n8776 = ~n8772 ^ n8775;
  assign n8777 = ~n8757 ^ n8776;
  assign n8778 = n8681 & ~n8684;
  assign n8779 = n8677 & n8680;
  assign n8780 = ~n8778 & ~n8779;
  assign n8781 = pi16 & pi59;
  assign n8782 = pi15 & pi60;
  assign n8783 = ~n8781 ^ ~n8782;
  assign n8784 = pi14 & pi61;
  assign n8785 = ~n8783 ^ n8784;
  assign n8786 = pi26 & pi49;
  assign n8787 = pi18 & pi57;
  assign n8788 = ~n8786 ^ ~n8787;
  assign n8789 = pi17 & pi58;
  assign n8790 = ~n8788 ^ n8789;
  assign n8791 = ~n8785 ^ ~n8790;
  assign n8792 = pi29 & pi46;
  assign n8793 = pi28 & pi47;
  assign n8794 = ~n8792 ^ ~n8793;
  assign n8795 = pi27 & pi48;
  assign n8796 = ~n8794 ^ n8795;
  assign n8797 = ~n8791 ^ n8796;
  assign n8798 = pi36 & pi39;
  assign n8799 = pi35 & pi40;
  assign n8800 = ~n8798 ^ ~n8799;
  assign n8801 = pi23 & pi52;
  assign n8802 = ~n8800 ^ n8801;
  assign n8803 = pi30 & pi45;
  assign n8804 = pi19 & pi56;
  assign n8805 = ~n8803 ^ ~n8804;
  assign n8806 = pi12 & pi63;
  assign n8807 = ~n8805 ^ n8806;
  assign n8808 = ~n8802 ^ ~n8807;
  assign n8809 = pi13 & pi62;
  assign n8810 = ~pi37 & pi38;
  assign n8811 = ~n8809 ^ ~n8810;
  assign n8812 = ~n8808 ^ ~n8811;
  assign n8813 = ~n8797 ^ ~n8812;
  assign n8814 = ~n8780 ^ ~n8813;
  assign n8815 = ~n8777 ^ n8814;
  assign n8816 = ~n8587 & n8601;
  assign n8817 = n8595 & ~n8600;
  assign n8818 = ~n8816 & ~n8817;
  assign n8819 = n8591 & n8594;
  assign n8820 = pi61 & pi62;
  assign n8821 = n1188 & n8820;
  assign n8822 = ~n8819 & ~n8821;
  assign n8823 = n8605 & ~n8606;
  assign n8824 = ~n8603 & ~n8604;
  assign n8825 = ~n8823 & ~n8824;
  assign n8826 = n8610 & ~n8611;
  assign n8827 = ~n8608 & ~n8609;
  assign n8828 = ~n8826 & ~n8827;
  assign n8829 = ~n8825 ^ ~n8828;
  assign n8830 = ~n8822 ^ ~n8829;
  assign n8831 = n8633 & ~n8634;
  assign n8832 = ~n8631 & ~n8632;
  assign n8833 = ~n8831 & ~n8832;
  assign n8834 = n8622 & ~n8623;
  assign n8835 = ~n8620 & ~n8621;
  assign n8836 = ~n8834 & ~n8835;
  assign n8837 = ~n8833 ^ ~n8836;
  assign n8838 = n8627 & ~n8628;
  assign n8839 = ~n8625 & ~n8626;
  assign n8840 = ~n8838 & ~n8839;
  assign n8841 = ~n8837 ^ ~n8840;
  assign n8842 = ~n8830 ^ n8841;
  assign n8843 = ~n8818 ^ n8842;
  assign n8844 = n8660 & n8663;
  assign n8845 = n8656 & n8659;
  assign n8846 = ~n8844 & ~n8845;
  assign n8847 = n8645 & n8648;
  assign n8848 = n8641 & n8644;
  assign n8849 = ~n8847 & ~n8848;
  assign n8850 = ~n8846 ^ ~n8849;
  assign n8851 = n8570 & ~n8573;
  assign n8852 = ~n8564 & n8569;
  assign n8853 = ~n8851 & ~n8852;
  assign n8854 = ~n8850 ^ n8853;
  assign n8855 = ~n8843 ^ n8854;
  assign n8856 = ~n8602 & n8637;
  assign n8857 = ~n8619 & ~n8636;
  assign n8858 = ~n8856 & ~n8857;
  assign n8859 = ~n8855 ^ n8858;
  assign n8860 = ~n8815 ^ ~n8859;
  assign n8861 = ~n8754 ^ n8860;
  assign n8862 = ~n8751 ^ ~n8861;
  assign n8863 = ~n8718 ^ n8862;
  assign n8864 = ~n8715 ^ n8863;
  assign po076 = ~n8711 ^ ~n8864;
  assign n8866 = n8715 & n8718;
  assign n8867 = n8751 & n8861;
  assign n8868 = ~n8866 & ~n8867;
  assign n8869 = ~n8751 & ~n8861;
  assign n8870 = ~n8868 & ~n8869;
  assign n8871 = ~n8715 & ~n8718;
  assign n8872 = n8870 & ~n8871;
  assign n8873 = n8711 & ~n8872;
  assign n8874 = ~n8871 & ~n8869;
  assign n8875 = n8868 & ~n8874;
  assign n8876 = ~n8711 & ~n8875;
  assign n8877 = ~n8873 & ~n8876;
  assign n8878 = n8871 & n8869;
  assign n8879 = n8866 & n8867;
  assign n8880 = ~n8878 & ~n8879;
  assign n8881 = ~n8877 & n8880;
  assign n8882 = ~n8754 & n8860;
  assign n8883 = ~n8815 & ~n8859;
  assign n8884 = ~n8882 & ~n8883;
  assign n8885 = n8777 & ~n8814;
  assign n8886 = n8757 & ~n8776;
  assign n8887 = ~n8885 & ~n8886;
  assign n8888 = ~n8843 & n8841;
  assign n8889 = ~n8818 & ~n8830;
  assign n8890 = ~n8888 & ~n8889;
  assign n8891 = n8772 & ~n8775;
  assign n8892 = ~n8760 & ~n8771;
  assign n8893 = ~n8891 & ~n8892;
  assign n8894 = ~n8890 ^ ~n8893;
  assign n8895 = pi32 & pi44;
  assign n8896 = pi31 & pi45;
  assign n8897 = ~n8895 ^ ~n8896;
  assign n8898 = pi13 & pi63;
  assign n8899 = ~n8897 ^ n8898;
  assign n8900 = pi33 & pi43;
  assign n8901 = pi23 & pi53;
  assign n8902 = ~n8900 ^ ~n8901;
  assign n8903 = pi19 & pi57;
  assign n8904 = ~n8902 ^ n8903;
  assign n8905 = ~n8899 ^ ~n8904;
  assign n8906 = pi22 & pi54;
  assign n8907 = pi21 & pi55;
  assign n8908 = ~n8906 ^ ~n8907;
  assign n8909 = pi20 & pi56;
  assign n8910 = ~n8908 ^ n8909;
  assign n8911 = ~n8905 ^ n8910;
  assign n8912 = ~n8894 ^ ~n8911;
  assign n8913 = ~n8887 ^ ~n8912;
  assign n8914 = n8855 & ~n8858;
  assign n8915 = ~n8843 & n8854;
  assign n8916 = ~n8914 & ~n8915;
  assign n8917 = ~n8913 ^ n8916;
  assign n8918 = ~n8884 ^ ~n8917;
  assign n8919 = n8747 & ~n8750;
  assign n8920 = ~n8721 & ~n8746;
  assign n8921 = ~n8919 & ~n8920;
  assign n8922 = n8728 & ~n8745;
  assign n8923 = ~n8724 & ~n8727;
  assign n8924 = ~n8922 & ~n8923;
  assign n8925 = n8808 & n8811;
  assign n8926 = ~n8802 & ~n8807;
  assign n8927 = ~n8925 & ~n8926;
  assign n8928 = n8791 & ~n8796;
  assign n8929 = ~n8785 & ~n8790;
  assign n8930 = ~n8928 & ~n8929;
  assign n8931 = ~n8927 ^ ~n8930;
  assign n8932 = n8731 & ~n8732;
  assign n8933 = ~n8729 & ~n8730;
  assign n8934 = ~n8932 & ~n8933;
  assign n8935 = n8788 & ~n8789;
  assign n8936 = ~n8786 & ~n8787;
  assign n8937 = ~n8935 & ~n8936;
  assign n8938 = ~n8934 ^ ~n8937;
  assign n8939 = n8783 & ~n8784;
  assign n8940 = ~n8781 & ~n8782;
  assign n8941 = ~n8939 & ~n8940;
  assign n8942 = ~n8938 ^ ~n8941;
  assign n8943 = ~n8931 ^ n8942;
  assign n8944 = ~n8924 ^ n8943;
  assign n8945 = n8850 & ~n8853;
  assign n8946 = n8846 & n8849;
  assign n8947 = ~n8945 & ~n8946;
  assign n8948 = pi36 & pi40;
  assign n8949 = pi35 & pi41;
  assign n8950 = ~n8948 ^ ~n8949;
  assign n8951 = pi34 & pi42;
  assign n8952 = ~n8950 ^ n8951;
  assign n8953 = pi37 & pi39;
  assign n8954 = pi25 & pi51;
  assign n8955 = ~n8953 ^ ~n8954;
  assign n8956 = pi24 & pi52;
  assign n8957 = ~n8955 ^ n8956;
  assign n8958 = ~n8952 ^ ~n8957;
  assign n8959 = pi30 & pi46;
  assign n8960 = pi29 & pi47;
  assign n8961 = ~n8959 ^ ~n8960;
  assign n8962 = pi28 & pi48;
  assign n8963 = ~n8961 ^ n8962;
  assign n8964 = ~n8958 ^ ~n8963;
  assign n8965 = ~n8947 ^ n8964;
  assign n8966 = n8736 & ~n8737;
  assign n8967 = ~n8734 & ~n8735;
  assign n8968 = ~n8966 & ~n8967;
  assign n8969 = pi27 & pi49;
  assign n8970 = ~n4492 ^ ~n8969;
  assign n8971 = pi18 & pi58;
  assign n8972 = ~n8970 ^ n8971;
  assign n8973 = ~n8968 ^ n8972;
  assign n8974 = pi17 & pi59;
  assign n8975 = pi16 & pi60;
  assign n8976 = ~n8974 ^ ~n8975;
  assign n8977 = pi15 & pi61;
  assign n8978 = ~n8976 ^ n8977;
  assign n8979 = ~n8973 ^ ~n8978;
  assign n8980 = ~n8965 ^ n8979;
  assign n8981 = ~n8944 ^ n8980;
  assign n8982 = n8780 & n8813;
  assign n8983 = n8797 & n8812;
  assign n8984 = ~n8982 & ~n8983;
  assign n8985 = n8822 & n8829;
  assign n8986 = ~n8825 & ~n8828;
  assign n8987 = ~n8985 & ~n8986;
  assign n8988 = n8767 & ~n8770;
  assign n8989 = ~n8763 & ~n8766;
  assign n8990 = ~n8988 & ~n8989;
  assign n8991 = ~n8987 ^ ~n8990;
  assign n8992 = n8837 & n8840;
  assign n8993 = n8833 & n8836;
  assign n8994 = ~n8992 & ~n8993;
  assign n8995 = ~n8991 ^ ~n8994;
  assign n8996 = n8742 & ~n8743;
  assign n8997 = ~n8740 & ~n8741;
  assign n8998 = ~n8996 & ~n8997;
  assign n8999 = n8794 & ~n8795;
  assign n9000 = ~n8792 & ~n8793;
  assign n9001 = ~n8999 & ~n9000;
  assign n9002 = ~n8998 ^ ~n9001;
  assign n9003 = n8805 & ~n8806;
  assign n9004 = ~n8803 & ~n8804;
  assign n9005 = ~n9003 & ~n9004;
  assign n9006 = ~n9002 ^ ~n9005;
  assign n9007 = n8800 & ~n8801;
  assign n9008 = ~n8798 & ~n8799;
  assign n9009 = ~n9007 & ~n9008;
  assign n9010 = ~n8809 & ~pi37;
  assign n9011 = ~n9010 & pi38;
  assign n9012 = pi14 & pi62;
  assign n9013 = ~n9011 ^ ~n9012;
  assign n9014 = ~n9009 ^ n9013;
  assign n9015 = ~n9006 ^ n9014;
  assign n9016 = n8739 & ~n8744;
  assign n9017 = ~n8733 & ~n8738;
  assign n9018 = ~n9016 & ~n9017;
  assign n9019 = ~n9015 ^ n9018;
  assign n9020 = ~n8995 ^ n9019;
  assign n9021 = ~n8984 ^ ~n9020;
  assign n9022 = ~n8981 ^ ~n9021;
  assign n9023 = ~n8921 ^ ~n9022;
  assign n9024 = ~n8918 ^ n9023;
  assign po077 = n8881 ^ n9024;
  assign n9026 = n8711 & ~n8871;
  assign n9027 = n9024 & ~n8869;
  assign n9028 = ~n8866 & ~n9027;
  assign n9029 = ~n9026 & n9028;
  assign n9030 = ~n8871 & n9024;
  assign n9031 = ~n9030 & ~n8867;
  assign n9032 = ~n8711 & n9031;
  assign n9033 = ~n8870 & ~n9024;
  assign n9034 = ~n9032 & ~n9033;
  assign n9035 = ~n9029 & n9034;
  assign n9036 = n8918 & ~n9023;
  assign n9037 = ~n8884 & ~n8917;
  assign n9038 = ~n9036 & ~n9037;
  assign n9039 = n8921 & n9022;
  assign n9040 = n8981 & n9021;
  assign n9041 = ~n9039 & ~n9040;
  assign n9042 = n8913 & ~n8916;
  assign n9043 = ~n8887 & ~n8912;
  assign n9044 = ~n9042 & ~n9043;
  assign n9045 = n8894 & n8911;
  assign n9046 = ~n8890 & ~n8893;
  assign n9047 = ~n9045 & ~n9046;
  assign n9048 = n8973 & n8978;
  assign n9049 = ~n8968 & n8972;
  assign n9050 = ~n9048 & ~n9049;
  assign n9051 = ~n9009 & n9013;
  assign n9052 = ~n9011 & ~n9012;
  assign n9053 = ~n9051 & ~n9052;
  assign n9054 = n8958 & n8963;
  assign n9055 = n8952 & n8957;
  assign n9056 = ~n9054 & ~n9055;
  assign n9057 = ~n9053 ^ ~n9056;
  assign n9058 = ~n9050 ^ n9057;
  assign n9059 = ~n9047 ^ ~n9058;
  assign n9060 = n8991 & n8994;
  assign n9061 = ~n8987 & ~n8990;
  assign n9062 = ~n9060 & ~n9061;
  assign n9063 = n8950 & ~n8951;
  assign n9064 = ~n8948 & ~n8949;
  assign n9065 = ~n9063 & ~n9064;
  assign n9066 = pi21 & pi56;
  assign n9067 = pi20 & pi57;
  assign n9068 = ~n9066 ^ ~n9067;
  assign n9069 = pi19 & pi58;
  assign n9070 = ~n9068 ^ n9069;
  assign n9071 = pi29 & pi48;
  assign n9072 = pi28 & pi49;
  assign n9073 = ~n9071 ^ ~n9072;
  assign n9074 = pi27 & pi50;
  assign n9075 = ~n9073 ^ n9074;
  assign n9076 = ~n9070 ^ ~n9075;
  assign n9077 = ~n9065 ^ ~n9076;
  assign n9078 = pi31 & pi46;
  assign n9079 = pi30 & pi47;
  assign n9080 = ~n9078 ^ ~n9079;
  assign n9081 = pi14 & pi63;
  assign n9082 = ~n9080 ^ n9081;
  assign n9083 = pi37 & pi40;
  assign n9084 = pi36 & pi41;
  assign n9085 = ~n9083 ^ ~n9084;
  assign n9086 = pi35 & pi42;
  assign n9087 = ~n9085 ^ n9086;
  assign n9088 = ~n9082 ^ ~n9087;
  assign n9089 = pi15 & pi62;
  assign n9090 = ~pi38 & pi39;
  assign n9091 = ~n9089 ^ ~n9090;
  assign n9092 = ~n9088 ^ ~n9091;
  assign n9093 = ~n9077 ^ ~n9092;
  assign n9094 = ~n9062 ^ n9093;
  assign n9095 = ~n9059 ^ ~n9094;
  assign n9096 = n8965 & ~n8979;
  assign n9097 = n8947 & ~n8964;
  assign n9098 = ~n9096 & ~n9097;
  assign n9099 = n9002 & n9005;
  assign n9100 = n8998 & n9001;
  assign n9101 = ~n9099 & ~n9100;
  assign n9102 = n8955 & ~n8956;
  assign n9103 = ~n8953 & ~n8954;
  assign n9104 = ~n9102 & ~n9103;
  assign n9105 = pi17 & pi60;
  assign n9106 = pi18 & pi59;
  assign n9107 = ~n9105 ^ ~n9106;
  assign n9108 = ~n9104 ^ ~n9107;
  assign n9109 = ~n9101 ^ n9108;
  assign n9110 = n8938 & n8941;
  assign n9111 = n8934 & n8937;
  assign n9112 = ~n9110 & ~n9111;
  assign n9113 = ~n9109 ^ ~n9112;
  assign n9114 = n8905 & ~n8910;
  assign n9115 = ~n8899 & ~n8904;
  assign n9116 = ~n9114 & ~n9115;
  assign n9117 = n8902 & ~n8903;
  assign n9118 = ~n8900 & ~n8901;
  assign n9119 = ~n9117 & ~n9118;
  assign n9120 = n8976 & ~n8977;
  assign n9121 = ~n8974 & ~n8975;
  assign n9122 = ~n9120 & ~n9121;
  assign n9123 = ~n9119 ^ ~n9122;
  assign n9124 = n8970 & ~n8971;
  assign n9125 = ~n4492 & ~n8969;
  assign n9126 = ~n9124 & ~n9125;
  assign n9127 = ~n9123 ^ n9126;
  assign n9128 = ~n9116 ^ ~n9127;
  assign n9129 = n8908 & ~n8909;
  assign n9130 = ~n8906 & ~n8907;
  assign n9131 = ~n9129 & ~n9130;
  assign n9132 = n8897 & ~n8898;
  assign n9133 = ~n8895 & ~n8896;
  assign n9134 = ~n9132 & ~n9133;
  assign n9135 = ~n9131 ^ ~n9134;
  assign n9136 = n8961 & ~n8962;
  assign n9137 = ~n8959 & ~n8960;
  assign n9138 = ~n9136 & ~n9137;
  assign n9139 = ~n9135 ^ n9138;
  assign n9140 = ~n9128 ^ n9139;
  assign n9141 = ~n9113 ^ n9140;
  assign n9142 = ~n9098 ^ n9141;
  assign n9143 = ~n9095 ^ n9142;
  assign n9144 = ~n9044 ^ n9143;
  assign n9145 = n8944 & ~n8980;
  assign n9146 = ~n8924 & n8943;
  assign n9147 = ~n9145 & ~n9146;
  assign n9148 = n8984 & n9020;
  assign n9149 = n8995 & ~n9019;
  assign n9150 = ~n9148 & ~n9149;
  assign n9151 = n8931 & ~n8942;
  assign n9152 = n8927 & n8930;
  assign n9153 = ~n9151 & ~n9152;
  assign n9154 = pi34 & pi43;
  assign n9155 = ~n4542 ^ ~n9154;
  assign n9156 = pi22 & pi55;
  assign n9157 = ~n9155 ^ n9156;
  assign n9158 = pi33 & pi44;
  assign n9159 = pi32 & pi45;
  assign n9160 = ~n9158 ^ ~n9159;
  assign n9161 = pi16 & pi61;
  assign n9162 = ~n9160 ^ n9161;
  assign n9163 = ~n9157 ^ ~n9162;
  assign n9164 = pi25 & pi52;
  assign n9165 = pi24 & pi53;
  assign n9166 = ~n9164 ^ ~n9165;
  assign n9167 = pi23 & pi54;
  assign n9168 = ~n9166 ^ n9167;
  assign n9169 = ~n9163 ^ n9168;
  assign n9170 = ~n9153 ^ ~n9169;
  assign n9171 = n9015 & ~n9018;
  assign n9172 = n9006 & ~n9014;
  assign n9173 = ~n9171 & ~n9172;
  assign n9174 = ~n9170 ^ ~n9173;
  assign n9175 = ~n9150 ^ n9174;
  assign n9176 = ~n9147 ^ n9175;
  assign n9177 = ~n9144 ^ ~n9176;
  assign n9178 = ~n9041 ^ n9177;
  assign n9179 = ~n9038 ^ n9178;
  assign po078 = n9035 ^ ~n9179;
  assign n9181 = ~n9038 & n9041;
  assign n9182 = ~n9144 & ~n9176;
  assign n9183 = ~n9181 & ~n9182;
  assign n9184 = n9038 & ~n9041;
  assign n9185 = n9144 & n9176;
  assign n9186 = ~n9184 & ~n9185;
  assign n9187 = ~n9183 & n9186;
  assign n9188 = n9035 & ~n9187;
  assign n9189 = n9183 & ~n9186;
  assign n9190 = ~n9035 & ~n9189;
  assign n9191 = ~n9188 & ~n9190;
  assign n9192 = n9181 & n9182;
  assign n9193 = n9184 & n9185;
  assign n9194 = ~n9192 & ~n9193;
  assign n9195 = ~n9191 & n9194;
  assign n9196 = ~n9147 & n9175;
  assign n9197 = ~n9150 & n9174;
  assign n9198 = ~n9196 & ~n9197;
  assign n9199 = ~n9094 & ~n9092;
  assign n9200 = ~n9062 & ~n9077;
  assign n9201 = ~n9199 & ~n9200;
  assign n9202 = n9170 & n9173;
  assign n9203 = ~n9153 & ~n9169;
  assign n9204 = ~n9202 & ~n9203;
  assign n9205 = n9109 & n9112;
  assign n9206 = n9101 & ~n9108;
  assign n9207 = ~n9205 & ~n9206;
  assign n9208 = n9135 & ~n9138;
  assign n9209 = ~n9131 & ~n9134;
  assign n9210 = ~n9208 & ~n9209;
  assign n9211 = pi36 & pi42;
  assign n9212 = pi35 & pi43;
  assign n9213 = ~n9211 ^ ~n9212;
  assign n9214 = pi23 & pi55;
  assign n9215 = ~n9213 ^ n9214;
  assign n9216 = pi38 & pi40;
  assign n9217 = pi37 & pi41;
  assign n9218 = ~n9216 ^ ~n9217;
  assign n9219 = pi26 & pi52;
  assign n9220 = ~n9218 ^ n9219;
  assign n9221 = ~n9215 ^ ~n9220;
  assign n9222 = ~n9210 ^ ~n9221;
  assign n9223 = n9104 & n9107;
  assign n9224 = pi59 & pi60;
  assign n9225 = n2143 & n9224;
  assign n9226 = ~n9223 & ~n9225;
  assign n9227 = n9068 & ~n9069;
  assign n9228 = ~n9066 & ~n9067;
  assign n9229 = ~n9227 & ~n9228;
  assign n9230 = n9155 & ~n9156;
  assign n9231 = ~n4542 & ~n9154;
  assign n9232 = ~n9230 & ~n9231;
  assign n9233 = ~n9229 ^ ~n9232;
  assign n9234 = ~n9226 ^ n9233;
  assign n9235 = ~n9222 ^ ~n9234;
  assign n9236 = ~n9207 ^ n9235;
  assign n9237 = ~n9204 ^ n9236;
  assign n9238 = ~n9201 ^ ~n9237;
  assign n9239 = n9123 & ~n9126;
  assign n9240 = ~n9119 & ~n9122;
  assign n9241 = ~n9239 & ~n9240;
  assign n9242 = n9166 & ~n9167;
  assign n9243 = ~n9164 & ~n9165;
  assign n9244 = ~n9242 & ~n9243;
  assign n9245 = n9085 & ~n9086;
  assign n9246 = ~n9083 & ~n9084;
  assign n9247 = ~n9245 & ~n9246;
  assign n9248 = ~n9244 ^ ~n9247;
  assign n9249 = ~n9089 & ~pi38;
  assign n9250 = ~n9249 & pi39;
  assign n9251 = ~n9248 ^ n9250;
  assign n9252 = ~n9241 ^ n9251;
  assign n9253 = n9080 & ~n9081;
  assign n9254 = ~n9078 & ~n9079;
  assign n9255 = ~n9253 & ~n9254;
  assign n9256 = n9073 & ~n9074;
  assign n9257 = ~n9071 & ~n9072;
  assign n9258 = ~n9256 & ~n9257;
  assign n9259 = ~n9255 ^ ~n9258;
  assign n9260 = n9160 & ~n9161;
  assign n9261 = ~n9158 & ~n9159;
  assign n9262 = ~n9260 & ~n9261;
  assign n9263 = ~n9259 ^ ~n9262;
  assign n9264 = ~n9252 ^ n9263;
  assign n9265 = n9163 & ~n9168;
  assign n9266 = ~n9157 & ~n9162;
  assign n9267 = ~n9265 & ~n9266;
  assign n9268 = n9088 & n9091;
  assign n9269 = ~n9082 & ~n9087;
  assign n9270 = ~n9268 & ~n9269;
  assign n9271 = ~n9267 ^ ~n9270;
  assign n9272 = n9065 & n9076;
  assign n9273 = ~n9070 & ~n9075;
  assign n9274 = ~n9272 & ~n9273;
  assign n9275 = ~n9271 ^ ~n9274;
  assign n9276 = ~n9264 ^ ~n9275;
  assign n9277 = n9128 & ~n9139;
  assign n9278 = ~n9116 & ~n9127;
  assign n9279 = ~n9277 & ~n9278;
  assign n9280 = ~n9276 ^ ~n9279;
  assign n9281 = ~n9238 ^ n9280;
  assign n9282 = ~n9198 ^ n9281;
  assign n9283 = n9059 & n9094;
  assign n9284 = n9047 & n9058;
  assign n9285 = ~n9283 & ~n9284;
  assign n9286 = ~n9098 & n9141;
  assign n9287 = ~n9113 & n9140;
  assign n9288 = ~n9286 & ~n9287;
  assign n9289 = ~n9285 ^ n9288;
  assign n9290 = ~n9050 & n9057;
  assign n9291 = ~n9053 & ~n9056;
  assign n9292 = ~n9290 & ~n9291;
  assign n9293 = pi34 & pi44;
  assign n9294 = pi33 & pi45;
  assign n9295 = ~n9293 ^ ~n9294;
  assign n9296 = pi32 & pi46;
  assign n9297 = ~n9295 ^ n9296;
  assign n9298 = pi31 & pi47;
  assign n9299 = pi30 & pi48;
  assign n9300 = ~n9298 ^ ~n9299;
  assign n9301 = pi20 & pi58;
  assign n9302 = ~n9300 ^ n9301;
  assign n9303 = ~n9297 ^ ~n9302;
  assign n9304 = pi25 & pi53;
  assign n9305 = pi24 & pi54;
  assign n9306 = ~n9304 ^ ~n9305;
  assign n9307 = pi22 & pi56;
  assign n9308 = ~n9306 ^ n9307;
  assign n9309 = ~n9303 ^ n9308;
  assign n9310 = pi21 & pi57;
  assign n9311 = pi19 & pi59;
  assign n9312 = ~n9310 ^ ~n9311;
  assign n9313 = pi18 & pi60;
  assign n9314 = ~n9312 ^ n9313;
  assign n9315 = pi17 & pi61;
  assign n9316 = pi16 & pi62;
  assign n9317 = ~n9315 ^ ~n9316;
  assign n9318 = pi15 & pi63;
  assign n9319 = ~n9317 ^ n9318;
  assign n9320 = ~n9314 ^ ~n9319;
  assign n9321 = pi29 & pi49;
  assign n9322 = pi28 & pi50;
  assign n9323 = ~n9321 ^ ~n9322;
  assign n9324 = pi27 & pi51;
  assign n9325 = ~n9323 ^ n9324;
  assign n9326 = ~n9320 ^ ~n9325;
  assign n9327 = ~n9309 ^ n9326;
  assign n9328 = ~n9292 ^ ~n9327;
  assign n9329 = ~n9289 ^ ~n9328;
  assign n9330 = ~n9282 ^ n9329;
  assign n9331 = ~n9044 & n9143;
  assign n9332 = n9095 & ~n9142;
  assign n9333 = ~n9331 & ~n9332;
  assign n9334 = ~n9330 ^ n9333;
  assign po079 = n9195 ^ ~n9334;
  assign n9336 = n9035 & ~n9184;
  assign n9337 = ~n9334 & ~n9185;
  assign n9338 = ~n9181 & ~n9337;
  assign n9339 = ~n9336 & n9338;
  assign n9340 = ~n9184 & ~n9334;
  assign n9341 = ~n9340 & ~n9182;
  assign n9342 = ~n9035 & n9341;
  assign n9343 = ~n9183 & ~n9185;
  assign n9344 = ~n9343 & n9334;
  assign n9345 = ~n9342 & ~n9344;
  assign n9346 = ~n9339 & n9345;
  assign n9347 = n9330 & ~n9333;
  assign n9348 = n9282 & ~n9329;
  assign n9349 = ~n9347 & ~n9348;
  assign n9350 = ~n9198 & n9281;
  assign n9351 = ~n9238 & n9280;
  assign n9352 = ~n9350 & ~n9351;
  assign n9353 = n9289 & n9328;
  assign n9354 = n9285 & ~n9288;
  assign n9355 = ~n9353 & ~n9354;
  assign n9356 = n9201 & n9237;
  assign n9357 = n9204 & ~n9236;
  assign n9358 = ~n9356 & ~n9357;
  assign n9359 = n9210 & n9221;
  assign n9360 = ~n9215 & ~n9220;
  assign n9361 = ~n9359 & ~n9360;
  assign n9362 = n9312 & ~n9313;
  assign n9363 = ~n9310 & ~n9311;
  assign n9364 = ~n9362 & ~n9363;
  assign n9365 = n9323 & ~n9324;
  assign n9366 = ~n9321 & ~n9322;
  assign n9367 = ~n9365 & ~n9366;
  assign n9368 = ~n9364 ^ ~n9367;
  assign n9369 = n9306 & ~n9307;
  assign n9370 = ~n9304 & ~n9305;
  assign n9371 = ~n9369 & ~n9370;
  assign n9372 = ~n9368 ^ ~n9371;
  assign n9373 = ~n9361 ^ n9372;
  assign n9374 = ~n9226 & n9233;
  assign n9375 = n9229 & n9232;
  assign n9376 = ~n9374 & ~n9375;
  assign n9377 = pi36 & pi43;
  assign n9378 = ~n4826 ^ ~n9377;
  assign n9379 = pi23 & pi56;
  assign n9380 = ~n9378 ^ n9379;
  assign n9381 = pi35 & pi44;
  assign n9382 = pi34 & pi45;
  assign n9383 = ~n9381 ^ ~n9382;
  assign n9384 = pi16 & pi63;
  assign n9385 = ~n9383 ^ n9384;
  assign n9386 = ~n9380 ^ ~n9385;
  assign n9387 = ~n9376 ^ n9386;
  assign n9388 = ~n9373 ^ n9387;
  assign n9389 = n9218 & ~n9219;
  assign n9390 = ~n9216 & ~n9217;
  assign n9391 = ~n9389 & ~n9390;
  assign n9392 = pi18 & pi61;
  assign n9393 = ~n9391 ^ ~n9392;
  assign n9394 = n9213 & ~n9214;
  assign n9395 = ~n9211 & ~n9212;
  assign n9396 = ~n9394 & ~n9395;
  assign n9397 = ~n9393 ^ ~n9396;
  assign n9398 = n9303 & ~n9308;
  assign n9399 = ~n9297 & ~n9302;
  assign n9400 = ~n9398 & ~n9399;
  assign n9401 = ~n9397 ^ n9400;
  assign n9402 = n9300 & ~n9301;
  assign n9403 = ~n9298 & ~n9299;
  assign n9404 = ~n9402 & ~n9403;
  assign n9405 = n9295 & ~n9296;
  assign n9406 = ~n9293 & ~n9294;
  assign n9407 = ~n9405 & ~n9406;
  assign n9408 = ~n9404 ^ ~n9407;
  assign n9409 = n9317 & ~n9318;
  assign n9410 = ~n9315 & ~n9316;
  assign n9411 = ~n9409 & ~n9410;
  assign n9412 = ~n9408 ^ ~n9411;
  assign n9413 = ~n9401 ^ n9412;
  assign n9414 = ~n9388 ^ ~n9413;
  assign n9415 = n9328 & n9326;
  assign n9416 = ~n9292 & ~n9309;
  assign n9417 = ~n9415 & ~n9416;
  assign n9418 = ~n9414 ^ n9417;
  assign n9419 = ~n9358 ^ n9418;
  assign n9420 = ~n9355 ^ ~n9419;
  assign n9421 = ~n9352 ^ ~n9420;
  assign n9422 = n9280 & ~n9264;
  assign n9423 = ~n9279 & ~n9275;
  assign n9424 = ~n9422 & ~n9423;
  assign n9425 = n9252 & ~n9263;
  assign n9426 = ~n9241 & n9251;
  assign n9427 = ~n9425 & ~n9426;
  assign n9428 = pi30 & pi49;
  assign n9429 = pi29 & pi50;
  assign n9430 = ~n9428 ^ ~n9429;
  assign n9431 = pi22 & pi57;
  assign n9432 = ~n9430 ^ n9431;
  assign n9433 = pi33 & pi46;
  assign n9434 = pi32 & pi47;
  assign n9435 = ~n9433 ^ ~n9434;
  assign n9436 = pi31 & pi48;
  assign n9437 = ~n9435 ^ n9436;
  assign n9438 = ~n9432 ^ ~n9437;
  assign n9439 = pi21 & pi58;
  assign n9440 = pi20 & pi59;
  assign n9441 = ~n9439 ^ ~n9440;
  assign n9442 = pi19 & pi60;
  assign n9443 = ~n9441 ^ n9442;
  assign n9444 = ~n9438 ^ n9443;
  assign n9445 = ~n9427 ^ ~n9444;
  assign n9446 = pi39 & pi40;
  assign n9447 = pi38 & pi41;
  assign n9448 = ~n9446 ^ ~n9447;
  assign n9449 = pi37 & pi42;
  assign n9450 = ~n9448 ^ n9449;
  assign n9451 = pi17 & pi62;
  assign n9452 = pi28 & pi51;
  assign n9453 = ~n9451 ^ n9452;
  assign n9454 = ~n9453 ^ pi40;
  assign n9455 = ~n9450 ^ n9454;
  assign n9456 = pi25 & pi54;
  assign n9457 = ~n4990 ^ ~n9456;
  assign n9458 = pi24 & pi55;
  assign n9459 = ~n9457 ^ n9458;
  assign n9460 = ~n9455 ^ n9459;
  assign n9461 = ~n9445 ^ n9460;
  assign n9462 = ~n9424 ^ ~n9461;
  assign n9463 = ~n9236 & ~n9234;
  assign n9464 = ~n9207 & ~n9222;
  assign n9465 = ~n9463 & ~n9464;
  assign n9466 = n9271 & n9274;
  assign n9467 = n9267 & n9270;
  assign n9468 = ~n9466 & ~n9467;
  assign n9469 = n9248 & ~n9250;
  assign n9470 = ~n9244 & ~n9247;
  assign n9471 = ~n9469 & ~n9470;
  assign n9472 = n9320 & n9325;
  assign n9473 = n9314 & n9319;
  assign n9474 = ~n9472 & ~n9473;
  assign n9475 = ~n9471 ^ ~n9474;
  assign n9476 = n9259 & n9262;
  assign n9477 = n9255 & n9258;
  assign n9478 = ~n9476 & ~n9477;
  assign n9479 = ~n9475 ^ n9478;
  assign n9480 = ~n9468 ^ ~n9479;
  assign n9481 = ~n9465 ^ ~n9480;
  assign n9482 = ~n9462 ^ n9481;
  assign n9483 = ~n9421 ^ n9482;
  assign n9484 = ~n9349 ^ ~n9483;
  assign po080 = n9346 ^ n9484;
  assign n9486 = n9349 & n9483;
  assign n9487 = ~n9346 & ~n9486;
  assign n9488 = ~n9349 & ~n9483;
  assign n9489 = ~n9487 & ~n9488;
  assign n9490 = n9421 & ~n9482;
  assign n9491 = n9352 & n9420;
  assign n9492 = ~n9490 & ~n9491;
  assign n9493 = ~n9420 & ~n9418;
  assign n9494 = ~n9355 & ~n9358;
  assign n9495 = ~n9493 & ~n9494;
  assign n9496 = n9462 & ~n9481;
  assign n9497 = n9424 & n9461;
  assign n9498 = ~n9496 & ~n9497;
  assign n9499 = n9445 & ~n9460;
  assign n9500 = ~n9427 & ~n9444;
  assign n9501 = ~n9499 & ~n9500;
  assign n9502 = ~n9376 & n9386;
  assign n9503 = ~n9380 & ~n9385;
  assign n9504 = ~n9502 & ~n9503;
  assign n9505 = n9475 & ~n9478;
  assign n9506 = n9471 & n9474;
  assign n9507 = ~n9505 & ~n9506;
  assign n9508 = ~n9504 ^ ~n9507;
  assign n9509 = n9457 & ~n9458;
  assign n9510 = ~n4990 & ~n9456;
  assign n9511 = ~n9509 & ~n9510;
  assign n9512 = n9383 & ~n9384;
  assign n9513 = ~n9381 & ~n9382;
  assign n9514 = ~n9512 & ~n9513;
  assign n9515 = ~n9511 ^ ~n9514;
  assign n9516 = n9378 & ~n9379;
  assign n9517 = ~n4826 & ~n9377;
  assign n9518 = ~n9516 & ~n9517;
  assign n9519 = ~n9515 ^ ~n9518;
  assign n9520 = ~n9508 ^ ~n9519;
  assign n9521 = n9430 & ~n9431;
  assign n9522 = ~n9428 & ~n9429;
  assign n9523 = ~n9521 & ~n9522;
  assign n9524 = n9435 & ~n9436;
  assign n9525 = ~n9433 & ~n9434;
  assign n9526 = ~n9524 & ~n9525;
  assign n9527 = ~n9523 ^ ~n9526;
  assign n9528 = n9441 & ~n9442;
  assign n9529 = ~n9439 & ~n9440;
  assign n9530 = ~n9528 & ~n9529;
  assign n9531 = ~n9527 ^ ~n9530;
  assign n9532 = n9455 & ~n9459;
  assign n9533 = ~n9450 & n9454;
  assign n9534 = ~n9532 & ~n9533;
  assign n9535 = ~n9531 ^ n9534;
  assign n9536 = n9438 & ~n9443;
  assign n9537 = ~n9432 & ~n9437;
  assign n9538 = ~n9536 & ~n9537;
  assign n9539 = ~n9535 ^ ~n9538;
  assign n9540 = ~n9520 ^ n9539;
  assign n9541 = ~n9501 ^ ~n9540;
  assign n9542 = n9373 & ~n9387;
  assign n9543 = n9361 & ~n9372;
  assign n9544 = ~n9542 & ~n9543;
  assign n9545 = n9401 & ~n9412;
  assign n9546 = ~n9397 & n9400;
  assign n9547 = ~n9545 & ~n9546;
  assign n9548 = n9368 & n9371;
  assign n9549 = n9364 & n9367;
  assign n9550 = ~n9548 & ~n9549;
  assign n9551 = n9408 & n9411;
  assign n9552 = n9404 & n9407;
  assign n9553 = ~n9551 & ~n9552;
  assign n9554 = ~n9550 ^ ~n9553;
  assign n9555 = n9393 & n9396;
  assign n9556 = n9391 & n9392;
  assign n9557 = ~n9555 & ~n9556;
  assign n9558 = ~n9554 ^ n9557;
  assign n9559 = ~n9547 ^ ~n9558;
  assign n9560 = ~n9544 ^ ~n9559;
  assign n9561 = ~n9541 ^ ~n9560;
  assign n9562 = ~n9498 ^ n9561;
  assign n9563 = n9465 & n9480;
  assign n9564 = n9468 & n9479;
  assign n9565 = ~n9563 & ~n9564;
  assign n9566 = n9414 & ~n9417;
  assign n9567 = n9388 & n9413;
  assign n9568 = ~n9566 & ~n9567;
  assign n9569 = n7524 & pi51;
  assign n9570 = ~n9569 & ~n9451;
  assign n9571 = ~n9452 & ~pi40;
  assign n9572 = ~n9570 & ~n9571;
  assign n9573 = pi18 & pi62;
  assign n9574 = pi19 & pi61;
  assign n9575 = ~n9573 ^ ~n9574;
  assign n9576 = ~n9572 ^ ~n9575;
  assign n9577 = pi36 & pi44;
  assign n9578 = pi35 & pi45;
  assign n9579 = ~n9577 ^ ~n9578;
  assign n9580 = pi34 & pi46;
  assign n9581 = ~n9579 ^ n9580;
  assign n9582 = pi33 & pi47;
  assign n9583 = pi29 & pi51;
  assign n9584 = ~n9582 ^ ~n9583;
  assign n9585 = pi17 & pi63;
  assign n9586 = ~n9584 ^ n9585;
  assign n9587 = ~n9581 ^ ~n9586;
  assign n9588 = ~n9576 ^ n9587;
  assign n9589 = pi39 & pi41;
  assign n9590 = pi28 & pi52;
  assign n9591 = ~n9589 ^ ~n9590;
  assign n9592 = pi27 & pi53;
  assign n9593 = ~n9591 ^ n9592;
  assign n9594 = pi38 & pi42;
  assign n9595 = pi37 & pi43;
  assign n9596 = ~n9594 ^ ~n9595;
  assign n9597 = pi25 & pi55;
  assign n9598 = ~n9596 ^ n9597;
  assign n9599 = ~n9593 ^ ~n9598;
  assign n9600 = pi26 & pi54;
  assign n9601 = pi24 & pi56;
  assign n9602 = ~n9600 ^ ~n9601;
  assign n9603 = pi23 & pi57;
  assign n9604 = ~n9602 ^ n9603;
  assign n9605 = ~n9599 ^ n9604;
  assign n9606 = ~n9588 ^ n9605;
  assign n9607 = n9448 & ~n9449;
  assign n9608 = ~n9446 & ~n9447;
  assign n9609 = ~n9607 & ~n9608;
  assign n9610 = pi22 & pi58;
  assign n9611 = pi21 & pi59;
  assign n9612 = ~n9610 ^ ~n9611;
  assign n9613 = pi20 & pi60;
  assign n9614 = ~n9612 ^ n9613;
  assign n9615 = pi32 & pi48;
  assign n9616 = pi31 & pi49;
  assign n9617 = ~n9615 ^ ~n9616;
  assign n9618 = pi30 & pi50;
  assign n9619 = ~n9617 ^ n9618;
  assign n9620 = ~n9614 ^ ~n9619;
  assign n9621 = ~n9609 ^ ~n9620;
  assign n9622 = ~n9606 ^ ~n9621;
  assign n9623 = ~n9568 ^ ~n9622;
  assign n9624 = ~n9565 ^ n9623;
  assign n9625 = ~n9562 ^ ~n9624;
  assign n9626 = ~n9495 ^ n9625;
  assign n9627 = ~n9492 ^ n9626;
  assign po081 = ~n9489 ^ n9627;
  assign n9629 = ~n9562 & n9624;
  assign n9630 = n9495 & ~n9629;
  assign n9631 = n9492 & n9630;
  assign n9632 = n9562 & ~n9624;
  assign n9633 = ~n9631 & ~n9632;
  assign n9634 = ~n9492 & ~n9495;
  assign n9635 = ~n9633 & ~n9634;
  assign n9636 = ~n9489 & n9635;
  assign n9637 = n9495 & n9632;
  assign n9638 = n9492 & n9637;
  assign n9639 = ~n9495 & n9629;
  assign n9640 = ~n9492 & n9639;
  assign n9641 = ~n9638 & ~n9640;
  assign n9642 = ~n9636 & n9641;
  assign n9643 = n9492 & ~n9639;
  assign n9644 = ~n9630 & ~n9632;
  assign n9645 = ~n9643 & n9644;
  assign n9646 = n9489 & n9645;
  assign n9647 = n9642 & ~n9646;
  assign n9648 = ~n9565 & n9623;
  assign n9649 = n9568 & n9622;
  assign n9650 = ~n9648 & ~n9649;
  assign n9651 = n9606 & n9621;
  assign n9652 = ~n9588 & n9605;
  assign n9653 = ~n9651 & ~n9652;
  assign n9654 = n9609 & n9620;
  assign n9655 = ~n9614 & ~n9619;
  assign n9656 = ~n9654 & ~n9655;
  assign n9657 = n9602 & ~n9603;
  assign n9658 = ~n9600 & ~n9601;
  assign n9659 = ~n9657 & ~n9658;
  assign n9660 = n9591 & ~n9592;
  assign n9661 = ~n9589 & ~n9590;
  assign n9662 = ~n9660 & ~n9661;
  assign n9663 = ~n9659 ^ ~n9662;
  assign n9664 = n9596 & ~n9597;
  assign n9665 = ~n9594 & ~n9595;
  assign n9666 = ~n9664 & ~n9665;
  assign n9667 = ~n9663 ^ ~n9666;
  assign n9668 = ~n9656 ^ n9667;
  assign n9669 = n9599 & ~n9604;
  assign n9670 = ~n9593 & ~n9598;
  assign n9671 = ~n9669 & ~n9670;
  assign n9672 = ~n9668 ^ n9671;
  assign n9673 = ~n9653 ^ n9672;
  assign n9674 = n9572 & n9575;
  assign n9675 = n2386 & n8820;
  assign n9676 = ~n9674 & ~n9675;
  assign n9677 = n9579 & ~n9580;
  assign n9678 = ~n9577 & ~n9578;
  assign n9679 = ~n9677 & ~n9678;
  assign n9680 = pi32 & pi49;
  assign n9681 = pi31 & pi50;
  assign n9682 = ~n9680 ^ ~n9681;
  assign n9683 = pi30 & pi51;
  assign n9684 = ~n9682 ^ n9683;
  assign n9685 = ~n9679 ^ n9684;
  assign n9686 = ~n9676 ^ ~n9685;
  assign n9687 = ~n9576 & n9587;
  assign n9688 = n9581 & n9586;
  assign n9689 = ~n9687 & ~n9688;
  assign n9690 = ~n9686 ^ n9689;
  assign n9691 = n9584 & ~n9585;
  assign n9692 = ~n9582 & ~n9583;
  assign n9693 = ~n9691 & ~n9692;
  assign n9694 = n9612 & ~n9613;
  assign n9695 = ~n9610 & ~n9611;
  assign n9696 = ~n9694 & ~n9695;
  assign n9697 = ~n9693 ^ ~n9696;
  assign n9698 = n9617 & ~n9618;
  assign n9699 = ~n9615 & ~n9616;
  assign n9700 = ~n9698 & ~n9699;
  assign n9701 = ~n9697 ^ ~n9700;
  assign n9702 = ~n9690 ^ ~n9701;
  assign n9703 = ~n9673 ^ n9702;
  assign n9704 = ~n9650 ^ ~n9703;
  assign n9705 = n9508 & n9519;
  assign n9706 = ~n9504 & ~n9507;
  assign n9707 = ~n9705 & ~n9706;
  assign n9708 = n9535 & n9538;
  assign n9709 = ~n9531 & n9534;
  assign n9710 = ~n9708 & ~n9709;
  assign n9711 = n9527 & n9530;
  assign n9712 = n9523 & n9526;
  assign n9713 = ~n9711 & ~n9712;
  assign n9714 = pi39 & pi42;
  assign n9715 = pi38 & pi43;
  assign n9716 = ~n9714 ^ ~n9715;
  assign n9717 = pi27 & pi54;
  assign n9718 = ~n9716 ^ n9717;
  assign n9719 = ~n9713 ^ ~n9718;
  assign n9720 = n9515 & n9518;
  assign n9721 = n9511 & n9514;
  assign n9722 = ~n9720 & ~n9721;
  assign n9723 = ~n9719 ^ ~n9722;
  assign n9724 = ~n9710 ^ n9723;
  assign n9725 = ~n9707 ^ n9724;
  assign n9726 = ~n9704 ^ n9725;
  assign n9727 = n9562 & n9541;
  assign n9728 = n9498 & n9560;
  assign n9729 = ~n9727 & ~n9728;
  assign n9730 = ~n9726 ^ ~n9729;
  assign n9731 = n9501 & n9540;
  assign n9732 = n9520 & ~n9539;
  assign n9733 = ~n9731 & ~n9732;
  assign n9734 = n9554 & ~n9557;
  assign n9735 = ~n9550 & ~n9553;
  assign n9736 = ~n9734 & ~n9735;
  assign n9737 = pi29 & pi52;
  assign n9738 = ~n5283 ^ ~n9737;
  assign n9739 = pi26 & pi55;
  assign n9740 = ~n9738 ^ n9739;
  assign n9741 = pi37 & pi44;
  assign n9742 = pi36 & pi45;
  assign n9743 = ~n9741 ^ ~n9742;
  assign n9744 = pi35 & pi46;
  assign n9745 = ~n9743 ^ n9744;
  assign n9746 = ~n9740 ^ ~n9745;
  assign n9747 = pi21 & pi60;
  assign n9748 = pi20 & pi61;
  assign n9749 = ~n9747 ^ ~n9748;
  assign n9750 = pi18 & pi63;
  assign n9751 = ~n9749 ^ n9750;
  assign n9752 = ~n9746 ^ n9751;
  assign n9753 = ~n9736 ^ n9752;
  assign n9754 = pi34 & pi47;
  assign n9755 = pi33 & pi48;
  assign n9756 = ~n9754 ^ ~n9755;
  assign n9757 = pi24 & pi57;
  assign n9758 = ~n9756 ^ n9757;
  assign n9759 = pi25 & pi56;
  assign n9760 = pi23 & pi58;
  assign n9761 = ~n9759 ^ ~n9760;
  assign n9762 = pi22 & pi59;
  assign n9763 = ~n9761 ^ n9762;
  assign n9764 = ~n9758 ^ ~n9763;
  assign n9765 = pi19 & pi62;
  assign n9766 = ~pi40 & pi41;
  assign n9767 = ~n9765 ^ ~n9766;
  assign n9768 = ~n9764 ^ ~n9767;
  assign n9769 = ~n9753 ^ n9768;
  assign n9770 = ~n9733 ^ ~n9769;
  assign n9771 = n9544 & n9559;
  assign n9772 = n9547 & n9558;
  assign n9773 = ~n9771 & ~n9772;
  assign n9774 = ~n9770 ^ n9773;
  assign n9775 = ~n9730 ^ ~n9774;
  assign po082 = n9647 ^ n9775;
  assign n9777 = n9492 & n9495;
  assign n9778 = ~n9777 & ~n9488;
  assign n9779 = ~n9487 & n9778;
  assign n9780 = ~n9779 & ~n9634;
  assign n9781 = ~n9775 & ~n9629;
  assign n9782 = ~n9780 & ~n9781;
  assign n9783 = ~n9634 & ~n9775;
  assign n9784 = ~n9783 & ~n9632;
  assign n9785 = n9489 & n9784;
  assign n9786 = n9633 & n9775;
  assign n9787 = ~n9785 & ~n9786;
  assign n9788 = ~n9782 & n9787;
  assign n9789 = n9730 & n9774;
  assign n9790 = ~n9726 & ~n9729;
  assign n9791 = ~n9789 & ~n9790;
  assign n9792 = n9704 & ~n9725;
  assign n9793 = n9650 & n9703;
  assign n9794 = ~n9792 & ~n9793;
  assign n9795 = n9770 & ~n9773;
  assign n9796 = ~n9733 & ~n9769;
  assign n9797 = ~n9795 & ~n9796;
  assign n9798 = n9753 & ~n9768;
  assign n9799 = n9736 & ~n9752;
  assign n9800 = ~n9798 & ~n9799;
  assign n9801 = n9676 & n9685;
  assign n9802 = ~n9679 & n9684;
  assign n9803 = ~n9801 & ~n9802;
  assign n9804 = n9716 & ~n9717;
  assign n9805 = ~n9714 & ~n9715;
  assign n9806 = ~n9804 & ~n9805;
  assign n9807 = pi19 & pi63;
  assign n9808 = ~n9806 ^ ~n9807;
  assign n9809 = ~n9765 & ~pi40;
  assign n9810 = ~n9809 & pi41;
  assign n9811 = ~n9808 ^ ~n9810;
  assign n9812 = n9764 & n9767;
  assign n9813 = ~n9758 & ~n9763;
  assign n9814 = ~n9812 & ~n9813;
  assign n9815 = ~n9811 ^ n9814;
  assign n9816 = ~n9803 ^ ~n9815;
  assign n9817 = ~n9800 ^ ~n9816;
  assign n9818 = n9761 & ~n9762;
  assign n9819 = ~n9759 & ~n9760;
  assign n9820 = ~n9818 & ~n9819;
  assign n9821 = n9749 & ~n9750;
  assign n9822 = ~n9747 & ~n9748;
  assign n9823 = ~n9821 & ~n9822;
  assign n9824 = ~n9820 ^ ~n9823;
  assign n9825 = n9743 & ~n9744;
  assign n9826 = ~n9741 & ~n9742;
  assign n9827 = ~n9825 & ~n9826;
  assign n9828 = ~n9824 ^ ~n9827;
  assign n9829 = n9746 & ~n9751;
  assign n9830 = ~n9740 & ~n9745;
  assign n9831 = ~n9829 & ~n9830;
  assign n9832 = ~n9828 ^ n9831;
  assign n9833 = n9738 & ~n9739;
  assign n9834 = ~n5283 & ~n9737;
  assign n9835 = ~n9833 & ~n9834;
  assign n9836 = n9756 & ~n9757;
  assign n9837 = ~n9754 & ~n9755;
  assign n9838 = ~n9836 & ~n9837;
  assign n9839 = ~n9835 ^ ~n9838;
  assign n9840 = n9682 & ~n9683;
  assign n9841 = ~n9680 & ~n9681;
  assign n9842 = ~n9840 & ~n9841;
  assign n9843 = ~n9839 ^ n9842;
  assign n9844 = ~n9832 ^ ~n9843;
  assign n9845 = ~n9817 ^ n9844;
  assign n9846 = n9690 & n9701;
  assign n9847 = ~n9686 & n9689;
  assign n9848 = ~n9846 & ~n9847;
  assign n9849 = n9668 & ~n9671;
  assign n9850 = ~n9656 & n9667;
  assign n9851 = ~n9849 & ~n9850;
  assign n9852 = n9663 & n9666;
  assign n9853 = n9659 & n9662;
  assign n9854 = ~n9852 & ~n9853;
  assign n9855 = ~n5286 ^ ~n5477;
  assign n9856 = pi25 & pi57;
  assign n9857 = ~n9855 ^ n9856;
  assign n9858 = ~n9854 ^ ~n9857;
  assign n9859 = n9697 & n9700;
  assign n9860 = n9693 & n9696;
  assign n9861 = ~n9859 & ~n9860;
  assign n9862 = ~n9858 ^ ~n9861;
  assign n9863 = ~n9851 ^ ~n9862;
  assign n9864 = ~n9848 ^ n9863;
  assign n9865 = ~n9845 ^ ~n9864;
  assign n9866 = ~n9797 ^ ~n9865;
  assign n9867 = ~n9707 & n9724;
  assign n9868 = n9710 & ~n9723;
  assign n9869 = ~n9867 & ~n9868;
  assign n9870 = n9719 & n9722;
  assign n9871 = n9713 & n9718;
  assign n9872 = ~n9870 & ~n9871;
  assign n9873 = pi40 & pi42;
  assign n9874 = pi30 & pi52;
  assign n9875 = ~n9873 ^ ~n9874;
  assign n9876 = pi29 & pi53;
  assign n9877 = ~n9875 ^ n9876;
  assign n9878 = pi37 & pi45;
  assign n9879 = pi36 & pi46;
  assign n9880 = ~n9878 ^ ~n9879;
  assign n9881 = pi35 & pi47;
  assign n9882 = ~n9880 ^ n9881;
  assign n9883 = ~n9877 ^ ~n9882;
  assign n9884 = pi39 & pi43;
  assign n9885 = pi38 & pi44;
  assign n9886 = ~n9884 ^ ~n9885;
  assign n9887 = pi26 & pi56;
  assign n9888 = ~n9886 ^ n9887;
  assign n9889 = ~n9883 ^ n9888;
  assign n9890 = pi31 & pi51;
  assign n9891 = pi21 & pi61;
  assign n9892 = ~n9890 ^ ~n9891;
  assign n9893 = pi20 & pi62;
  assign n9894 = ~n9892 ^ n9893;
  assign n9895 = pi24 & pi58;
  assign n9896 = pi23 & pi59;
  assign n9897 = ~n9895 ^ ~n9896;
  assign n9898 = pi22 & pi60;
  assign n9899 = ~n9897 ^ n9898;
  assign n9900 = ~n9894 ^ ~n9899;
  assign n9901 = pi34 & pi48;
  assign n9902 = pi33 & pi49;
  assign n9903 = ~n9901 ^ ~n9902;
  assign n9904 = pi32 & pi50;
  assign n9905 = ~n9903 ^ n9904;
  assign n9906 = ~n9900 ^ n9905;
  assign n9907 = ~n9889 ^ ~n9906;
  assign n9908 = ~n9872 ^ ~n9907;
  assign n9909 = ~n9869 ^ n9908;
  assign n9910 = n9673 & ~n9702;
  assign n9911 = n9653 & ~n9672;
  assign n9912 = ~n9910 & ~n9911;
  assign n9913 = ~n9909 ^ n9912;
  assign n9914 = ~n9866 ^ n9913;
  assign n9915 = ~n9794 ^ n9914;
  assign n9916 = ~n9791 ^ n9915;
  assign po083 = ~n9788 ^ n9916;
  assign n9918 = ~n9794 & n9913;
  assign n9919 = ~n9918 & ~n9866;
  assign n9920 = n9794 & ~n9913;
  assign n9921 = ~n9919 & ~n9920;
  assign n9922 = n9918 & n9866;
  assign n9923 = ~n9791 & ~n9922;
  assign n9924 = n9921 & ~n9923;
  assign n9925 = n9788 & n9924;
  assign n9926 = n9791 & n9922;
  assign n9927 = n9920 & ~n9866;
  assign n9928 = ~n9791 & n9927;
  assign n9929 = ~n9926 & ~n9928;
  assign n9930 = ~n9925 & n9929;
  assign n9931 = n9791 & ~n9927;
  assign n9932 = ~n9921 & ~n9931;
  assign n9933 = ~n9788 & n9932;
  assign n9934 = n9930 & ~n9933;
  assign n9935 = n9797 & n9865;
  assign n9936 = ~n9845 & ~n9864;
  assign n9937 = ~n9935 & ~n9936;
  assign n9938 = n9909 & ~n9912;
  assign n9939 = n9869 & ~n9908;
  assign n9940 = ~n9938 & ~n9939;
  assign n9941 = n9872 & n9907;
  assign n9942 = n9889 & n9906;
  assign n9943 = ~n9941 & ~n9942;
  assign n9944 = n9832 & n9843;
  assign n9945 = ~n9828 & n9831;
  assign n9946 = ~n9944 & ~n9945;
  assign n9947 = n9892 & ~n9893;
  assign n9948 = ~n9890 & ~n9891;
  assign n9949 = ~n9947 & ~n9948;
  assign n9950 = n9903 & ~n9904;
  assign n9951 = ~n9901 & ~n9902;
  assign n9952 = ~n9950 & ~n9951;
  assign n9953 = ~n9949 ^ ~n9952;
  assign n9954 = n9855 & ~n9856;
  assign n9955 = ~n5286 & ~n5477;
  assign n9956 = ~n9954 & ~n9955;
  assign n9957 = ~n9953 ^ ~n9956;
  assign n9958 = n9880 & ~n9881;
  assign n9959 = ~n9878 & ~n9879;
  assign n9960 = ~n9958 & ~n9959;
  assign n9961 = n9886 & ~n9887;
  assign n9962 = ~n9884 & ~n9885;
  assign n9963 = ~n9961 & ~n9962;
  assign n9964 = ~n9960 ^ ~n9963;
  assign n9965 = n9897 & ~n9898;
  assign n9966 = ~n9895 & ~n9896;
  assign n9967 = ~n9965 & ~n9966;
  assign n9968 = ~n9964 ^ n9967;
  assign n9969 = ~n9957 ^ n9968;
  assign n9970 = n9883 & ~n9888;
  assign n9971 = ~n9877 & ~n9882;
  assign n9972 = ~n9970 & ~n9971;
  assign n9973 = ~n9969 ^ ~n9972;
  assign n9974 = ~n9946 ^ n9973;
  assign n9975 = ~n9943 ^ ~n9974;
  assign n9976 = n9803 & n9815;
  assign n9977 = n9811 & ~n9814;
  assign n9978 = ~n9976 & ~n9977;
  assign n9979 = n9839 & ~n9842;
  assign n9980 = ~n9835 & ~n9838;
  assign n9981 = ~n9979 & ~n9980;
  assign n9982 = n9900 & ~n9905;
  assign n9983 = ~n9894 & ~n9899;
  assign n9984 = ~n9982 & ~n9983;
  assign n9985 = ~n9981 ^ n9984;
  assign n9986 = n9824 & n9827;
  assign n9987 = n9820 & n9823;
  assign n9988 = ~n9986 & ~n9987;
  assign n9989 = ~n9985 ^ n9988;
  assign n9990 = ~n9978 ^ n9989;
  assign n9991 = n9808 & n9810;
  assign n9992 = n9806 & n9807;
  assign n9993 = ~n9991 & ~n9992;
  assign n9994 = n9875 & ~n9876;
  assign n9995 = ~n9873 & ~n9874;
  assign n9996 = ~n9994 & ~n9995;
  assign n9997 = pi23 & pi60;
  assign n9998 = pi24 & pi59;
  assign n9999 = ~n9997 ^ ~n9998;
  assign n10000 = ~n9996 ^ ~n9999;
  assign n10001 = pi31 & pi52;
  assign n10002 = pi30 & pi53;
  assign n10003 = ~n10001 ^ ~n10002;
  assign n10004 = pi28 & pi55;
  assign n10005 = ~n10003 ^ n10004;
  assign n10006 = ~n10000 ^ n10005;
  assign n10007 = ~n9993 ^ n10006;
  assign n10008 = ~n9990 ^ ~n10007;
  assign n10009 = ~n9975 ^ n10008;
  assign n10010 = ~n9940 ^ n10009;
  assign n10011 = ~n9937 ^ n10010;
  assign n10012 = n9817 & ~n9844;
  assign n10013 = n9800 & n9816;
  assign n10014 = ~n10012 & ~n10013;
  assign n10015 = ~n9848 & n9863;
  assign n10016 = ~n9851 & ~n9862;
  assign n10017 = ~n10015 & ~n10016;
  assign n10018 = n9858 & n9861;
  assign n10019 = n9854 & n9857;
  assign n10020 = ~n10018 & ~n10019;
  assign n10021 = pi32 & pi51;
  assign n10022 = pi26 & pi57;
  assign n10023 = ~n10021 ^ ~n10022;
  assign n10024 = pi25 & pi58;
  assign n10025 = ~n10023 ^ n10024;
  assign n10026 = pi38 & pi45;
  assign n10027 = pi37 & pi46;
  assign n10028 = ~n10026 ^ ~n10027;
  assign n10029 = pi36 & pi47;
  assign n10030 = ~n10028 ^ n10029;
  assign n10031 = ~n10025 ^ ~n10030;
  assign n10032 = pi27 & pi56;
  assign n10033 = pi22 & pi61;
  assign n10034 = ~n10032 ^ ~n10033;
  assign n10035 = pi20 & pi63;
  assign n10036 = ~n10034 ^ n10035;
  assign n10037 = ~n10031 ^ n10036;
  assign n10038 = pi40 & pi43;
  assign n10039 = pi39 & pi44;
  assign n10040 = ~n10038 ^ ~n10039;
  assign n10041 = pi29 & pi54;
  assign n10042 = ~n10040 ^ n10041;
  assign n10043 = pi35 & pi48;
  assign n10044 = pi34 & pi49;
  assign n10045 = ~n10043 ^ ~n10044;
  assign n10046 = pi33 & pi50;
  assign n10047 = ~n10045 ^ n10046;
  assign n10048 = ~n10042 ^ ~n10047;
  assign n10049 = pi21 & pi62;
  assign n10050 = ~pi41 & pi42;
  assign n10051 = ~n10049 ^ ~n10050;
  assign n10052 = ~n10048 ^ ~n10051;
  assign n10053 = ~n10037 ^ ~n10052;
  assign n10054 = ~n10020 ^ ~n10053;
  assign n10055 = ~n10017 ^ n10054;
  assign n10056 = ~n10014 ^ n10055;
  assign n10057 = ~n10011 ^ n10056;
  assign po084 = n9934 ^ ~n10057;
  assign n10059 = ~n9791 & ~n9866;
  assign n10060 = n9788 & ~n10059;
  assign n10061 = n9791 & n9866;
  assign n10062 = n10057 & ~n9920;
  assign n10063 = ~n10061 & ~n10062;
  assign n10064 = ~n10060 & n10063;
  assign n10065 = n10061 & ~n9920;
  assign n10066 = ~n10065 & ~n10057;
  assign n10067 = n9788 & ~n10066;
  assign n10068 = ~n10059 & n10057;
  assign n10069 = ~n10068 & ~n9918;
  assign n10070 = ~n10067 & n10069;
  assign n10071 = ~n10064 & ~n10070;
  assign n10072 = n10011 & ~n10056;
  assign n10073 = ~n9937 & n10010;
  assign n10074 = ~n10072 & ~n10073;
  assign n10075 = ~n9940 & n10009;
  assign n10076 = n9975 & ~n10008;
  assign n10077 = ~n10075 & ~n10076;
  assign n10078 = n9990 & n10007;
  assign n10079 = ~n9978 & n9989;
  assign n10080 = ~n10078 & ~n10079;
  assign n10081 = n9985 & ~n9988;
  assign n10082 = n9981 & ~n9984;
  assign n10083 = ~n10081 & ~n10082;
  assign n10084 = ~n9993 & n10006;
  assign n10085 = n10000 & ~n10005;
  assign n10086 = ~n10084 & ~n10085;
  assign n10087 = ~n10083 ^ ~n10086;
  assign n10088 = n9996 & n9999;
  assign n10089 = n3804 & n9224;
  assign n10090 = ~n10088 & ~n10089;
  assign n10091 = n10034 & ~n10035;
  assign n10092 = ~n10032 & ~n10033;
  assign n10093 = ~n10091 & ~n10092;
  assign n10094 = pi32 & pi52;
  assign n10095 = pi31 & pi53;
  assign n10096 = ~n10094 ^ ~n10095;
  assign n10097 = pi26 & pi58;
  assign n10098 = ~n10096 ^ n10097;
  assign n10099 = ~n10093 ^ n10098;
  assign n10100 = ~n10090 ^ n10099;
  assign n10101 = ~n10087 ^ n10100;
  assign n10102 = ~n10080 ^ ~n10101;
  assign n10103 = n9964 & ~n9967;
  assign n10104 = ~n9960 & ~n9963;
  assign n10105 = ~n10103 & ~n10104;
  assign n10106 = n10023 & ~n10024;
  assign n10107 = ~n10021 & ~n10022;
  assign n10108 = ~n10106 & ~n10107;
  assign n10109 = n10045 & ~n10046;
  assign n10110 = ~n10043 & ~n10044;
  assign n10111 = ~n10109 & ~n10110;
  assign n10112 = ~n10108 ^ ~n10111;
  assign n10113 = n10028 & ~n10029;
  assign n10114 = ~n10026 & ~n10027;
  assign n10115 = ~n10113 & ~n10114;
  assign n10116 = ~n10112 ^ ~n10115;
  assign n10117 = ~n10105 ^ ~n10116;
  assign n10118 = n9953 & n9956;
  assign n10119 = n9949 & n9952;
  assign n10120 = ~n10118 & ~n10119;
  assign n10121 = ~n10117 ^ n10120;
  assign n10122 = pi41 & pi43;
  assign n10123 = pi40 & pi44;
  assign n10124 = ~n10122 ^ ~n10123;
  assign n10125 = pi39 & pi45;
  assign n10126 = ~n10124 ^ n10125;
  assign n10127 = pi38 & pi46;
  assign n10128 = pi29 & pi55;
  assign n10129 = ~n10127 ^ ~n10128;
  assign n10130 = pi28 & pi56;
  assign n10131 = ~n10129 ^ n10130;
  assign n10132 = ~n10126 ^ ~n10131;
  assign n10133 = pi37 & pi47;
  assign n10134 = pi30 & pi54;
  assign n10135 = ~n10133 ^ ~n10134;
  assign n10136 = pi27 & pi57;
  assign n10137 = ~n10135 ^ n10136;
  assign n10138 = ~n10132 ^ n10137;
  assign n10139 = pi36 & pi48;
  assign n10140 = pi35 & pi49;
  assign n10141 = ~n10139 ^ ~n10140;
  assign n10142 = pi34 & pi50;
  assign n10143 = ~n10141 ^ n10142;
  assign n10144 = pi33 & pi51;
  assign n10145 = pi25 & pi59;
  assign n10146 = ~n10144 ^ ~n10145;
  assign n10147 = pi24 & pi60;
  assign n10148 = ~n10146 ^ n10147;
  assign n10149 = ~n10143 ^ ~n10148;
  assign n10150 = pi23 & pi61;
  assign n10151 = pi22 & pi62;
  assign n10152 = ~n10150 ^ ~n10151;
  assign n10153 = pi21 & pi63;
  assign n10154 = ~n10152 ^ n10153;
  assign n10155 = ~n10149 ^ n10154;
  assign n10156 = ~n10138 ^ ~n10155;
  assign n10157 = ~n10121 ^ ~n10156;
  assign n10158 = ~n10102 ^ ~n10157;
  assign n10159 = ~n10077 ^ ~n10158;
  assign n10160 = ~n10014 & n10055;
  assign n10161 = ~n10017 & n10054;
  assign n10162 = ~n10160 & ~n10161;
  assign n10163 = n9943 & n9974;
  assign n10164 = ~n9946 & n9973;
  assign n10165 = ~n10163 & ~n10164;
  assign n10166 = ~n10162 ^ n10165;
  assign n10167 = n10020 & n10053;
  assign n10168 = n10037 & n10052;
  assign n10169 = ~n10167 & ~n10168;
  assign n10170 = n9973 & n9957;
  assign n10171 = ~n9972 & ~n9968;
  assign n10172 = ~n10170 & ~n10171;
  assign n10173 = n10048 & n10051;
  assign n10174 = ~n10042 & ~n10047;
  assign n10175 = ~n10173 & ~n10174;
  assign n10176 = n10040 & ~n10041;
  assign n10177 = ~n10038 & ~n10039;
  assign n10178 = ~n10176 & ~n10177;
  assign n10179 = n10003 & ~n10004;
  assign n10180 = ~n10001 & ~n10002;
  assign n10181 = ~n10179 & ~n10180;
  assign n10182 = ~n10178 ^ ~n10181;
  assign n10183 = ~n10049 & ~pi41;
  assign n10184 = ~n10183 & pi42;
  assign n10185 = ~n10182 ^ n10184;
  assign n10186 = ~n10175 ^ ~n10185;
  assign n10187 = n10031 & ~n10036;
  assign n10188 = ~n10025 & ~n10030;
  assign n10189 = ~n10187 & ~n10188;
  assign n10190 = ~n10186 ^ ~n10189;
  assign n10191 = ~n10172 ^ ~n10190;
  assign n10192 = ~n10169 ^ n10191;
  assign n10193 = ~n10166 ^ n10192;
  assign n10194 = ~n10159 ^ n10193;
  assign n10195 = ~n10074 ^ n10194;
  assign po085 = n10071 ^ n10195;
  assign n10197 = n10074 & n10194;
  assign n10198 = n10071 & ~n10197;
  assign n10199 = ~n10074 & ~n10194;
  assign n10200 = ~n10198 & ~n10199;
  assign n10201 = n10159 & ~n10193;
  assign n10202 = n10077 & n10158;
  assign n10203 = ~n10201 & ~n10202;
  assign n10204 = n10166 & ~n10192;
  assign n10205 = n10162 & ~n10165;
  assign n10206 = ~n10204 & ~n10205;
  assign n10207 = n10102 & n10157;
  assign n10208 = ~n10080 & ~n10101;
  assign n10209 = ~n10207 & ~n10208;
  assign n10210 = n10087 & ~n10100;
  assign n10211 = n10083 & n10086;
  assign n10212 = ~n10210 & ~n10211;
  assign n10213 = ~n10090 & n10099;
  assign n10214 = n10093 & ~n10098;
  assign n10215 = ~n10213 & ~n10214;
  assign n10216 = n10182 & ~n10184;
  assign n10217 = ~n10178 & ~n10181;
  assign n10218 = ~n10216 & ~n10217;
  assign n10219 = n10112 & n10115;
  assign n10220 = n10108 & n10111;
  assign n10221 = ~n10219 & ~n10220;
  assign n10222 = ~n10218 ^ n10221;
  assign n10223 = ~n10215 ^ n10222;
  assign n10224 = ~n10212 ^ ~n10223;
  assign n10225 = n10121 & n10156;
  assign n10226 = n10138 & n10155;
  assign n10227 = ~n10225 & ~n10226;
  assign n10228 = ~n10224 ^ ~n10227;
  assign n10229 = ~n10209 ^ ~n10228;
  assign n10230 = ~n10169 & n10191;
  assign n10231 = ~n10172 & ~n10190;
  assign n10232 = ~n10230 & ~n10231;
  assign n10233 = ~n10229 ^ n10232;
  assign n10234 = n10117 & ~n10120;
  assign n10235 = n10105 & n10116;
  assign n10236 = ~n10234 & ~n10235;
  assign n10237 = n10124 & ~n10125;
  assign n10238 = ~n10122 & ~n10123;
  assign n10239 = ~n10237 & ~n10238;
  assign n10240 = pi24 & pi61;
  assign n10241 = ~n10239 ^ ~n10240;
  assign n10242 = n10129 & ~n10130;
  assign n10243 = ~n10127 & ~n10128;
  assign n10244 = ~n10242 & ~n10243;
  assign n10245 = ~n10241 ^ ~n10244;
  assign n10246 = n10096 & ~n10097;
  assign n10247 = ~n10094 & ~n10095;
  assign n10248 = ~n10246 & ~n10247;
  assign n10249 = pi27 & pi58;
  assign n10250 = pi26 & pi59;
  assign n10251 = ~n10249 ^ ~n10250;
  assign n10252 = pi25 & pi60;
  assign n10253 = ~n10251 ^ n10252;
  assign n10254 = ~n10248 ^ n10253;
  assign n10255 = n10135 & ~n10136;
  assign n10256 = ~n10133 & ~n10134;
  assign n10257 = ~n10255 & ~n10256;
  assign n10258 = ~n10254 ^ n10257;
  assign n10259 = ~n10245 ^ n10258;
  assign n10260 = ~n10236 ^ n10259;
  assign n10261 = n10149 & ~n10154;
  assign n10262 = ~n10143 & ~n10148;
  assign n10263 = ~n10261 & ~n10262;
  assign n10264 = n10132 & ~n10137;
  assign n10265 = ~n10126 & ~n10131;
  assign n10266 = ~n10264 & ~n10265;
  assign n10267 = ~n10263 ^ ~n10266;
  assign n10268 = n10146 & ~n10147;
  assign n10269 = ~n10144 & ~n10145;
  assign n10270 = ~n10268 & ~n10269;
  assign n10271 = n10152 & ~n10153;
  assign n10272 = ~n10150 & ~n10151;
  assign n10273 = ~n10271 & ~n10272;
  assign n10274 = ~n10270 ^ ~n10273;
  assign n10275 = n10141 & ~n10142;
  assign n10276 = ~n10139 & ~n10140;
  assign n10277 = ~n10275 & ~n10276;
  assign n10278 = ~n10274 ^ ~n10277;
  assign n10279 = ~n10267 ^ n10278;
  assign n10280 = ~n10260 ^ n10279;
  assign n10281 = n10186 & n10189;
  assign n10282 = n10175 & n10185;
  assign n10283 = ~n10281 & ~n10282;
  assign n10284 = pi31 & pi54;
  assign n10285 = ~n5612 ^ ~n10284;
  assign n10286 = pi30 & pi55;
  assign n10287 = ~n10285 ^ n10286;
  assign n10288 = pi38 & pi47;
  assign n10289 = pi37 & pi48;
  assign n10290 = ~n10288 ^ ~n10289;
  assign n10291 = pi36 & pi49;
  assign n10292 = ~n10290 ^ n10291;
  assign n10293 = ~n10287 ^ ~n10292;
  assign n10294 = pi23 & pi62;
  assign n10295 = ~pi42 & pi43;
  assign n10296 = ~n10294 ^ ~n10295;
  assign n10297 = ~n10293 ^ ~n10296;
  assign n10298 = ~n10283 ^ ~n10297;
  assign n10299 = pi35 & pi50;
  assign n10300 = pi28 & pi57;
  assign n10301 = ~n10299 ^ ~n10300;
  assign n10302 = pi22 & pi63;
  assign n10303 = ~n10301 ^ n10302;
  assign n10304 = pi34 & pi51;
  assign n10305 = pi33 & pi52;
  assign n10306 = ~n10304 ^ ~n10305;
  assign n10307 = pi32 & pi53;
  assign n10308 = ~n10306 ^ n10307;
  assign n10309 = ~n10303 ^ ~n10308;
  assign n10310 = pi41 & pi44;
  assign n10311 = pi40 & pi45;
  assign n10312 = ~n10310 ^ ~n10311;
  assign n10313 = pi39 & pi46;
  assign n10314 = ~n10312 ^ n10313;
  assign n10315 = ~n10309 ^ n10314;
  assign n10316 = ~n10298 ^ ~n10315;
  assign n10317 = ~n10280 ^ ~n10316;
  assign n10318 = ~n10233 ^ ~n10317;
  assign n10319 = ~n10206 ^ n10318;
  assign n10320 = ~n10203 ^ n10319;
  assign po086 = n10200 ^ ~n10320;
  assign n10322 = n10203 & ~n10206;
  assign n10323 = ~n10322 & n10317;
  assign n10324 = ~n10203 & n10206;
  assign n10325 = ~n10323 & ~n10324;
  assign n10326 = n10322 & ~n10317;
  assign n10327 = ~n10326 & n10233;
  assign n10328 = n10325 & ~n10327;
  assign n10329 = ~n10200 & n10328;
  assign n10330 = n10324 & n10317;
  assign n10331 = ~n10330 & ~n10326;
  assign n10332 = ~n10331 & ~n10318;
  assign n10333 = ~n10329 & ~n10332;
  assign n10334 = ~n10330 & ~n10233;
  assign n10335 = ~n10325 & ~n10334;
  assign n10336 = n10200 & n10335;
  assign n10337 = n10333 & ~n10336;
  assign n10338 = n10229 & ~n10232;
  assign n10339 = ~n10209 & ~n10228;
  assign n10340 = ~n10338 & ~n10339;
  assign n10341 = ~n10215 & n10222;
  assign n10342 = n10218 & ~n10221;
  assign n10343 = ~n10341 & ~n10342;
  assign n10344 = n10301 & ~n10302;
  assign n10345 = ~n10299 & ~n10300;
  assign n10346 = ~n10344 & ~n10345;
  assign n10347 = n10251 & ~n10252;
  assign n10348 = ~n10249 & ~n10250;
  assign n10349 = ~n10347 & ~n10348;
  assign n10350 = ~n10346 ^ ~n10349;
  assign n10351 = n10306 & ~n10307;
  assign n10352 = ~n10304 & ~n10305;
  assign n10353 = ~n10351 & ~n10352;
  assign n10354 = ~n10350 ^ ~n10353;
  assign n10355 = ~n10343 ^ n10354;
  assign n10356 = n10290 & ~n10291;
  assign n10357 = ~n10288 & ~n10289;
  assign n10358 = ~n10356 & ~n10357;
  assign n10359 = n10312 & ~n10313;
  assign n10360 = ~n10310 & ~n10311;
  assign n10361 = ~n10359 & ~n10360;
  assign n10362 = ~n10358 ^ ~n10361;
  assign n10363 = n10285 & ~n10286;
  assign n10364 = ~n5612 & ~n10284;
  assign n10365 = ~n10363 & ~n10364;
  assign n10366 = ~n10362 ^ n10365;
  assign n10367 = ~n10355 ^ n10366;
  assign n10368 = n10267 & ~n10278;
  assign n10369 = n10263 & n10266;
  assign n10370 = ~n10368 & ~n10369;
  assign n10371 = pi38 & pi48;
  assign n10372 = pi31 & pi55;
  assign n10373 = ~n10371 ^ ~n10372;
  assign n10374 = ~n10373 ^ n5565;
  assign n10375 = pi37 & pi49;
  assign n10376 = pi36 & pi50;
  assign n10377 = ~n10375 ^ ~n10376;
  assign n10378 = pi23 & pi63;
  assign n10379 = ~n10377 ^ n10378;
  assign n10380 = ~n10374 ^ ~n10379;
  assign n10381 = pi35 & pi51;
  assign n10382 = pi34 & pi52;
  assign n10383 = ~n10381 ^ ~n10382;
  assign n10384 = pi33 & pi53;
  assign n10385 = ~n10383 ^ n10384;
  assign n10386 = ~n10380 ^ n10385;
  assign n10387 = pi40 & pi46;
  assign n10388 = pi39 & pi47;
  assign n10389 = ~n10387 ^ ~n10388;
  assign n10390 = pi30 & pi56;
  assign n10391 = ~n10389 ^ n10390;
  assign n10392 = pi28 & pi58;
  assign n10393 = pi27 & pi59;
  assign n10394 = ~n10392 ^ ~n10393;
  assign n10395 = pi26 & pi60;
  assign n10396 = ~n10394 ^ n10395;
  assign n10397 = ~n10391 ^ n10396;
  assign n10398 = pi42 & pi44;
  assign n10399 = pi41 & pi45;
  assign n10400 = ~n10398 ^ ~n10399;
  assign n10401 = pi32 & pi54;
  assign n10402 = ~n10400 ^ n10401;
  assign n10403 = ~n10397 ^ ~n10402;
  assign n10404 = ~n10386 ^ ~n10403;
  assign n10405 = ~n10370 ^ ~n10404;
  assign n10406 = n10254 & ~n10257;
  assign n10407 = ~n10248 & n10253;
  assign n10408 = ~n10406 & ~n10407;
  assign n10409 = n10293 & n10296;
  assign n10410 = ~n10287 & ~n10292;
  assign n10411 = ~n10409 & ~n10410;
  assign n10412 = ~n10408 ^ n10411;
  assign n10413 = n10309 & ~n10314;
  assign n10414 = ~n10303 & ~n10308;
  assign n10415 = ~n10413 & ~n10414;
  assign n10416 = ~n10412 ^ n10415;
  assign n10417 = ~n10405 ^ ~n10416;
  assign n10418 = ~n10367 ^ n10417;
  assign n10419 = ~n10340 ^ ~n10418;
  assign n10420 = n10224 & n10227;
  assign n10421 = ~n10212 & ~n10223;
  assign n10422 = ~n10420 & ~n10421;
  assign n10423 = ~n10236 & n10259;
  assign n10424 = n10245 & ~n10258;
  assign n10425 = ~n10423 & ~n10424;
  assign n10426 = n10298 & n10315;
  assign n10427 = n10283 & n10297;
  assign n10428 = ~n10426 & ~n10427;
  assign n10429 = ~n10425 ^ ~n10428;
  assign n10430 = n10274 & n10277;
  assign n10431 = n10270 & n10273;
  assign n10432 = ~n10430 & ~n10431;
  assign n10433 = ~n10294 & ~pi42;
  assign n10434 = ~n10433 & pi43;
  assign n10435 = pi25 & pi61;
  assign n10436 = pi24 & pi62;
  assign n10437 = ~n10435 ^ ~n10436;
  assign n10438 = ~n10434 ^ n10437;
  assign n10439 = ~n10432 ^ ~n10438;
  assign n10440 = n10241 & n10244;
  assign n10441 = n10239 & n10240;
  assign n10442 = ~n10440 & ~n10441;
  assign n10443 = ~n10439 ^ n10442;
  assign n10444 = ~n10429 ^ ~n10443;
  assign n10445 = ~n10422 ^ ~n10444;
  assign n10446 = n10280 & n10316;
  assign n10447 = n10260 & ~n10279;
  assign n10448 = ~n10446 & ~n10447;
  assign n10449 = ~n10445 ^ ~n10448;
  assign n10450 = ~n10419 ^ n10449;
  assign po087 = n10337 ^ n10450;
  assign n10452 = ~n10199 & ~n10322;
  assign n10453 = ~n10198 & n10452;
  assign n10454 = ~n10453 & ~n10324;
  assign n10455 = n10233 & n10317;
  assign n10456 = ~n10450 & ~n10455;
  assign n10457 = ~n10454 & ~n10456;
  assign n10458 = ~n10324 & ~n10450;
  assign n10459 = ~n10233 & ~n10317;
  assign n10460 = ~n10458 & ~n10459;
  assign n10461 = n10200 & n10460;
  assign n10462 = ~n10327 & ~n10323;
  assign n10463 = ~n10462 & n10450;
  assign n10464 = ~n10461 & ~n10463;
  assign n10465 = ~n10457 & n10464;
  assign n10466 = n10419 & ~n10449;
  assign n10467 = ~n10340 & ~n10418;
  assign n10468 = ~n10466 & ~n10467;
  assign n10469 = n10445 & n10448;
  assign n10470 = ~n10422 & ~n10444;
  assign n10471 = ~n10469 & ~n10470;
  assign n10472 = n10355 & ~n10366;
  assign n10473 = ~n10343 & n10354;
  assign n10474 = ~n10472 & ~n10473;
  assign n10475 = n10412 & ~n10415;
  assign n10476 = n10408 & ~n10411;
  assign n10477 = ~n10475 & ~n10476;
  assign n10478 = ~n10474 ^ ~n10477;
  assign n10479 = n10439 & ~n10442;
  assign n10480 = ~n10432 & ~n10438;
  assign n10481 = ~n10479 & ~n10480;
  assign n10482 = n10394 & ~n10395;
  assign n10483 = ~n10392 & ~n10393;
  assign n10484 = ~n10482 & ~n10483;
  assign n10485 = n10377 & ~n10378;
  assign n10486 = ~n10375 & ~n10376;
  assign n10487 = ~n10485 & ~n10486;
  assign n10488 = ~n10484 ^ ~n10487;
  assign n10489 = n10383 & ~n10384;
  assign n10490 = ~n10381 & ~n10382;
  assign n10491 = ~n10489 & ~n10490;
  assign n10492 = ~n10488 ^ n10491;
  assign n10493 = ~n10481 ^ ~n10492;
  assign n10494 = n10373 & ~n5565;
  assign n10495 = ~n10371 & ~n10372;
  assign n10496 = ~n10494 & ~n10495;
  assign n10497 = n10389 & ~n10390;
  assign n10498 = ~n10387 & ~n10388;
  assign n10499 = ~n10497 & ~n10498;
  assign n10500 = ~n10496 ^ ~n10499;
  assign n10501 = n10400 & ~n10401;
  assign n10502 = ~n10398 & ~n10399;
  assign n10503 = ~n10501 & ~n10502;
  assign n10504 = ~n10500 ^ ~n10503;
  assign n10505 = ~n10493 ^ n10504;
  assign n10506 = ~n10478 ^ n10505;
  assign n10507 = ~n10367 & n10417;
  assign n10508 = ~n10405 & ~n10416;
  assign n10509 = ~n10507 & ~n10508;
  assign n10510 = ~n10506 ^ ~n10509;
  assign n10511 = n10350 & n10353;
  assign n10512 = n10346 & n10349;
  assign n10513 = ~n10511 & ~n10512;
  assign n10514 = pi40 & pi47;
  assign n10515 = pi33 & pi54;
  assign n10516 = ~n10514 ^ ~n10515;
  assign n10517 = pi31 & pi56;
  assign n10518 = ~n10516 ^ n10517;
  assign n10519 = pi25 & pi62;
  assign n10520 = ~pi43 & pi44;
  assign n10521 = ~n10519 ^ ~n10520;
  assign n10522 = ~n10518 ^ n10521;
  assign n10523 = ~n10513 ^ n10522;
  assign n10524 = pi42 & pi45;
  assign n10525 = pi41 & pi46;
  assign n10526 = ~n10524 ^ ~n10525;
  assign n10527 = pi32 & pi55;
  assign n10528 = ~n10526 ^ n10527;
  assign n10529 = pi27 & pi60;
  assign n10530 = pi26 & pi61;
  assign n10531 = ~n10529 ^ ~n10530;
  assign n10532 = pi24 & pi63;
  assign n10533 = ~n10531 ^ n10532;
  assign n10534 = ~n10528 ^ ~n10533;
  assign n10535 = pi39 & pi48;
  assign n10536 = pi38 & pi49;
  assign n10537 = ~n10535 ^ ~n10536;
  assign n10538 = pi37 & pi50;
  assign n10539 = ~n10537 ^ n10538;
  assign n10540 = ~n10534 ^ n10539;
  assign n10541 = ~n10523 ^ ~n10540;
  assign n10542 = ~n10435 & ~pi24;
  assign n10543 = pi43 & pi62;
  assign n10544 = ~n10542 & n10543;
  assign n10545 = n10544 & ~n7410;
  assign n10546 = n10435 & n10436;
  assign n10547 = pi42 & pi61;
  assign n10548 = n7511 & n10547;
  assign n10549 = ~n10546 & ~n10548;
  assign n10550 = ~n10545 & n10549;
  assign n10551 = pi36 & pi51;
  assign n10552 = pi35 & pi52;
  assign n10553 = ~n10551 ^ ~n10552;
  assign n10554 = pi29 & pi58;
  assign n10555 = ~n10553 ^ n10554;
  assign n10556 = pi34 & pi53;
  assign n10557 = pi30 & pi57;
  assign n10558 = ~n10556 ^ ~n10557;
  assign n10559 = pi28 & pi59;
  assign n10560 = ~n10558 ^ n10559;
  assign n10561 = ~n10555 ^ ~n10560;
  assign n10562 = ~n10550 ^ n10561;
  assign n10563 = ~n10541 ^ n10562;
  assign n10564 = ~n10510 ^ ~n10563;
  assign n10565 = n10429 & n10443;
  assign n10566 = ~n10425 & ~n10428;
  assign n10567 = ~n10565 & ~n10566;
  assign n10568 = ~n10391 & ~n10396;
  assign n10569 = ~n10568 & n10402;
  assign n10570 = n10391 & n10396;
  assign n10571 = ~n10569 & ~n10570;
  assign n10572 = n10571 & n10404;
  assign n10573 = n10370 & n10572;
  assign n10574 = n10568 & ~n10402;
  assign n10575 = n10386 & n10574;
  assign n10576 = ~n10573 & ~n10575;
  assign n10577 = n10570 & n10402;
  assign n10578 = ~n10370 & n10577;
  assign n10579 = n10576 & ~n10578;
  assign n10580 = ~n10571 & ~n10386;
  assign n10581 = n10580 & n10405;
  assign n10582 = n10579 & ~n10581;
  assign n10583 = n10362 & ~n10365;
  assign n10584 = ~n10358 & ~n10361;
  assign n10585 = ~n10583 & ~n10584;
  assign n10586 = n10380 & ~n10385;
  assign n10587 = ~n10374 & ~n10379;
  assign n10588 = ~n10586 & ~n10587;
  assign n10589 = ~n10585 ^ n10588;
  assign n10590 = ~n10582 ^ ~n10589;
  assign n10591 = ~n10567 ^ ~n10590;
  assign n10592 = ~n10564 ^ ~n10591;
  assign n10593 = ~n10471 ^ n10592;
  assign n10594 = ~n10468 ^ ~n10593;
  assign po088 = n10465 ^ ~n10594;
  assign n10596 = n10468 & n10593;
  assign n10597 = ~n10465 & ~n10596;
  assign n10598 = ~n10468 & ~n10593;
  assign n10599 = ~n10597 & ~n10598;
  assign n10600 = ~n10593 & n10591;
  assign n10601 = ~n10471 & n10564;
  assign n10602 = ~n10600 & ~n10601;
  assign n10603 = n10478 & ~n10505;
  assign n10604 = ~n10474 & ~n10477;
  assign n10605 = ~n10603 & ~n10604;
  assign n10606 = n10541 & ~n10562;
  assign n10607 = ~n10523 & ~n10540;
  assign n10608 = ~n10606 & ~n10607;
  assign n10609 = ~n10605 ^ n10608;
  assign n10610 = ~n10550 & n10561;
  assign n10611 = ~n10555 & ~n10560;
  assign n10612 = ~n10610 & ~n10611;
  assign n10613 = n10488 & ~n10491;
  assign n10614 = ~n10484 & ~n10487;
  assign n10615 = ~n10613 & ~n10614;
  assign n10616 = ~n10612 ^ n10615;
  assign n10617 = n10534 & ~n10539;
  assign n10618 = ~n10528 & ~n10533;
  assign n10619 = ~n10617 & ~n10618;
  assign n10620 = ~n10616 ^ ~n10619;
  assign n10621 = ~n10609 ^ ~n10620;
  assign n10622 = n10510 & n10563;
  assign n10623 = ~n10506 & ~n10509;
  assign n10624 = ~n10622 & ~n10623;
  assign n10625 = ~n10621 ^ n10624;
  assign n10626 = n10567 & n10590;
  assign n10627 = n10589 & ~n10571;
  assign n10628 = n10576 & ~n10627;
  assign n10629 = ~n10590 & n10628;
  assign n10630 = ~n10626 & ~n10629;
  assign n10631 = n10500 & n10503;
  assign n10632 = n10496 & n10499;
  assign n10633 = ~n10631 & ~n10632;
  assign n10634 = pi40 & pi48;
  assign n10635 = pi32 & pi56;
  assign n10636 = ~n10634 ^ ~n10635;
  assign n10637 = pi30 & pi58;
  assign n10638 = ~n10636 ^ n10637;
  assign n10639 = pi39 & pi49;
  assign n10640 = pi38 & pi50;
  assign n10641 = ~n10639 ^ ~n10640;
  assign n10642 = ~n10641 ^ n6130;
  assign n10643 = ~n10638 ^ ~n10642;
  assign n10644 = ~n10633 ^ n10643;
  assign n10645 = ~n10519 & ~pi43;
  assign n10646 = ~n10645 & pi44;
  assign n10647 = pi25 & pi63;
  assign n10648 = ~n10646 & ~n10647;
  assign n10649 = pi62 & pi63;
  assign n10650 = pi43 & pi63;
  assign n10651 = ~n10649 & ~n10650;
  assign n10652 = ~n10651 & n7758;
  assign n10653 = ~n10648 & ~n10652;
  assign n10654 = n10526 & ~n10527;
  assign n10655 = ~n10524 & ~n10525;
  assign n10656 = ~n10654 & ~n10655;
  assign n10657 = ~n10653 ^ ~n10656;
  assign n10658 = ~n10644 ^ ~n10657;
  assign n10659 = pi42 & pi46;
  assign n10660 = pi41 & pi47;
  assign n10661 = ~n10659 ^ ~n10660;
  assign n10662 = pi31 & pi57;
  assign n10663 = ~n10661 ^ n10662;
  assign n10664 = pi28 & pi60;
  assign n10665 = pi27 & pi61;
  assign n10666 = ~n10664 ^ ~n10665;
  assign n10667 = pi26 & pi62;
  assign n10668 = ~n10666 ^ n10667;
  assign n10669 = ~n10663 ^ ~n10668;
  assign n10670 = pi37 & pi51;
  assign n10671 = pi36 & pi52;
  assign n10672 = ~n10670 ^ ~n10671;
  assign n10673 = pi35 & pi53;
  assign n10674 = ~n10672 ^ n10673;
  assign n10675 = ~n10669 ^ n10674;
  assign n10676 = ~n10658 ^ n10675;
  assign n10677 = ~n10630 ^ n10676;
  assign n10678 = n10493 & ~n10504;
  assign n10679 = n10481 & n10492;
  assign n10680 = ~n10678 & ~n10679;
  assign n10681 = ~n10585 & n10588;
  assign n10682 = ~n10627 & ~n10681;
  assign n10683 = ~n10680 ^ ~n10682;
  assign n10684 = ~n10513 & n10522;
  assign n10685 = ~n10518 & n10521;
  assign n10686 = ~n10684 & ~n10685;
  assign n10687 = n10516 & ~n10517;
  assign n10688 = ~n10514 & ~n10515;
  assign n10689 = ~n10687 & ~n10688;
  assign n10690 = pi43 & pi45;
  assign n10691 = pi34 & pi54;
  assign n10692 = ~n10690 ^ ~n10691;
  assign n10693 = pi33 & pi55;
  assign n10694 = ~n10692 ^ n10693;
  assign n10695 = ~n10689 ^ n10694;
  assign n10696 = n10553 & ~n10554;
  assign n10697 = ~n10551 & ~n10552;
  assign n10698 = ~n10696 & ~n10697;
  assign n10699 = ~n10695 ^ n10698;
  assign n10700 = ~n10686 ^ ~n10699;
  assign n10701 = n10531 & ~n10532;
  assign n10702 = ~n10529 & ~n10530;
  assign n10703 = ~n10701 & ~n10702;
  assign n10704 = n10537 & ~n10538;
  assign n10705 = ~n10535 & ~n10536;
  assign n10706 = ~n10704 & ~n10705;
  assign n10707 = ~n10703 ^ ~n10706;
  assign n10708 = n10558 & ~n10559;
  assign n10709 = ~n10556 & ~n10557;
  assign n10710 = ~n10708 & ~n10709;
  assign n10711 = ~n10707 ^ ~n10710;
  assign n10712 = ~n10700 ^ n10711;
  assign n10713 = ~n10683 ^ n10712;
  assign n10714 = ~n10677 ^ ~n10713;
  assign n10715 = ~n10625 ^ n10714;
  assign n10716 = ~n10602 ^ n10715;
  assign po089 = n10599 ^ ~n10716;
  assign n10718 = n10602 & ~n10715;
  assign n10719 = ~n10598 & ~n10718;
  assign n10720 = ~n10597 & n10719;
  assign n10721 = ~n10602 & n10715;
  assign n10722 = ~n10720 & ~n10721;
  assign n10723 = n10609 & n10620;
  assign n10724 = n10605 & ~n10608;
  assign n10725 = ~n10723 & ~n10724;
  assign n10726 = n10700 & ~n10711;
  assign n10727 = n10686 & n10699;
  assign n10728 = ~n10726 & ~n10727;
  assign n10729 = n10616 & n10619;
  assign n10730 = n10612 & ~n10615;
  assign n10731 = ~n10729 & ~n10730;
  assign n10732 = n10695 & ~n10698;
  assign n10733 = ~n10689 & n10694;
  assign n10734 = ~n10732 & ~n10733;
  assign n10735 = ~n10648 & n10656;
  assign n10736 = ~n10735 & ~n10652;
  assign n10737 = ~n10734 ^ n10736;
  assign n10738 = n10707 & n10710;
  assign n10739 = n10703 & n10706;
  assign n10740 = ~n10738 & ~n10739;
  assign n10741 = ~n10737 ^ ~n10740;
  assign n10742 = ~n10731 ^ n10741;
  assign n10743 = ~n10728 ^ ~n10742;
  assign n10744 = ~n10725 ^ ~n10743;
  assign n10745 = n10692 & ~n10693;
  assign n10746 = ~n10690 & ~n10691;
  assign n10747 = ~n10745 & ~n10746;
  assign n10748 = pi28 & pi61;
  assign n10749 = pi29 & pi60;
  assign n10750 = ~n10748 ^ ~n10749;
  assign n10751 = ~n10747 ^ ~n10750;
  assign n10752 = pi43 & pi46;
  assign n10753 = pi42 & pi47;
  assign n10754 = ~n10752 ^ ~n10753;
  assign n10755 = pi34 & pi55;
  assign n10756 = ~n10754 ^ n10755;
  assign n10757 = ~n10751 ^ n10756;
  assign n10758 = pi27 & pi62;
  assign n10759 = ~pi44 & pi45;
  assign n10760 = ~n10758 ^ ~n10759;
  assign n10761 = ~n10757 ^ ~n10760;
  assign n10762 = pi32 & pi57;
  assign n10763 = pi31 & pi58;
  assign n10764 = ~n10762 ^ ~n10763;
  assign n10765 = pi30 & pi59;
  assign n10766 = ~n10764 ^ n10765;
  assign n10767 = pi38 & pi51;
  assign n10768 = pi37 & pi52;
  assign n10769 = ~n10767 ^ ~n10768;
  assign n10770 = pi36 & pi53;
  assign n10771 = ~n10769 ^ n10770;
  assign n10772 = ~n10766 ^ ~n10771;
  assign n10773 = pi41 & pi48;
  assign n10774 = pi35 & pi54;
  assign n10775 = ~n10773 ^ ~n10774;
  assign n10776 = pi33 & pi56;
  assign n10777 = ~n10775 ^ n10776;
  assign n10778 = ~n10772 ^ n10777;
  assign n10779 = ~n10761 ^ ~n10778;
  assign n10780 = n10636 & ~n10637;
  assign n10781 = ~n10634 & ~n10635;
  assign n10782 = ~n10780 & ~n10781;
  assign n10783 = n10672 & ~n10673;
  assign n10784 = ~n10670 & ~n10671;
  assign n10785 = ~n10783 & ~n10784;
  assign n10786 = ~n10782 ^ ~n10785;
  assign n10787 = n10666 & ~n10667;
  assign n10788 = ~n10664 & ~n10665;
  assign n10789 = ~n10787 & ~n10788;
  assign n10790 = ~n10786 ^ ~n10789;
  assign n10791 = ~n10779 ^ n10790;
  assign n10792 = ~n10744 ^ ~n10791;
  assign n10793 = n10683 & ~n10712;
  assign n10794 = n10680 & n10682;
  assign n10795 = ~n10793 & ~n10794;
  assign n10796 = n10658 & ~n10675;
  assign n10797 = ~n10644 & ~n10657;
  assign n10798 = ~n10796 & ~n10797;
  assign n10799 = ~n10795 ^ n10798;
  assign n10800 = ~n10633 & n10643;
  assign n10801 = ~n10638 & ~n10642;
  assign n10802 = ~n10800 & ~n10801;
  assign n10803 = n10641 & ~n6130;
  assign n10804 = ~n10639 & ~n10640;
  assign n10805 = ~n10803 & ~n10804;
  assign n10806 = pi40 & pi49;
  assign n10807 = pi39 & pi50;
  assign n10808 = ~n10806 ^ ~n10807;
  assign n10809 = pi26 & pi63;
  assign n10810 = ~n10808 ^ n10809;
  assign n10811 = ~n10805 ^ n10810;
  assign n10812 = n10661 & ~n10662;
  assign n10813 = ~n10659 & ~n10660;
  assign n10814 = ~n10812 & ~n10813;
  assign n10815 = ~n10811 ^ ~n10814;
  assign n10816 = ~n10802 ^ n10815;
  assign n10817 = n10669 & ~n10674;
  assign n10818 = ~n10663 & ~n10668;
  assign n10819 = ~n10817 & ~n10818;
  assign n10820 = ~n10816 ^ n10819;
  assign n10821 = ~n10799 ^ n10820;
  assign n10822 = ~n10792 ^ ~n10821;
  assign n10823 = n10677 & n10713;
  assign n10824 = n10630 & ~n10676;
  assign n10825 = ~n10823 & ~n10824;
  assign n10826 = ~n10822 ^ ~n10825;
  assign n10827 = n10625 & ~n10714;
  assign n10828 = n10621 & ~n10624;
  assign n10829 = ~n10827 & ~n10828;
  assign n10830 = ~n10826 ^ n10829;
  assign po090 = n10722 ^ n10830;
  assign n10832 = ~n10826 & n10829;
  assign n10833 = ~n10722 & ~n10832;
  assign n10834 = n10826 & ~n10829;
  assign n10835 = ~n10833 & ~n10834;
  assign n10836 = n10822 & n10825;
  assign n10837 = n10792 & n10821;
  assign n10838 = ~n10836 & ~n10837;
  assign n10839 = n10744 & n10791;
  assign n10840 = ~n10725 & ~n10743;
  assign n10841 = ~n10839 & ~n10840;
  assign n10842 = n10799 & ~n10820;
  assign n10843 = n10795 & ~n10798;
  assign n10844 = ~n10842 & ~n10843;
  assign n10845 = n10816 & ~n10819;
  assign n10846 = ~n10802 & n10815;
  assign n10847 = ~n10845 & ~n10846;
  assign n10848 = n10747 & n10750;
  assign n10849 = n5371 & n7772;
  assign n10850 = ~n10848 & ~n10849;
  assign n10851 = pi32 & pi58;
  assign n10852 = ~n6365 ^ ~n10851;
  assign n10853 = pi30 & pi60;
  assign n10854 = ~n10852 ^ n10853;
  assign n10855 = pi29 & pi61;
  assign n10856 = pi28 & pi62;
  assign n10857 = ~n10855 ^ ~n10856;
  assign n10858 = pi27 & pi63;
  assign n10859 = ~n10857 ^ n10858;
  assign n10860 = ~n10854 ^ ~n10859;
  assign n10861 = ~n10850 ^ n10860;
  assign n10862 = ~n10847 ^ n10861;
  assign n10863 = n10811 & n10814;
  assign n10864 = n10805 & ~n10810;
  assign n10865 = ~n10863 & ~n10864;
  assign n10866 = pi41 & pi49;
  assign n10867 = pi40 & pi50;
  assign n10868 = ~n10866 ^ ~n10867;
  assign n10869 = pi39 & pi51;
  assign n10870 = ~n10868 ^ n10869;
  assign n10871 = ~n10865 ^ ~n10870;
  assign n10872 = n10786 & n10789;
  assign n10873 = n10782 & n10785;
  assign n10874 = ~n10872 & ~n10873;
  assign n10875 = ~n10871 ^ ~n10874;
  assign n10876 = ~n10862 ^ n10875;
  assign n10877 = ~n10844 ^ ~n10876;
  assign n10878 = n10737 & n10740;
  assign n10879 = ~n10734 & n10736;
  assign n10880 = ~n10878 & ~n10879;
  assign n10881 = n10764 & ~n10765;
  assign n10882 = ~n10762 & ~n10763;
  assign n10883 = ~n10881 & ~n10882;
  assign n10884 = n10808 & ~n10809;
  assign n10885 = ~n10806 & ~n10807;
  assign n10886 = ~n10884 & ~n10885;
  assign n10887 = ~n10883 ^ ~n10886;
  assign n10888 = n10769 & ~n10770;
  assign n10889 = ~n10767 & ~n10768;
  assign n10890 = ~n10888 & ~n10889;
  assign n10891 = ~n10887 ^ n10890;
  assign n10892 = pi35 & pi55;
  assign n10893 = pi34 & pi56;
  assign n10894 = ~n10892 ^ ~n10893;
  assign n10895 = pi33 & pi57;
  assign n10896 = ~n10894 ^ n10895;
  assign n10897 = pi38 & pi52;
  assign n10898 = pi37 & pi53;
  assign n10899 = ~n10897 ^ ~n10898;
  assign n10900 = pi36 & pi54;
  assign n10901 = ~n10899 ^ n10900;
  assign n10902 = ~n10896 ^ ~n10901;
  assign n10903 = pi44 & pi46;
  assign n10904 = pi43 & pi47;
  assign n10905 = ~n10903 ^ ~n10904;
  assign n10906 = pi42 & pi48;
  assign n10907 = ~n10905 ^ n10906;
  assign n10908 = ~n10902 ^ n10907;
  assign n10909 = ~n10891 ^ n10908;
  assign n10910 = ~n10880 ^ n10909;
  assign n10911 = ~n10877 ^ ~n10910;
  assign n10912 = ~n10841 ^ n10911;
  assign n10913 = ~n10743 & ~n10741;
  assign n10914 = n10728 & n10731;
  assign n10915 = ~n10913 & ~n10914;
  assign n10916 = n10779 & ~n10790;
  assign n10917 = ~n10761 & ~n10778;
  assign n10918 = ~n10916 & ~n10917;
  assign n10919 = n10757 & n10760;
  assign n10920 = n10751 & ~n10756;
  assign n10921 = ~n10919 & ~n10920;
  assign n10922 = n10754 & ~n10755;
  assign n10923 = ~n10752 & ~n10753;
  assign n10924 = ~n10922 & ~n10923;
  assign n10925 = n10775 & ~n10776;
  assign n10926 = ~n10773 & ~n10774;
  assign n10927 = ~n10925 & ~n10926;
  assign n10928 = ~n10924 ^ ~n10927;
  assign n10929 = ~n10758 & ~pi44;
  assign n10930 = ~n10929 & pi45;
  assign n10931 = ~n10928 ^ n10930;
  assign n10932 = ~n10921 ^ ~n10931;
  assign n10933 = n10772 & ~n10777;
  assign n10934 = ~n10766 & ~n10771;
  assign n10935 = ~n10933 & ~n10934;
  assign n10936 = ~n10932 ^ ~n10935;
  assign n10937 = ~n10918 ^ n10936;
  assign n10938 = ~n10915 ^ ~n10937;
  assign n10939 = ~n10912 ^ n10938;
  assign n10940 = ~n10838 ^ ~n10939;
  assign po091 = n10835 ^ n10940;
  assign n10942 = n10838 & n10939;
  assign n10943 = ~n10835 & ~n10942;
  assign n10944 = ~n10838 & ~n10939;
  assign n10945 = ~n10943 & ~n10944;
  assign n10946 = n10912 & ~n10938;
  assign n10947 = n10841 & ~n10911;
  assign n10948 = ~n10946 & ~n10947;
  assign n10949 = n10877 & n10910;
  assign n10950 = ~n10844 & ~n10876;
  assign n10951 = ~n10949 & ~n10950;
  assign n10952 = n10915 & n10937;
  assign n10953 = ~n10918 & n10936;
  assign n10954 = ~n10952 & ~n10953;
  assign n10955 = n10871 & n10874;
  assign n10956 = n10865 & n10870;
  assign n10957 = ~n10955 & ~n10956;
  assign n10958 = pi44 & pi47;
  assign n10959 = pi43 & pi48;
  assign n10960 = ~n10958 ^ ~n10959;
  assign n10961 = pi35 & pi56;
  assign n10962 = ~n10960 ^ n10961;
  assign n10963 = pi41 & pi50;
  assign n10964 = pi40 & pi51;
  assign n10965 = ~n10963 ^ ~n10964;
  assign n10966 = pi28 & pi63;
  assign n10967 = ~n10965 ^ n10966;
  assign n10968 = ~n10962 ^ ~n10967;
  assign n10969 = pi29 & pi62;
  assign n10970 = ~pi45 & pi46;
  assign n10971 = ~n10969 ^ ~n10970;
  assign n10972 = ~n10968 ^ ~n10971;
  assign n10973 = ~n10957 ^ ~n10972;
  assign n10974 = n10852 & ~n10853;
  assign n10975 = ~n6365 & ~n10851;
  assign n10976 = ~n10974 & ~n10975;
  assign n10977 = n10899 & ~n10900;
  assign n10978 = ~n10897 & ~n10898;
  assign n10979 = ~n10977 & ~n10978;
  assign n10980 = ~n10976 ^ ~n10979;
  assign n10981 = n10857 & ~n10858;
  assign n10982 = ~n10855 & ~n10856;
  assign n10983 = ~n10981 & ~n10982;
  assign n10984 = ~n10980 ^ ~n10983;
  assign n10985 = ~n10973 ^ n10984;
  assign n10986 = ~n10954 ^ n10985;
  assign n10987 = n10932 & n10935;
  assign n10988 = n10921 & n10931;
  assign n10989 = ~n10987 & ~n10988;
  assign n10990 = n10928 & ~n10930;
  assign n10991 = ~n10924 & ~n10927;
  assign n10992 = ~n10990 & ~n10991;
  assign n10993 = pi42 & pi49;
  assign n10994 = pi36 & pi55;
  assign n10995 = ~n10993 ^ ~n10994;
  assign n10996 = pi34 & pi57;
  assign n10997 = ~n10995 ^ n10996;
  assign n10998 = ~n10992 ^ n10997;
  assign n10999 = n10887 & ~n10890;
  assign n11000 = ~n10883 & ~n10886;
  assign n11001 = ~n10999 & ~n11000;
  assign n11002 = ~n10998 ^ ~n11001;
  assign n11003 = ~n10989 ^ ~n11002;
  assign n11004 = n10868 & ~n10869;
  assign n11005 = ~n10866 & ~n10867;
  assign n11006 = ~n11004 & ~n11005;
  assign n11007 = pi33 & pi58;
  assign n11008 = pi32 & pi59;
  assign n11009 = ~n11007 ^ ~n11008;
  assign n11010 = ~n11009 ^ n6368;
  assign n11011 = pi39 & pi52;
  assign n11012 = pi38 & pi53;
  assign n11013 = ~n11011 ^ ~n11012;
  assign n11014 = pi37 & pi54;
  assign n11015 = ~n11013 ^ n11014;
  assign n11016 = ~n11010 ^ ~n11015;
  assign n11017 = ~n11006 ^ ~n11016;
  assign n11018 = ~n11003 ^ n11017;
  assign n11019 = ~n10986 ^ n11018;
  assign n11020 = n10862 & ~n10875;
  assign n11021 = ~n10847 & n10861;
  assign n11022 = ~n11020 & ~n11021;
  assign n11023 = ~n10850 & n10860;
  assign n11024 = ~n10854 & ~n10859;
  assign n11025 = ~n11023 & ~n11024;
  assign n11026 = n10902 & ~n10907;
  assign n11027 = ~n10896 & ~n10901;
  assign n11028 = ~n11026 & ~n11027;
  assign n11029 = n10905 & ~n10906;
  assign n11030 = ~n10903 & ~n10904;
  assign n11031 = ~n11029 & ~n11030;
  assign n11032 = n10894 & ~n10895;
  assign n11033 = ~n10892 & ~n10893;
  assign n11034 = ~n11032 & ~n11033;
  assign n11035 = ~n11031 ^ ~n11034;
  assign n11036 = ~n11035 ^ ~n6626;
  assign n11037 = ~n11028 ^ n11036;
  assign n11038 = ~n11025 ^ n11037;
  assign n11039 = ~n11022 ^ n11038;
  assign n11040 = ~n10880 & n10909;
  assign n11041 = n10891 & ~n10908;
  assign n11042 = ~n11040 & ~n11041;
  assign n11043 = ~n11039 ^ ~n11042;
  assign n11044 = ~n11019 ^ ~n11043;
  assign n11045 = ~n10951 ^ ~n11044;
  assign n11046 = ~n10948 ^ n11045;
  assign po092 = n10945 ^ n11046;
  assign n11048 = ~n11019 & ~n11043;
  assign n11049 = n10951 & ~n11048;
  assign n11050 = ~n10948 & n11049;
  assign n11051 = n11019 & n11043;
  assign n11052 = ~n11050 & ~n11051;
  assign n11053 = n10948 & ~n10951;
  assign n11054 = ~n11052 & ~n11053;
  assign n11055 = n10945 & ~n11054;
  assign n11056 = ~n11049 & ~n11051;
  assign n11057 = n10948 & n11056;
  assign n11058 = ~n10951 & n11048;
  assign n11059 = ~n11057 & ~n11058;
  assign n11060 = ~n10945 & n11059;
  assign n11061 = ~n11055 & ~n11060;
  assign n11062 = ~n10948 & n10951;
  assign n11063 = n11062 & n11051;
  assign n11064 = n10948 & n11058;
  assign n11065 = ~n11063 & ~n11064;
  assign n11066 = ~n11061 & n11065;
  assign n11067 = n10986 & ~n11018;
  assign n11068 = n10954 & ~n10985;
  assign n11069 = ~n11067 & ~n11068;
  assign n11070 = n11039 & n11042;
  assign n11071 = ~n11022 & n11038;
  assign n11072 = ~n11070 & ~n11071;
  assign n11073 = n11003 & ~n11017;
  assign n11074 = ~n10989 & ~n11002;
  assign n11075 = ~n11073 & ~n11074;
  assign n11076 = ~n11072 ^ n11075;
  assign n11077 = ~n11038 & n11036;
  assign n11078 = ~n11025 & ~n11028;
  assign n11079 = ~n11077 & ~n11078;
  assign n11080 = n11035 & n6626;
  assign n11081 = n11031 & n11034;
  assign n11082 = ~n11080 & ~n11081;
  assign n11083 = ~n10969 & ~pi45;
  assign n11084 = ~n11083 & pi46;
  assign n11085 = pi31 & pi61;
  assign n11086 = pi30 & pi62;
  assign n11087 = ~n11085 ^ ~n11086;
  assign n11088 = ~n11084 ^ n11087;
  assign n11089 = pi41 & pi51;
  assign n11090 = pi40 & pi52;
  assign n11091 = ~n11089 ^ ~n11090;
  assign n11092 = pi39 & pi53;
  assign n11093 = ~n11091 ^ n11092;
  assign n11094 = ~n11088 ^ ~n11093;
  assign n11095 = ~n11082 ^ ~n11094;
  assign n11096 = pi42 & pi50;
  assign n11097 = pi35 & pi57;
  assign n11098 = ~n11096 ^ ~n11097;
  assign n11099 = pi34 & pi58;
  assign n11100 = ~n11098 ^ n11099;
  assign n11101 = pi45 & pi47;
  assign n11102 = pi44 & pi48;
  assign n11103 = ~n11101 ^ ~n11102;
  assign n11104 = pi43 & pi49;
  assign n11105 = ~n11103 ^ n11104;
  assign n11106 = ~n11100 ^ ~n11105;
  assign n11107 = pi36 & pi56;
  assign n11108 = pi33 & pi59;
  assign n11109 = ~n11107 ^ ~n11108;
  assign n11110 = pi29 & pi63;
  assign n11111 = ~n11109 ^ n11110;
  assign n11112 = ~n11106 ^ n11111;
  assign n11113 = ~n11095 ^ n11112;
  assign n11114 = ~n11079 ^ ~n11113;
  assign n11115 = ~n11076 ^ ~n11114;
  assign n11116 = ~n11069 ^ ~n11115;
  assign n11117 = n10973 & ~n10984;
  assign n11118 = ~n10957 & ~n10972;
  assign n11119 = ~n11117 & ~n11118;
  assign n11120 = n10998 & n11001;
  assign n11121 = n10992 & ~n10997;
  assign n11122 = ~n11120 & ~n11121;
  assign n11123 = n11013 & ~n11014;
  assign n11124 = ~n11011 & ~n11012;
  assign n11125 = ~n11123 & ~n11124;
  assign n11126 = n10965 & ~n10966;
  assign n11127 = ~n10963 & ~n10964;
  assign n11128 = ~n11126 & ~n11127;
  assign n11129 = ~n11125 ^ ~n11128;
  assign n11130 = n11009 & ~n6368;
  assign n11131 = ~n11007 & ~n11008;
  assign n11132 = ~n11130 & ~n11131;
  assign n11133 = ~n11129 ^ n11132;
  assign n11134 = ~n11122 ^ ~n11133;
  assign n11135 = n10960 & ~n10961;
  assign n11136 = ~n10958 & ~n10959;
  assign n11137 = ~n11135 & ~n11136;
  assign n11138 = pi38 & pi54;
  assign n11139 = pi37 & pi55;
  assign n11140 = ~n11138 ^ ~n11139;
  assign n11141 = pi32 & pi60;
  assign n11142 = ~n11140 ^ n11141;
  assign n11143 = ~n11137 ^ n11142;
  assign n11144 = n10995 & ~n10996;
  assign n11145 = ~n10993 & ~n10994;
  assign n11146 = ~n11144 & ~n11145;
  assign n11147 = ~n11143 ^ ~n11146;
  assign n11148 = ~n11134 ^ ~n11147;
  assign n11149 = n10980 & n10983;
  assign n11150 = n10976 & n10979;
  assign n11151 = ~n11149 & ~n11150;
  assign n11152 = n10968 & n10971;
  assign n11153 = ~n10962 & ~n10967;
  assign n11154 = ~n11152 & ~n11153;
  assign n11155 = n11006 & n11016;
  assign n11156 = ~n11010 & ~n11015;
  assign n11157 = ~n11155 & ~n11156;
  assign n11158 = ~n11154 ^ ~n11157;
  assign n11159 = ~n11151 ^ ~n11158;
  assign n11160 = ~n11148 ^ n11159;
  assign n11161 = ~n11119 ^ n11160;
  assign n11162 = ~n11116 ^ ~n11161;
  assign po093 = ~n11066 ^ n11162;
  assign n11164 = n10945 & ~n11053;
  assign n11165 = ~n11162 & ~n11048;
  assign n11166 = ~n11062 & ~n11165;
  assign n11167 = ~n11164 & n11166;
  assign n11168 = ~n11053 & ~n11162;
  assign n11169 = ~n11168 & ~n11051;
  assign n11170 = ~n10945 & n11169;
  assign n11171 = n11052 & n11162;
  assign n11172 = ~n11170 & ~n11171;
  assign n11173 = ~n11167 & n11172;
  assign n11174 = n11116 & n11161;
  assign n11175 = n11069 & n11115;
  assign n11176 = ~n11174 & ~n11175;
  assign n11177 = n11076 & n11114;
  assign n11178 = n11072 & ~n11075;
  assign n11179 = ~n11177 & ~n11178;
  assign n11180 = n11134 & n11147;
  assign n11181 = ~n11122 & ~n11133;
  assign n11182 = ~n11180 & ~n11181;
  assign n11183 = n11082 & n11094;
  assign n11184 = n11088 & n11093;
  assign n11185 = ~n11183 & ~n11184;
  assign n11186 = n11098 & ~n11099;
  assign n11187 = ~n11096 & ~n11097;
  assign n11188 = ~n11186 & ~n11187;
  assign n11189 = n11103 & ~n11104;
  assign n11190 = ~n11101 & ~n11102;
  assign n11191 = ~n11189 & ~n11190;
  assign n11192 = ~n11188 ^ ~n11191;
  assign n11193 = n11091 & ~n11092;
  assign n11194 = ~n11089 & ~n11090;
  assign n11195 = ~n11193 & ~n11194;
  assign n11196 = ~n11192 ^ ~n11195;
  assign n11197 = ~n11185 ^ ~n11196;
  assign n11198 = n11109 & ~n11110;
  assign n11199 = ~n11107 & ~n11108;
  assign n11200 = ~n11198 & ~n11199;
  assign n11201 = n11140 & ~n11141;
  assign n11202 = ~n11138 & ~n11139;
  assign n11203 = ~n11201 & ~n11202;
  assign n11204 = ~n11200 ^ ~n11203;
  assign n11205 = pi45 & pi46;
  assign n11206 = ~n11205 & ~n11086;
  assign n11207 = ~n11206 & n11085;
  assign n11208 = ~n8803 & ~pi29;
  assign n11209 = pi46 & pi62;
  assign n11210 = ~n11208 & n11209;
  assign n11211 = ~n11207 & ~n11210;
  assign n11212 = ~n11085 & ~pi30;
  assign n11213 = ~n11211 & ~n11212;
  assign n11214 = ~n11204 ^ ~n11213;
  assign n11215 = ~n11197 ^ n11214;
  assign n11216 = n11129 & ~n11132;
  assign n11217 = ~n11125 & ~n11128;
  assign n11218 = ~n11216 & ~n11217;
  assign n11219 = n11106 & ~n11111;
  assign n11220 = ~n11100 & ~n11105;
  assign n11221 = ~n11219 & ~n11220;
  assign n11222 = ~n11218 ^ n11221;
  assign n11223 = n11143 & n11146;
  assign n11224 = n11137 & ~n11142;
  assign n11225 = ~n11223 & ~n11224;
  assign n11226 = ~n11222 ^ n11225;
  assign n11227 = ~n11215 ^ n11226;
  assign n11228 = ~n11182 ^ ~n11227;
  assign n11229 = ~n11179 ^ n11228;
  assign n11230 = ~n11119 & n11160;
  assign n11231 = ~n11148 & n11159;
  assign n11232 = ~n11230 & ~n11231;
  assign n11233 = n11079 & n11113;
  assign n11234 = n11095 & ~n11112;
  assign n11235 = ~n11233 & ~n11234;
  assign n11236 = n11151 & n11158;
  assign n11237 = n11154 & n11157;
  assign n11238 = ~n11236 & ~n11237;
  assign n11239 = pi45 & pi48;
  assign n11240 = pi38 & pi55;
  assign n11241 = ~n11239 ^ ~n11240;
  assign n11242 = pi37 & pi56;
  assign n11243 = ~n11241 ^ n11242;
  assign n11244 = pi44 & pi49;
  assign n11245 = pi43 & pi50;
  assign n11246 = ~n11244 ^ ~n11245;
  assign n11247 = pi42 & pi51;
  assign n11248 = ~n11246 ^ n11247;
  assign n11249 = ~n11243 ^ ~n11248;
  assign n11250 = pi31 & pi62;
  assign n11251 = ~pi46 & pi47;
  assign n11252 = ~n11250 ^ ~n11251;
  assign n11253 = ~n11249 ^ ~n11252;
  assign n11254 = pi39 & pi54;
  assign n11255 = pi36 & pi57;
  assign n11256 = ~n11254 ^ ~n11255;
  assign n11257 = pi35 & pi58;
  assign n11258 = ~n11256 ^ n11257;
  assign n11259 = pi33 & pi60;
  assign n11260 = ~n6762 ^ ~n11259;
  assign n11261 = pi30 & pi63;
  assign n11262 = ~n11260 ^ n11261;
  assign n11263 = ~n11258 ^ ~n11262;
  assign n11264 = pi41 & pi52;
  assign n11265 = pi40 & pi53;
  assign n11266 = ~n11264 ^ ~n11265;
  assign n11267 = pi34 & pi59;
  assign n11268 = ~n11266 ^ n11267;
  assign n11269 = ~n11263 ^ ~n11268;
  assign n11270 = ~n11253 ^ n11269;
  assign n11271 = ~n11238 ^ n11270;
  assign n11272 = ~n11235 ^ n11271;
  assign n11273 = ~n11232 ^ n11272;
  assign n11274 = ~n11229 ^ ~n11273;
  assign n11275 = ~n11176 ^ n11274;
  assign po094 = ~n11173 ^ ~n11275;
  assign n11277 = n11176 & ~n11274;
  assign n11278 = ~n11173 & ~n11277;
  assign n11279 = ~n11176 & n11274;
  assign n11280 = ~n11278 & ~n11279;
  assign n11281 = n11229 & n11273;
  assign n11282 = ~n11179 & n11228;
  assign n11283 = ~n11281 & ~n11282;
  assign n11284 = n11197 & ~n11214;
  assign n11285 = ~n11185 & ~n11196;
  assign n11286 = ~n11284 & ~n11285;
  assign n11287 = n11204 & n11213;
  assign n11288 = n11200 & n11203;
  assign n11289 = ~n11287 & ~n11288;
  assign n11290 = n11263 & n11268;
  assign n11291 = n11258 & n11262;
  assign n11292 = ~n11290 & ~n11291;
  assign n11293 = ~n11289 ^ n11292;
  assign n11294 = n11192 & n11195;
  assign n11295 = n11188 & n11191;
  assign n11296 = ~n11294 & ~n11295;
  assign n11297 = ~n11293 ^ ~n11296;
  assign n11298 = ~n11286 ^ n11297;
  assign n11299 = ~n11253 & n11269;
  assign n11300 = ~n11298 & ~n11299;
  assign n11301 = n11253 & ~n11269;
  assign n11302 = ~n11238 & ~n11301;
  assign n11303 = n11300 & ~n11302;
  assign n11304 = n11298 & n11299;
  assign n11305 = ~n11303 & ~n11304;
  assign n11306 = ~n11305 & n11238;
  assign n11307 = ~n11238 & n11270;
  assign n11308 = ~n11306 & ~n11307;
  assign n11309 = ~n11232 & ~n11235;
  assign n11310 = ~n11298 & ~n11301;
  assign n11311 = ~n11309 & ~n11310;
  assign n11312 = ~n11308 & n11311;
  assign n11313 = n11232 & n11235;
  assign n11314 = n11313 & ~n11305;
  assign n11315 = ~n11312 & ~n11314;
  assign n11316 = ~n11300 & n11271;
  assign n11317 = n11298 & n11302;
  assign n11318 = n11316 & ~n11317;
  assign n11319 = ~n11313 & n11318;
  assign n11320 = n11298 & ~n11301;
  assign n11321 = ~n11303 & ~n11320;
  assign n11322 = n11309 & n11321;
  assign n11323 = ~n11319 & ~n11322;
  assign n11324 = n11315 & n11323;
  assign n11325 = n11182 & n11227;
  assign n11326 = n11215 & ~n11226;
  assign n11327 = ~n11325 & ~n11326;
  assign n11328 = n11222 & ~n11225;
  assign n11329 = n11218 & ~n11221;
  assign n11330 = ~n11328 & ~n11329;
  assign n11331 = pi44 & pi50;
  assign n11332 = pi43 & pi51;
  assign n11333 = ~n11331 ^ ~n11332;
  assign n11334 = pi36 & pi58;
  assign n11335 = ~n11333 ^ n11334;
  assign n11336 = pi42 & pi52;
  assign n11337 = pi41 & pi53;
  assign n11338 = ~n11336 ^ ~n11337;
  assign n11339 = pi40 & pi54;
  assign n11340 = ~n11338 ^ n11339;
  assign n11341 = ~n11335 ^ ~n11340;
  assign n11342 = pi46 & pi48;
  assign n11343 = pi45 & pi49;
  assign n11344 = ~n11342 ^ ~n11343;
  assign n11345 = pi38 & pi56;
  assign n11346 = ~n11344 ^ n11345;
  assign n11347 = ~n11341 ^ ~n11346;
  assign n11348 = ~n11330 ^ ~n11347;
  assign n11349 = n11246 & ~n11247;
  assign n11350 = ~n11244 & ~n11245;
  assign n11351 = ~n11349 & ~n11350;
  assign n11352 = pi39 & pi55;
  assign n11353 = pi37 & pi57;
  assign n11354 = ~n11352 ^ ~n11353;
  assign n11355 = pi34 & pi60;
  assign n11356 = ~n11354 ^ n11355;
  assign n11357 = ~n11351 ^ n11356;
  assign n11358 = pi35 & pi59;
  assign n11359 = ~n6695 ^ ~n11358;
  assign n11360 = pi33 & pi61;
  assign n11361 = ~n11359 ^ n11360;
  assign n11362 = ~n11357 ^ n11361;
  assign n11363 = ~n11348 ^ n11362;
  assign n11364 = n11249 & n11252;
  assign n11365 = ~n11243 & ~n11248;
  assign n11366 = ~n11364 & ~n11365;
  assign n11367 = pi47 & pi62;
  assign n11368 = ~n11367 & ~pi63;
  assign n11369 = ~n11368 & pi31;
  assign n11370 = pi46 & pi47;
  assign n11371 = ~n11369 & ~n11370;
  assign n11372 = pi46 & pi63;
  assign n11373 = ~n10649 & ~n11372;
  assign n11374 = ~n11373 & n9298;
  assign n11375 = ~n11371 & ~n11374;
  assign n11376 = n11241 & ~n11242;
  assign n11377 = ~n11239 & ~n11240;
  assign n11378 = ~n11376 & ~n11377;
  assign n11379 = ~n11375 ^ ~n11378;
  assign n11380 = ~n11366 ^ n11379;
  assign n11381 = n11260 & ~n11261;
  assign n11382 = ~n6762 & ~n11259;
  assign n11383 = ~n11381 & ~n11382;
  assign n11384 = n11256 & ~n11257;
  assign n11385 = ~n11254 & ~n11255;
  assign n11386 = ~n11384 & ~n11385;
  assign n11387 = ~n11383 ^ ~n11386;
  assign n11388 = n11266 & ~n11267;
  assign n11389 = ~n11264 & ~n11265;
  assign n11390 = ~n11388 & ~n11389;
  assign n11391 = ~n11387 ^ ~n11390;
  assign n11392 = ~n11380 ^ n11391;
  assign n11393 = ~n11363 ^ ~n11392;
  assign n11394 = ~n11327 ^ ~n11393;
  assign n11395 = ~n11324 ^ ~n11394;
  assign n11396 = ~n11283 ^ n11395;
  assign po095 = ~n11280 ^ n11396;
  assign n11398 = ~n11280 & ~n11283;
  assign n11399 = ~n11286 & n11297;
  assign n11400 = ~n11317 & ~n11399;
  assign n11401 = n11400 & ~n11304;
  assign n11402 = n11293 & n11296;
  assign n11403 = n11289 & ~n11292;
  assign n11404 = ~n11402 & ~n11403;
  assign n11405 = pi44 & pi51;
  assign n11406 = pi43 & pi52;
  assign n11407 = ~n11405 ^ ~n11406;
  assign n11408 = pi42 & pi53;
  assign n11409 = ~n11407 ^ n11408;
  assign n11410 = pi46 & pi49;
  assign n11411 = pi45 & pi50;
  assign n11412 = ~n11410 ^ ~n11411;
  assign n11413 = pi39 & pi56;
  assign n11414 = ~n11412 ^ n11413;
  assign n11415 = ~n11409 ^ ~n11414;
  assign n11416 = pi33 & pi62;
  assign n11417 = ~pi47 & pi48;
  assign n11418 = ~n11416 ^ ~n11417;
  assign n11419 = ~n11415 ^ ~n11418;
  assign n11420 = ~n11404 ^ ~n11419;
  assign n11421 = n11333 & ~n11334;
  assign n11422 = ~n11331 & ~n11332;
  assign n11423 = ~n11421 & ~n11422;
  assign n11424 = pi41 & pi54;
  assign n11425 = pi34 & pi61;
  assign n11426 = ~n11424 ^ ~n11425;
  assign n11427 = ~n11426 ^ n6698;
  assign n11428 = pi40 & pi55;
  assign n11429 = pi38 & pi57;
  assign n11430 = ~n11428 ^ ~n11429;
  assign n11431 = pi37 & pi58;
  assign n11432 = ~n11430 ^ n11431;
  assign n11433 = ~n11427 ^ ~n11432;
  assign n11434 = ~n11423 ^ n11433;
  assign n11435 = ~n11420 ^ n11434;
  assign n11436 = ~n11401 ^ ~n11435;
  assign n11437 = n11357 & ~n11361;
  assign n11438 = n11351 & ~n11356;
  assign n11439 = ~n11437 & ~n11438;
  assign n11440 = n11354 & ~n11355;
  assign n11441 = ~n11352 & ~n11353;
  assign n11442 = ~n11440 & ~n11441;
  assign n11443 = n11338 & ~n11339;
  assign n11444 = ~n11336 & ~n11337;
  assign n11445 = ~n11443 & ~n11444;
  assign n11446 = ~n11442 ^ ~n11445;
  assign n11447 = n11359 & ~n11360;
  assign n11448 = ~n6695 & ~n11358;
  assign n11449 = ~n11447 & ~n11448;
  assign n11450 = ~n11446 ^ n11449;
  assign n11451 = ~n11439 ^ ~n11450;
  assign n11452 = n11341 & n11346;
  assign n11453 = n11335 & n11340;
  assign n11454 = ~n11452 & ~n11453;
  assign n11455 = ~n11451 ^ n11454;
  assign n11456 = ~n11436 ^ ~n11455;
  assign n11457 = n11327 & n11393;
  assign n11458 = ~n11363 & ~n11392;
  assign n11459 = ~n11457 & ~n11458;
  assign n11460 = ~n11456 ^ ~n11459;
  assign n11461 = n11348 & ~n11362;
  assign n11462 = n11330 & n11347;
  assign n11463 = ~n11461 & ~n11462;
  assign n11464 = n11380 & ~n11391;
  assign n11465 = n11366 & ~n11379;
  assign n11466 = ~n11464 & ~n11465;
  assign n11467 = n11387 & n11390;
  assign n11468 = n11383 & n11386;
  assign n11469 = ~n11467 & ~n11468;
  assign n11470 = ~n11378 & ~n11374;
  assign n11471 = ~n11470 & ~n11371;
  assign n11472 = n11344 & ~n11345;
  assign n11473 = ~n11342 & ~n11343;
  assign n11474 = ~n11472 & ~n11473;
  assign n11475 = pi35 & pi60;
  assign n11476 = pi36 & pi59;
  assign n11477 = ~n11475 ^ ~n11476;
  assign n11478 = ~n11474 ^ ~n11477;
  assign n11479 = ~n11471 ^ ~n11478;
  assign n11480 = ~n11469 ^ n11479;
  assign n11481 = ~n11466 ^ ~n11480;
  assign n11482 = ~n11463 ^ ~n11481;
  assign n11483 = ~n11460 ^ ~n11482;
  assign n11484 = n11398 & ~n11483;
  assign n11485 = ~n11279 & n11283;
  assign n11486 = ~n11278 & n11485;
  assign n11487 = n11486 & n11483;
  assign n11488 = ~n11484 & ~n11487;
  assign n11489 = ~n11488 & ~n11315;
  assign n11490 = ~n11398 & n11483;
  assign n11491 = ~n11486 & ~n11483;
  assign n11492 = ~n11491 & ~n11323;
  assign n11493 = ~n11490 & n11492;
  assign n11494 = ~n11489 & ~n11493;
  assign n11495 = n11315 & ~n11394;
  assign n11496 = n11495 & n11483;
  assign n11497 = n11398 & n11496;
  assign n11498 = n11323 & n11394;
  assign n11499 = n11487 & n11498;
  assign n11500 = ~n11497 & ~n11499;
  assign n11501 = n11315 & ~n11483;
  assign n11502 = n11483 & n11323;
  assign n11503 = ~n11501 & ~n11502;
  assign n11504 = n11395 & ~n11503;
  assign n11505 = n11504 & ~n11496;
  assign n11506 = ~n11398 & n11505;
  assign n11507 = n11503 & ~n11394;
  assign n11508 = ~n11507 & ~n11501;
  assign n11509 = ~n11486 & ~n11508;
  assign n11510 = ~n11507 & ~n11498;
  assign n11511 = n11509 & ~n11510;
  assign n11512 = ~n11506 & ~n11511;
  assign n11513 = n11500 & n11512;
  assign po096 = ~n11494 | ~n11513;
  assign n11515 = ~n11495 & n11323;
  assign n11516 = ~n11490 & ~n11515;
  assign n11517 = ~n11484 & ~n11509;
  assign n11518 = ~n11516 & n11517;
  assign n11519 = n11460 & n11482;
  assign n11520 = ~n11456 & ~n11459;
  assign n11521 = ~n11519 & ~n11520;
  assign n11522 = n11436 & n11455;
  assign n11523 = ~n11401 & ~n11435;
  assign n11524 = ~n11522 & ~n11523;
  assign n11525 = n11463 & n11481;
  assign n11526 = n11466 & n11480;
  assign n11527 = ~n11525 & ~n11526;
  assign n11528 = ~n11469 & n11479;
  assign n11529 = n11471 & n11478;
  assign n11530 = ~n11528 & ~n11529;
  assign n11531 = n11446 & ~n11449;
  assign n11532 = ~n11442 & ~n11445;
  assign n11533 = ~n11531 & ~n11532;
  assign n11534 = pi35 & pi61;
  assign n11535 = pi34 & pi62;
  assign n11536 = ~n11534 ^ ~n11535;
  assign n11537 = pi33 & pi63;
  assign n11538 = ~n11536 ^ n11537;
  assign n11539 = pi43 & pi53;
  assign n11540 = pi42 & pi54;
  assign n11541 = ~n11539 ^ ~n11540;
  assign n11542 = pi41 & pi55;
  assign n11543 = ~n11541 ^ n11542;
  assign n11544 = ~n11538 ^ ~n11543;
  assign n11545 = ~n11533 ^ ~n11544;
  assign n11546 = ~n11530 ^ n11545;
  assign n11547 = n11474 & n11477;
  assign n11548 = n8125 & n9224;
  assign n11549 = ~n11547 & ~n11548;
  assign n11550 = n11430 & ~n11431;
  assign n11551 = ~n11428 & ~n11429;
  assign n11552 = ~n11550 & ~n11551;
  assign n11553 = n11426 & ~n6698;
  assign n11554 = ~n11424 & ~n11425;
  assign n11555 = ~n11553 & ~n11554;
  assign n11556 = ~n11552 ^ ~n11555;
  assign n11557 = ~n11549 ^ n11556;
  assign n11558 = ~n11546 ^ n11557;
  assign n11559 = n11415 & n11418;
  assign n11560 = ~n11409 & ~n11414;
  assign n11561 = ~n11559 & ~n11560;
  assign n11562 = n11407 & ~n11408;
  assign n11563 = ~n11405 & ~n11406;
  assign n11564 = ~n11562 & ~n11563;
  assign n11565 = n11412 & ~n11413;
  assign n11566 = ~n11410 & ~n11411;
  assign n11567 = ~n11565 & ~n11566;
  assign n11568 = ~n11564 ^ ~n11567;
  assign n11569 = ~n11416 & ~pi47;
  assign n11570 = ~n11569 & pi48;
  assign n11571 = ~n11568 ^ n11570;
  assign n11572 = ~n11561 ^ ~n11571;
  assign n11573 = ~n11423 & n11433;
  assign n11574 = n11427 & n11432;
  assign n11575 = ~n11573 & ~n11574;
  assign n11576 = ~n11572 ^ ~n11575;
  assign n11577 = ~n11558 ^ n11576;
  assign n11578 = ~n11527 ^ n11577;
  assign n11579 = n11420 & ~n11434;
  assign n11580 = n11404 & n11419;
  assign n11581 = ~n11579 & ~n11580;
  assign n11582 = n11451 & ~n11454;
  assign n11583 = n11439 & n11450;
  assign n11584 = ~n11582 & ~n11583;
  assign n11585 = pi47 & pi49;
  assign n11586 = pi46 & pi50;
  assign n11587 = ~n11585 ^ ~n11586;
  assign n11588 = pi45 & pi51;
  assign n11589 = ~n11587 ^ n11588;
  assign n11590 = pi44 & pi52;
  assign n11591 = pi39 & pi57;
  assign n11592 = ~n11590 ^ ~n11591;
  assign n11593 = pi38 & pi58;
  assign n11594 = ~n11592 ^ n11593;
  assign n11595 = ~n11589 ^ ~n11594;
  assign n11596 = pi40 & pi56;
  assign n11597 = pi37 & pi59;
  assign n11598 = ~n11596 ^ ~n11597;
  assign n11599 = pi36 & pi60;
  assign n11600 = ~n11598 ^ n11599;
  assign n11601 = ~n11595 ^ n11600;
  assign n11602 = ~n11584 ^ ~n11601;
  assign n11603 = ~n11581 ^ ~n11602;
  assign n11604 = ~n11578 ^ n11603;
  assign n11605 = ~n11524 ^ n11604;
  assign n11606 = ~n11521 ^ ~n11605;
  assign po097 = n11518 ^ n11606;
  assign n11608 = ~n11578 & n11603;
  assign n11609 = n11524 & ~n11608;
  assign n11610 = n11578 & ~n11603;
  assign n11611 = ~n11609 & ~n11610;
  assign n11612 = ~n11521 & ~n11611;
  assign n11613 = n11524 & n11610;
  assign n11614 = ~n11612 & ~n11613;
  assign n11615 = n11518 & n11614;
  assign n11616 = n11521 & n11611;
  assign n11617 = ~n11524 & n11608;
  assign n11618 = ~n11616 & ~n11617;
  assign n11619 = ~n11518 & n11618;
  assign n11620 = ~n11615 & ~n11619;
  assign n11621 = n11521 & n11617;
  assign n11622 = ~n11521 & n11613;
  assign n11623 = ~n11621 & ~n11622;
  assign n11624 = ~n11620 & n11623;
  assign n11625 = ~n11527 & n11577;
  assign n11626 = ~n11558 & n11576;
  assign n11627 = ~n11625 & ~n11626;
  assign n11628 = n11581 & n11602;
  assign n11629 = ~n11584 & ~n11601;
  assign n11630 = ~n11628 & ~n11629;
  assign n11631 = n11533 & n11544;
  assign n11632 = ~n11538 & ~n11543;
  assign n11633 = ~n11631 & ~n11632;
  assign n11634 = n11568 & ~n11570;
  assign n11635 = ~n11564 & ~n11567;
  assign n11636 = ~n11634 & ~n11635;
  assign n11637 = pi47 & pi50;
  assign n11638 = pi46 & pi51;
  assign n11639 = ~n11637 ^ ~n11638;
  assign n11640 = pi40 & pi57;
  assign n11641 = ~n11639 ^ n11640;
  assign n11642 = ~n11636 ^ n11641;
  assign n11643 = pi35 & pi62;
  assign n11644 = ~pi48 & pi49;
  assign n11645 = ~n11643 ^ ~n11644;
  assign n11646 = ~n11642 ^ ~n11645;
  assign n11647 = ~n11633 ^ n11646;
  assign n11648 = n11598 & ~n11599;
  assign n11649 = ~n11596 & ~n11597;
  assign n11650 = ~n11648 & ~n11649;
  assign n11651 = n11536 & ~n11537;
  assign n11652 = ~n11534 & ~n11535;
  assign n11653 = ~n11651 & ~n11652;
  assign n11654 = ~n11650 ^ ~n11653;
  assign n11655 = n11541 & ~n11542;
  assign n11656 = ~n11539 & ~n11540;
  assign n11657 = ~n11655 & ~n11656;
  assign n11658 = ~n11654 ^ ~n11657;
  assign n11659 = ~n11647 ^ ~n11658;
  assign n11660 = ~n11549 & n11556;
  assign n11661 = n11552 & n11555;
  assign n11662 = ~n11660 & ~n11661;
  assign n11663 = n11592 & ~n11593;
  assign n11664 = ~n11590 & ~n11591;
  assign n11665 = ~n11663 & ~n11664;
  assign n11666 = pi36 & pi61;
  assign n11667 = ~n11665 ^ ~n11666;
  assign n11668 = n11587 & ~n11588;
  assign n11669 = ~n11585 & ~n11586;
  assign n11670 = ~n11668 & ~n11669;
  assign n11671 = ~n11667 ^ ~n11670;
  assign n11672 = ~n11662 ^ n11671;
  assign n11673 = n11595 & ~n11600;
  assign n11674 = ~n11589 & ~n11594;
  assign n11675 = ~n11673 & ~n11674;
  assign n11676 = ~n11672 ^ n11675;
  assign n11677 = ~n11659 ^ ~n11676;
  assign n11678 = ~n11630 ^ n11677;
  assign n11679 = ~n11627 ^ ~n11678;
  assign n11680 = n11546 & ~n11557;
  assign n11681 = n11530 & ~n11545;
  assign n11682 = ~n11680 & ~n11681;
  assign n11683 = n11572 & n11575;
  assign n11684 = ~n11561 & ~n11571;
  assign n11685 = ~n11683 & ~n11684;
  assign n11686 = ~n11682 ^ n11685;
  assign n11687 = pi42 & pi55;
  assign n11688 = pi41 & pi56;
  assign n11689 = ~n11687 ^ ~n11688;
  assign n11690 = pi34 & pi63;
  assign n11691 = ~n11689 ^ n11690;
  assign n11692 = pi39 & pi58;
  assign n11693 = pi38 & pi59;
  assign n11694 = ~n11692 ^ ~n11693;
  assign n11695 = pi37 & pi60;
  assign n11696 = ~n11694 ^ n11695;
  assign n11697 = ~n11691 ^ ~n11696;
  assign n11698 = pi43 & pi54;
  assign n11699 = pi44 & pi53;
  assign n11700 = ~n11698 ^ ~n11699;
  assign n11701 = pi45 & pi52;
  assign n11702 = ~n11700 ^ ~n11701;
  assign n11703 = ~n11697 ^ n11702;
  assign n11704 = ~n11686 ^ n11703;
  assign n11705 = ~n11679 ^ ~n11704;
  assign po098 = n11624 ^ n11705;
  assign n11707 = n11521 & ~n11524;
  assign n11708 = n11517 & ~n11707;
  assign n11709 = n11708 & ~n11516;
  assign n11710 = ~n11521 & n11524;
  assign n11711 = ~n11709 & ~n11710;
  assign n11712 = ~n11705 & ~n11610;
  assign n11713 = ~n11711 & ~n11712;
  assign n11714 = n11705 & ~n11608;
  assign n11715 = ~n11616 & n11714;
  assign n11716 = ~n11518 & ~n11715;
  assign n11717 = ~n11521 & n11609;
  assign n11718 = ~n11717 & ~n11714;
  assign n11719 = ~n11716 & ~n11718;
  assign n11720 = ~n11713 & ~n11719;
  assign n11721 = n11679 & n11704;
  assign n11722 = ~n11627 & ~n11678;
  assign n11723 = ~n11721 & ~n11722;
  assign n11724 = ~n11630 & n11677;
  assign n11725 = ~n11659 & ~n11676;
  assign n11726 = ~n11724 & ~n11725;
  assign n11727 = n11686 & ~n11703;
  assign n11728 = n11682 & ~n11685;
  assign n11729 = ~n11727 & ~n11728;
  assign n11730 = n11642 & n11645;
  assign n11731 = n11636 & ~n11641;
  assign n11732 = ~n11730 & ~n11731;
  assign n11733 = n11694 & ~n11695;
  assign n11734 = ~n11692 & ~n11693;
  assign n11735 = ~n11733 & ~n11734;
  assign n11736 = n11689 & ~n11690;
  assign n11737 = ~n11687 & ~n11688;
  assign n11738 = ~n11736 & ~n11737;
  assign n11739 = ~n11735 ^ ~n11738;
  assign n11740 = n11700 & n11701;
  assign n11741 = pi44 & pi54;
  assign n11742 = n11539 & n11741;
  assign n11743 = ~n11740 & ~n11742;
  assign n11744 = ~n11739 ^ n11743;
  assign n11745 = ~n11732 ^ n11744;
  assign n11746 = pi48 & pi50;
  assign n11747 = pi47 & pi51;
  assign n11748 = ~n11746 ^ ~n11747;
  assign n11749 = pi46 & pi52;
  assign n11750 = ~n11748 ^ n11749;
  assign n11751 = pi45 & pi53;
  assign n11752 = pi40 & pi58;
  assign n11753 = ~n11751 ^ ~n11752;
  assign n11754 = pi39 & pi59;
  assign n11755 = ~n11753 ^ n11754;
  assign n11756 = ~n11750 ^ ~n11755;
  assign n11757 = ~n11643 & ~pi48;
  assign n11758 = ~n11757 & pi49;
  assign n11759 = pi37 & pi61;
  assign n11760 = pi36 & pi62;
  assign n11761 = ~n11759 ^ ~n11760;
  assign n11762 = ~n11758 ^ n11761;
  assign n11763 = ~n11756 ^ n11762;
  assign n11764 = ~n11745 ^ n11763;
  assign n11765 = n11667 & n11670;
  assign n11766 = n11665 & n11666;
  assign n11767 = ~n11765 & ~n11766;
  assign n11768 = n11697 & ~n11702;
  assign n11769 = n11691 & n11696;
  assign n11770 = ~n11768 & ~n11769;
  assign n11771 = ~n11767 ^ n11770;
  assign n11772 = n11654 & n11657;
  assign n11773 = n11650 & n11653;
  assign n11774 = ~n11772 & ~n11773;
  assign n11775 = ~n11771 ^ n11774;
  assign n11776 = ~n11764 ^ n11775;
  assign n11777 = ~n11729 ^ ~n11776;
  assign n11778 = n11647 & n11658;
  assign n11779 = ~n11633 & n11646;
  assign n11780 = ~n11778 & ~n11779;
  assign n11781 = n11672 & ~n11675;
  assign n11782 = ~n11662 & n11671;
  assign n11783 = ~n11781 & ~n11782;
  assign n11784 = ~n11780 ^ ~n11783;
  assign n11785 = n11639 & ~n11640;
  assign n11786 = ~n11637 & ~n11638;
  assign n11787 = ~n11785 & ~n11786;
  assign n11788 = pi42 & pi56;
  assign n11789 = pi41 & pi57;
  assign n11790 = ~n11788 ^ ~n11789;
  assign n11791 = pi38 & pi60;
  assign n11792 = ~n11790 ^ n11791;
  assign n11793 = pi43 & pi55;
  assign n11794 = ~n11741 ^ ~n11793;
  assign n11795 = pi35 & pi63;
  assign n11796 = ~n11794 ^ n11795;
  assign n11797 = ~n11792 ^ ~n11796;
  assign n11798 = ~n11787 ^ ~n11797;
  assign n11799 = ~n11784 ^ n11798;
  assign n11800 = ~n11777 ^ ~n11799;
  assign n11801 = ~n11726 ^ ~n11800;
  assign n11802 = ~n11723 ^ n11801;
  assign po099 = n11720 ^ ~n11802;
  assign n11804 = ~n11723 & n11801;
  assign n11805 = n11720 & ~n11804;
  assign n11806 = n11723 & ~n11801;
  assign n11807 = ~n11805 & ~n11806;
  assign n11808 = n11726 & n11800;
  assign n11809 = ~n11777 & ~n11799;
  assign n11810 = ~n11808 & ~n11809;
  assign n11811 = n11784 & ~n11798;
  assign n11812 = n11780 & n11783;
  assign n11813 = ~n11811 & ~n11812;
  assign n11814 = n11756 & ~n11762;
  assign n11815 = ~n11750 & ~n11755;
  assign n11816 = ~n11814 & ~n11815;
  assign n11817 = ~n10139 & ~pi35;
  assign n11818 = pi49 & pi62;
  assign n11819 = ~n11817 & n11818;
  assign n11820 = ~n11759 & ~pi36;
  assign n11821 = n11819 & ~n11820;
  assign n11822 = pi48 & pi49;
  assign n11823 = ~n11760 & ~n11822;
  assign n11824 = ~n11823 & n11759;
  assign n11825 = ~n11821 & ~n11824;
  assign n11826 = n11790 & ~n11791;
  assign n11827 = ~n11788 & ~n11789;
  assign n11828 = ~n11826 & ~n11827;
  assign n11829 = pi39 & pi60;
  assign n11830 = pi38 & pi61;
  assign n11831 = ~n11829 ^ ~n11830;
  assign n11832 = pi36 & pi63;
  assign n11833 = ~n11831 ^ n11832;
  assign n11834 = ~n11828 ^ n11833;
  assign n11835 = ~n11825 ^ ~n11834;
  assign n11836 = ~n11816 ^ ~n11835;
  assign n11837 = n11753 & ~n11754;
  assign n11838 = ~n11751 & ~n11752;
  assign n11839 = ~n11837 & ~n11838;
  assign n11840 = n11794 & ~n11795;
  assign n11841 = ~n11741 & ~n11793;
  assign n11842 = ~n11840 & ~n11841;
  assign n11843 = ~n11839 ^ ~n11842;
  assign n11844 = n11748 & ~n11749;
  assign n11845 = ~n11746 & ~n11747;
  assign n11846 = ~n11844 & ~n11845;
  assign n11847 = ~n11843 ^ ~n11846;
  assign n11848 = ~n11836 ^ n11847;
  assign n11849 = n11739 & ~n11743;
  assign n11850 = n11735 & n11738;
  assign n11851 = ~n11849 & ~n11850;
  assign n11852 = n11787 & n11797;
  assign n11853 = ~n11792 & ~n11796;
  assign n11854 = ~n11852 & ~n11853;
  assign n11855 = pi37 & pi62;
  assign n11856 = ~pi49 & pi50;
  assign n11857 = ~n11855 ^ ~n11856;
  assign n11858 = ~n11854 ^ n11857;
  assign n11859 = ~n11851 ^ n11858;
  assign n11860 = ~n11848 ^ n11859;
  assign n11861 = ~n11813 ^ n11860;
  assign n11862 = n11745 & ~n11763;
  assign n11863 = n11732 & ~n11744;
  assign n11864 = ~n11862 & ~n11863;
  assign n11865 = pi48 & pi51;
  assign n11866 = pi43 & pi56;
  assign n11867 = ~n11865 ^ ~n11866;
  assign n11868 = pi42 & pi57;
  assign n11869 = ~n11867 ^ n11868;
  assign n11870 = pi44 & pi55;
  assign n11871 = pi41 & pi58;
  assign n11872 = ~n11870 ^ ~n11871;
  assign n11873 = pi40 & pi59;
  assign n11874 = ~n11872 ^ n11873;
  assign n11875 = ~n11869 ^ ~n11874;
  assign n11876 = pi47 & pi52;
  assign n11877 = pi46 & pi53;
  assign n11878 = ~n11876 ^ ~n11877;
  assign n11879 = pi45 & pi54;
  assign n11880 = ~n11878 ^ n11879;
  assign n11881 = ~n11875 ^ n11880;
  assign n11882 = ~n11864 ^ ~n11881;
  assign n11883 = n11771 & ~n11774;
  assign n11884 = ~n11767 & n11770;
  assign n11885 = ~n11883 & ~n11884;
  assign n11886 = ~n11882 ^ ~n11885;
  assign n11887 = ~n11861 ^ ~n11886;
  assign n11888 = n11729 & n11776;
  assign n11889 = n11764 & ~n11775;
  assign n11890 = ~n11888 & ~n11889;
  assign n11891 = ~n11887 ^ ~n11890;
  assign n11892 = ~n11810 ^ n11891;
  assign po100 = ~n11807 ^ ~n11892;
  assign n11894 = ~n11810 & n11890;
  assign n11895 = ~n11807 & ~n11894;
  assign n11896 = n11810 & ~n11890;
  assign n11897 = ~n11861 & ~n11886;
  assign n11898 = n11896 & ~n11897;
  assign n11899 = n11861 & n11886;
  assign n11900 = ~n11898 & ~n11899;
  assign n11901 = n11895 & ~n11900;
  assign n11902 = ~n11810 & ~n11886;
  assign n11903 = n11902 & ~n11891;
  assign n11904 = n11810 & n11886;
  assign n11905 = n11890 & ~n11861;
  assign n11906 = ~n11904 & n11905;
  assign n11907 = ~n11903 & ~n11906;
  assign n11908 = n11807 & ~n11907;
  assign n11909 = n11894 & n11897;
  assign n11910 = n11896 & n11899;
  assign n11911 = ~n11909 & ~n11910;
  assign n11912 = ~n11908 & n11911;
  assign n11913 = ~n11901 & n11912;
  assign n11914 = ~n11813 & n11860;
  assign n11915 = n11848 & ~n11859;
  assign n11916 = ~n11914 & ~n11915;
  assign n11917 = n11882 & n11885;
  assign n11918 = ~n11864 & ~n11881;
  assign n11919 = ~n11917 & ~n11918;
  assign n11920 = n11843 & n11846;
  assign n11921 = n11839 & n11842;
  assign n11922 = ~n11920 & ~n11921;
  assign n11923 = pi49 & pi51;
  assign n11924 = pi48 & pi52;
  assign n11925 = ~n11923 ^ ~n11924;
  assign n11926 = pi47 & pi53;
  assign n11927 = ~n11925 ^ n11926;
  assign n11928 = ~n11922 ^ ~n11927;
  assign n11929 = n11825 & n11834;
  assign n11930 = ~n11828 & n11833;
  assign n11931 = ~n11929 & ~n11930;
  assign n11932 = ~n11928 ^ n11931;
  assign n11933 = n11875 & ~n11880;
  assign n11934 = ~n11869 & ~n11874;
  assign n11935 = ~n11933 & ~n11934;
  assign n11936 = ~n11855 & ~pi49;
  assign n11937 = ~n11936 & pi50;
  assign n11938 = pi37 & pi63;
  assign n11939 = ~n11937 & ~n11938;
  assign n11940 = pi49 & pi63;
  assign n11941 = ~n10649 & ~n11940;
  assign n11942 = ~n11941 & n10538;
  assign n11943 = ~n11939 & ~n11942;
  assign n11944 = n11867 & ~n11868;
  assign n11945 = ~n11865 & ~n11866;
  assign n11946 = ~n11944 & ~n11945;
  assign n11947 = ~n11943 ^ ~n11946;
  assign n11948 = ~n11935 ^ n11947;
  assign n11949 = n11878 & ~n11879;
  assign n11950 = ~n11876 & ~n11877;
  assign n11951 = ~n11949 & ~n11950;
  assign n11952 = n11872 & ~n11873;
  assign n11953 = ~n11870 & ~n11871;
  assign n11954 = ~n11952 & ~n11953;
  assign n11955 = ~n11951 ^ ~n11954;
  assign n11956 = n11831 & ~n11832;
  assign n11957 = ~n11829 & ~n11830;
  assign n11958 = ~n11956 & ~n11957;
  assign n11959 = ~n11955 ^ ~n11958;
  assign n11960 = ~n11948 ^ n11959;
  assign n11961 = ~n11932 ^ ~n11960;
  assign n11962 = ~n11919 ^ ~n11961;
  assign n11963 = ~n11916 ^ ~n11962;
  assign n11964 = ~n11851 & n11858;
  assign n11965 = ~n11854 & n11857;
  assign n11966 = ~n11964 & ~n11965;
  assign n11967 = pi45 & pi55;
  assign n11968 = pi44 & pi56;
  assign n11969 = ~n11967 ^ ~n11968;
  assign n11970 = pi43 & pi57;
  assign n11971 = ~n11969 ^ n11970;
  assign n11972 = pi46 & pi54;
  assign n11973 = pi42 & pi58;
  assign n11974 = ~n11972 ^ ~n11973;
  assign n11975 = pi41 & pi59;
  assign n11976 = ~n11974 ^ n11975;
  assign n11977 = ~n11971 ^ ~n11976;
  assign n11978 = pi40 & pi60;
  assign n11979 = pi39 & pi61;
  assign n11980 = ~n11978 ^ ~n11979;
  assign n11981 = pi38 & pi62;
  assign n11982 = ~n11980 ^ n11981;
  assign n11983 = ~n11977 ^ ~n11982;
  assign n11984 = ~n11966 ^ ~n11983;
  assign n11985 = n11836 & ~n11847;
  assign n11986 = n11816 & n11835;
  assign n11987 = ~n11985 & ~n11986;
  assign n11988 = ~n11984 ^ ~n11987;
  assign n11989 = ~n11963 ^ ~n11988;
  assign po101 = ~n11913 ^ ~n11989;
  assign n11991 = ~n11989 & ~n11897;
  assign n11992 = ~n11896 & ~n11991;
  assign n11993 = ~n11895 & n11992;
  assign n11994 = ~n11894 & ~n11989;
  assign n11995 = ~n11994 & ~n11899;
  assign n11996 = n11807 & n11995;
  assign n11997 = n11900 & n11989;
  assign n11998 = ~n11996 & ~n11997;
  assign n11999 = ~n11993 & n11998;
  assign n12000 = n11963 & n11988;
  assign n12001 = n11916 & n11962;
  assign n12002 = ~n12000 & ~n12001;
  assign n12003 = n11919 & n11961;
  assign n12004 = ~n11932 & ~n11960;
  assign n12005 = ~n12003 & ~n12004;
  assign n12006 = n11984 & n11987;
  assign n12007 = ~n11966 & ~n11983;
  assign n12008 = ~n12006 & ~n12007;
  assign n12009 = n11948 & ~n11959;
  assign n12010 = n11935 & ~n11947;
  assign n12011 = ~n12009 & ~n12010;
  assign n12012 = n11955 & n11958;
  assign n12013 = n11951 & n11954;
  assign n12014 = ~n12012 & ~n12013;
  assign n12015 = n11977 & n11982;
  assign n12016 = n11971 & n11976;
  assign n12017 = ~n12015 & ~n12016;
  assign n12018 = n11974 & ~n11975;
  assign n12019 = ~n11972 & ~n11973;
  assign n12020 = ~n12018 & ~n12019;
  assign n12021 = n11980 & ~n11981;
  assign n12022 = ~n11978 & ~n11979;
  assign n12023 = ~n12021 & ~n12022;
  assign n12024 = ~n12020 ^ ~n12023;
  assign n12025 = n11969 & ~n11970;
  assign n12026 = ~n11967 & ~n11968;
  assign n12027 = ~n12025 & ~n12026;
  assign n12028 = ~n12024 ^ n12027;
  assign n12029 = ~n12017 ^ n12028;
  assign n12030 = ~n12014 ^ n12029;
  assign n12031 = ~n12011 ^ ~n12030;
  assign n12032 = ~n12008 ^ n12031;
  assign n12033 = n11928 & ~n11931;
  assign n12034 = n11922 & n11927;
  assign n12035 = ~n12033 & ~n12034;
  assign n12036 = pi49 & pi52;
  assign n12037 = pi48 & pi53;
  assign n12038 = ~n12036 ^ ~n12037;
  assign n12039 = pi44 & pi57;
  assign n12040 = ~n12038 ^ n12039;
  assign n12041 = pi47 & pi54;
  assign n12042 = pi46 & pi55;
  assign n12043 = ~n12041 ^ ~n12042;
  assign n12044 = pi38 & pi63;
  assign n12045 = ~n12043 ^ n12044;
  assign n12046 = ~n12040 ^ ~n12045;
  assign n12047 = pi45 & pi56;
  assign n12048 = pi43 & pi58;
  assign n12049 = ~n12047 ^ ~n12048;
  assign n12050 = pi42 & pi59;
  assign n12051 = ~n12049 ^ n12050;
  assign n12052 = ~n12046 ^ n12051;
  assign n12053 = ~n12035 ^ ~n12052;
  assign n12054 = ~n11946 & ~n11942;
  assign n12055 = ~n12054 & ~n11939;
  assign n12056 = n11925 & ~n11926;
  assign n12057 = ~n11923 & ~n11924;
  assign n12058 = ~n12056 & ~n12057;
  assign n12059 = pi40 & pi61;
  assign n12060 = pi41 & pi60;
  assign n12061 = ~n12059 ^ ~n12060;
  assign n12062 = ~n12058 ^ ~n12061;
  assign n12063 = ~n12055 ^ ~n12062;
  assign n12064 = pi39 & pi62;
  assign n12065 = ~pi50 & pi51;
  assign n12066 = ~n12064 ^ ~n12065;
  assign n12067 = ~n12063 ^ n12066;
  assign n12068 = ~n12053 ^ ~n12067;
  assign n12069 = ~n12032 ^ n12068;
  assign n12070 = ~n12005 ^ n12069;
  assign n12071 = ~n12002 ^ ~n12070;
  assign po102 = ~n11999 ^ ~n12071;
  assign n12073 = ~n12032 & n12068;
  assign n12074 = ~n12005 & ~n12073;
  assign n12075 = n12032 & ~n12068;
  assign n12076 = ~n12074 & ~n12075;
  assign n12077 = n12002 & n12076;
  assign n12078 = n12005 & n12073;
  assign n12079 = ~n12077 & ~n12078;
  assign n12080 = n11999 & ~n12079;
  assign n12081 = n12002 & n12078;
  assign n12082 = ~n12005 & n12075;
  assign n12083 = ~n12002 & n12082;
  assign n12084 = ~n12081 & ~n12083;
  assign n12085 = ~n12080 & n12084;
  assign n12086 = ~n12002 & ~n12076;
  assign n12087 = ~n12086 & ~n12082;
  assign n12088 = ~n11999 & ~n12087;
  assign n12089 = n12085 & ~n12088;
  assign n12090 = n12053 & n12067;
  assign n12091 = ~n12035 & ~n12052;
  assign n12092 = ~n12090 & ~n12091;
  assign n12093 = ~n12014 & n12029;
  assign n12094 = n12017 & ~n12028;
  assign n12095 = ~n12093 & ~n12094;
  assign n12096 = ~n12092 ^ n12095;
  assign n12097 = n12024 & ~n12027;
  assign n12098 = ~n12020 & ~n12023;
  assign n12099 = ~n12097 & ~n12098;
  assign n12100 = n12046 & ~n12051;
  assign n12101 = ~n12040 & ~n12045;
  assign n12102 = ~n12100 & ~n12101;
  assign n12103 = ~n12099 ^ n12102;
  assign n12104 = n12043 & ~n12044;
  assign n12105 = ~n12041 & ~n12042;
  assign n12106 = ~n12104 & ~n12105;
  assign n12107 = n12038 & ~n12039;
  assign n12108 = ~n12036 & ~n12037;
  assign n12109 = ~n12107 & ~n12108;
  assign n12110 = ~n12106 ^ ~n12109;
  assign n12111 = ~n12064 & ~pi50;
  assign n12112 = ~n12111 & pi51;
  assign n12113 = ~n12110 ^ n12112;
  assign n12114 = ~n12103 ^ ~n12113;
  assign n12115 = ~n12096 ^ n12114;
  assign n12116 = n12063 & ~n12066;
  assign n12117 = ~n12055 & ~n12062;
  assign n12118 = ~n12116 & ~n12117;
  assign n12119 = n12058 & n12061;
  assign n12120 = pi41 & pi61;
  assign n12121 = n11978 & n12120;
  assign n12122 = ~n12119 & ~n12121;
  assign n12123 = n12049 & ~n12050;
  assign n12124 = ~n12047 & ~n12048;
  assign n12125 = ~n12123 & ~n12124;
  assign n12126 = pi42 & pi60;
  assign n12127 = ~n12120 ^ ~n12126;
  assign n12128 = pi39 & pi63;
  assign n12129 = ~n12127 ^ n12128;
  assign n12130 = ~n12125 ^ n12129;
  assign n12131 = ~n12122 ^ n12130;
  assign n12132 = pi50 & pi52;
  assign n12133 = pi49 & pi53;
  assign n12134 = ~n12132 ^ ~n12133;
  assign n12135 = pi48 & pi54;
  assign n12136 = ~n12134 ^ n12135;
  assign n12137 = pi44 & pi58;
  assign n12138 = pi43 & pi59;
  assign n12139 = ~n12137 ^ ~n12138;
  assign n12140 = pi40 & pi62;
  assign n12141 = ~n12139 ^ n12140;
  assign n12142 = ~n12136 ^ ~n12141;
  assign n12143 = pi47 & pi55;
  assign n12144 = pi46 & pi56;
  assign n12145 = ~n12143 ^ ~n12144;
  assign n12146 = pi45 & pi57;
  assign n12147 = ~n12145 ^ n12146;
  assign n12148 = ~n12142 ^ n12147;
  assign n12149 = ~n12131 ^ ~n12148;
  assign n12150 = ~n12118 ^ n12149;
  assign n12151 = ~n12115 ^ n12150;
  assign n12152 = ~n12008 & n12031;
  assign n12153 = n12011 & n12030;
  assign n12154 = ~n12152 & ~n12153;
  assign n12155 = ~n12151 ^ n12154;
  assign po103 = ~n12089 ^ ~n12155;
  assign n12157 = ~n12078 & n12155;
  assign n12158 = ~n12157 & ~n12082;
  assign n12159 = ~n12158 & ~n12002;
  assign n12160 = ~n12076 & n12155;
  assign n12161 = ~n12159 & ~n12160;
  assign n12162 = n11999 & n12161;
  assign n12163 = n12158 & n12002;
  assign n12164 = n12076 & ~n12155;
  assign n12165 = ~n12163 & ~n12164;
  assign n12166 = ~n12162 & n12165;
  assign n12167 = n12151 & ~n12154;
  assign n12168 = n12115 & ~n12150;
  assign n12169 = ~n12167 & ~n12168;
  assign n12170 = n12096 & ~n12114;
  assign n12171 = n12092 & ~n12095;
  assign n12172 = ~n12170 & ~n12171;
  assign n12173 = ~n12150 & ~n12131;
  assign n12174 = ~n12118 & ~n12148;
  assign n12175 = ~n12173 & ~n12174;
  assign n12176 = n12103 & n12113;
  assign n12177 = ~n12099 & n12102;
  assign n12178 = ~n12176 & ~n12177;
  assign n12179 = ~n12122 & n12130;
  assign n12180 = n12125 & ~n12129;
  assign n12181 = ~n12179 & ~n12180;
  assign n12182 = n12110 & ~n12112;
  assign n12183 = ~n12106 & ~n12109;
  assign n12184 = ~n12182 & ~n12183;
  assign n12185 = n12142 & ~n12147;
  assign n12186 = ~n12136 & ~n12141;
  assign n12187 = ~n12185 & ~n12186;
  assign n12188 = ~n12184 ^ n12187;
  assign n12189 = ~n12181 ^ ~n12188;
  assign n12190 = ~n12178 ^ n12189;
  assign n12191 = ~n12175 ^ n12190;
  assign n12192 = n12145 & ~n12146;
  assign n12193 = ~n12143 & ~n12144;
  assign n12194 = ~n12192 & ~n12193;
  assign n12195 = pi40 & pi63;
  assign n12196 = ~n12194 ^ ~n12195;
  assign n12197 = n12134 & ~n12135;
  assign n12198 = ~n12132 & ~n12133;
  assign n12199 = ~n12197 & ~n12198;
  assign n12200 = ~n12196 ^ ~n12199;
  assign n12201 = pi50 & pi53;
  assign n12202 = pi49 & pi54;
  assign n12203 = ~n12201 ^ ~n12202;
  assign n12204 = pi48 & pi55;
  assign n12205 = ~n12203 ^ n12204;
  assign n12206 = pi47 & pi56;
  assign n12207 = pi46 & pi57;
  assign n12208 = ~n12206 ^ ~n12207;
  assign n12209 = pi43 & pi60;
  assign n12210 = ~n12208 ^ n12209;
  assign n12211 = ~n12205 ^ ~n12210;
  assign n12212 = pi41 & pi62;
  assign n12213 = ~pi51 & pi52;
  assign n12214 = ~n12212 ^ n12213;
  assign n12215 = ~n12211 ^ n12214;
  assign n12216 = ~n12200 ^ ~n12215;
  assign n12217 = n12139 & ~n12140;
  assign n12218 = ~n12137 & ~n12138;
  assign n12219 = ~n12217 & ~n12218;
  assign n12220 = pi45 & pi58;
  assign n12221 = pi44 & pi59;
  assign n12222 = ~n12220 ^ ~n12221;
  assign n12223 = ~n12222 ^ n10547;
  assign n12224 = ~n12219 ^ n12223;
  assign n12225 = n12127 & ~n12128;
  assign n12226 = ~n12120 & ~n12126;
  assign n12227 = ~n12225 & ~n12226;
  assign n12228 = ~n12224 ^ ~n12227;
  assign n12229 = ~n12216 ^ ~n12228;
  assign n12230 = ~n12191 ^ n12229;
  assign n12231 = ~n12172 ^ n12230;
  assign n12232 = ~n12169 ^ n12231;
  assign po104 = ~n12166 ^ ~n12232;
  assign n12234 = n12169 & ~n12231;
  assign n12235 = n12165 & ~n12234;
  assign n12236 = ~n12162 & n12235;
  assign n12237 = ~n12169 & n12231;
  assign n12238 = ~n12236 & ~n12237;
  assign n12239 = n12231 & n12191;
  assign n12240 = n12172 & ~n12229;
  assign n12241 = ~n12239 & ~n12240;
  assign n12242 = ~n12175 & n12190;
  assign n12243 = ~n12178 & n12189;
  assign n12244 = ~n12242 & ~n12243;
  assign n12245 = ~n12241 ^ ~n12244;
  assign n12246 = n12181 & n12188;
  assign n12247 = ~n12184 & n12187;
  assign n12248 = ~n12246 & ~n12247;
  assign n12249 = n12216 & n12228;
  assign n12250 = n12200 & n12215;
  assign n12251 = ~n12249 & ~n12250;
  assign n12252 = n12196 & n12199;
  assign n12253 = n12194 & n12195;
  assign n12254 = ~n12252 & ~n12253;
  assign n12255 = pi42 & pi62;
  assign n12256 = ~n12255 & ~pi41;
  assign n12257 = ~pi62 & ~pi63;
  assign n12258 = ~n12256 & ~n12257;
  assign n12259 = pi51 & pi52;
  assign n12260 = ~n12258 & ~n12259;
  assign n12261 = ~pi42 ^ ~pi63;
  assign n12262 = n12261 & ~pi52;
  assign n12263 = n12258 & ~n12262;
  assign n12264 = ~n12260 & ~n12263;
  assign n12265 = ~pi62 & pi63;
  assign n12266 = ~n12265 & pi41;
  assign n12267 = ~n12256 & ~n12266;
  assign n12268 = n12267 & ~n12259;
  assign n12269 = pi52 & pi62;
  assign n12270 = n12269 & pi41;
  assign n12271 = n12270 & ~n12261;
  assign n12272 = ~n12268 & ~n12271;
  assign n12273 = ~n12264 & n12272;
  assign n12274 = ~n12254 ^ ~n12273;
  assign n12275 = n12224 & n12227;
  assign n12276 = n12219 & ~n12223;
  assign n12277 = ~n12275 & ~n12276;
  assign n12278 = ~n12274 ^ n12277;
  assign n12279 = ~n12251 ^ n12278;
  assign n12280 = ~n12248 ^ ~n12279;
  assign n12281 = n12211 & ~n12214;
  assign n12282 = ~n12205 & ~n12210;
  assign n12283 = ~n12281 & ~n12282;
  assign n12284 = pi45 & pi59;
  assign n12285 = pi44 & pi60;
  assign n12286 = ~n12284 ^ ~n12285;
  assign n12287 = pi43 & pi61;
  assign n12288 = ~n12286 ^ n12287;
  assign n12289 = pi51 & pi53;
  assign n12290 = pi50 & pi54;
  assign n12291 = ~n12289 ^ ~n12290;
  assign n12292 = pi49 & pi55;
  assign n12293 = ~n12291 ^ n12292;
  assign n12294 = ~n12288 ^ ~n12293;
  assign n12295 = pi48 & pi56;
  assign n12296 = pi47 & pi57;
  assign n12297 = ~n12295 ^ ~n12296;
  assign n12298 = pi46 & pi58;
  assign n12299 = ~n12297 ^ n12298;
  assign n12300 = ~n12294 ^ ~n12299;
  assign n12301 = ~n12283 ^ ~n12300;
  assign n12302 = n12222 & ~n10547;
  assign n12303 = ~n12220 & ~n12221;
  assign n12304 = ~n12302 & ~n12303;
  assign n12305 = n12208 & ~n12209;
  assign n12306 = ~n12206 & ~n12207;
  assign n12307 = ~n12305 & ~n12306;
  assign n12308 = ~n12304 ^ ~n12307;
  assign n12309 = n12203 & ~n12204;
  assign n12310 = ~n12201 & ~n12202;
  assign n12311 = ~n12309 & ~n12310;
  assign n12312 = ~n12308 ^ ~n12311;
  assign n12313 = ~n12301 ^ ~n12312;
  assign n12314 = ~n12280 ^ ~n12313;
  assign n12315 = ~n12245 ^ n12314;
  assign po105 = ~n12238 ^ ~n12315;
  assign n12317 = n12280 & n12313;
  assign n12318 = ~n12244 & ~n12317;
  assign n12319 = ~n12280 & ~n12313;
  assign n12320 = ~n12318 & ~n12319;
  assign n12321 = ~n12241 & ~n12320;
  assign n12322 = ~n12244 & n12319;
  assign n12323 = ~n12321 & ~n12322;
  assign n12324 = n12238 & n12323;
  assign n12325 = n12244 & n12317;
  assign n12326 = ~n12241 & ~n12325;
  assign n12327 = ~n12326 & n12320;
  assign n12328 = ~n12238 & ~n12327;
  assign n12329 = ~n12324 & ~n12328;
  assign n12330 = ~n12322 & ~n12325;
  assign n12331 = ~n12245 & ~n12330;
  assign n12332 = ~n12329 & ~n12331;
  assign n12333 = n12274 & ~n12277;
  assign n12334 = ~n12254 & ~n12273;
  assign n12335 = ~n12333 & ~n12334;
  assign n12336 = n12294 & n12299;
  assign n12337 = n12288 & n12293;
  assign n12338 = ~n12336 & ~n12337;
  assign n12339 = ~n12335 ^ n12338;
  assign n12340 = n12297 & ~n12298;
  assign n12341 = ~n12295 & ~n12296;
  assign n12342 = ~n12340 & ~n12341;
  assign n12343 = n12291 & ~n12292;
  assign n12344 = ~n12289 & ~n12290;
  assign n12345 = ~n12343 & ~n12344;
  assign n12346 = ~n12342 ^ ~n12345;
  assign n12347 = n12286 & ~n12287;
  assign n12348 = ~n12284 & ~n12285;
  assign n12349 = ~n12347 & ~n12348;
  assign n12350 = ~n12346 ^ ~n12349;
  assign n12351 = ~n12339 ^ n12350;
  assign n12352 = n12301 & n12312;
  assign n12353 = ~n12283 & ~n12300;
  assign n12354 = ~n12352 & ~n12353;
  assign n12355 = ~n11247 & ~pi41;
  assign n12356 = ~pi42 & ~pi63;
  assign n12357 = ~n12356 & n12269;
  assign n12358 = ~n12355 & n12357;
  assign n12359 = pi52 & pi63;
  assign n12360 = n11089 & n12359;
  assign n12361 = pi42 & pi63;
  assign n12362 = n12212 & n12361;
  assign n12363 = ~n12360 & ~n12362;
  assign n12364 = ~n12358 & n12363;
  assign n12365 = pi48 & pi57;
  assign n12366 = pi47 & pi58;
  assign n12367 = ~n12365 ^ ~n12366;
  assign n12368 = pi46 & pi59;
  assign n12369 = ~n12367 ^ n12368;
  assign n12370 = pi45 & pi60;
  assign n12371 = pi44 & pi61;
  assign n12372 = ~n12370 ^ ~n12371;
  assign n12373 = ~n12372 ^ n12361;
  assign n12374 = ~n12369 ^ ~n12373;
  assign n12375 = ~n12364 ^ ~n12374;
  assign n12376 = ~n12354 ^ ~n12375;
  assign n12377 = n12308 & n12311;
  assign n12378 = n12304 & n12307;
  assign n12379 = ~n12377 & ~n12378;
  assign n12380 = pi51 & pi54;
  assign n12381 = pi50 & pi55;
  assign n12382 = ~n12380 ^ ~n12381;
  assign n12383 = pi49 & pi56;
  assign n12384 = ~n12382 ^ n12383;
  assign n12385 = ~n12379 ^ ~n12384;
  assign n12386 = ~pi52 & pi53;
  assign n12387 = ~n10543 ^ ~n12386;
  assign n12388 = ~n12385 ^ n12387;
  assign n12389 = ~n12376 ^ n12388;
  assign n12390 = ~n12351 ^ n12389;
  assign n12391 = n12248 & n12279;
  assign n12392 = ~n12251 & n12278;
  assign n12393 = ~n12391 & ~n12392;
  assign n12394 = ~n12390 ^ n12393;
  assign po106 = n12332 ^ n12394;
  assign n12396 = ~n12331 & n12394;
  assign n12397 = ~n12396 & ~n12327;
  assign n12398 = ~n12238 & ~n12397;
  assign n12399 = n12323 & n12394;
  assign n12400 = n12241 & n12325;
  assign n12401 = ~n12399 & ~n12400;
  assign n12402 = ~n12398 & n12401;
  assign n12403 = n12339 & ~n12350;
  assign n12404 = n12335 & ~n12338;
  assign n12405 = ~n12403 & ~n12404;
  assign n12406 = n12346 & n12349;
  assign n12407 = n12342 & n12345;
  assign n12408 = ~n12406 & ~n12407;
  assign n12409 = pi52 & pi54;
  assign n12410 = pi51 & pi55;
  assign n12411 = ~n12409 ^ ~n12410;
  assign n12412 = pi50 & pi56;
  assign n12413 = ~n12411 ^ n12412;
  assign n12414 = pi49 & pi57;
  assign n12415 = pi48 & pi58;
  assign n12416 = ~n12414 ^ ~n12415;
  assign n12417 = pi47 & pi59;
  assign n12418 = ~n12416 ^ n12417;
  assign n12419 = ~n12413 ^ ~n12418;
  assign n12420 = ~n12408 ^ ~n12419;
  assign n12421 = ~n12405 ^ n12420;
  assign n12422 = n12367 & ~n12368;
  assign n12423 = ~n12365 & ~n12366;
  assign n12424 = ~n12422 & ~n12423;
  assign n12425 = pi46 & pi60;
  assign n12426 = pi45 & pi61;
  assign n12427 = ~n12425 ^ ~n12426;
  assign n12428 = pi44 & pi62;
  assign n12429 = ~n12427 ^ n12428;
  assign n12430 = ~n12424 ^ n12429;
  assign n12431 = n12372 & ~n12361;
  assign n12432 = ~n12370 & ~n12371;
  assign n12433 = ~n12431 & ~n12432;
  assign n12434 = ~n12430 ^ ~n12433;
  assign n12435 = ~n12421 ^ ~n12434;
  assign n12436 = n12376 & ~n12388;
  assign n12437 = ~n12354 & ~n12375;
  assign n12438 = ~n12436 & ~n12437;
  assign n12439 = n12385 & ~n12387;
  assign n12440 = n12379 & n12384;
  assign n12441 = ~n12439 & ~n12440;
  assign n12442 = n12364 & n12374;
  assign n12443 = n12369 & n12373;
  assign n12444 = ~n12442 & ~n12443;
  assign n12445 = ~n12441 ^ ~n12444;
  assign n12446 = n12382 & ~n12383;
  assign n12447 = ~n12380 & ~n12381;
  assign n12448 = ~n12446 & ~n12447;
  assign n12449 = ~n10543 & ~pi52;
  assign n12450 = ~n12449 & pi53;
  assign n12451 = ~n12450 ^ n10650;
  assign n12452 = ~n12448 ^ n12451;
  assign n12453 = ~n12445 ^ n12452;
  assign n12454 = ~n12438 ^ ~n12453;
  assign n12455 = ~n12435 ^ ~n12454;
  assign n12456 = n12390 & ~n12393;
  assign n12457 = ~n12351 & n12389;
  assign n12458 = ~n12456 & ~n12457;
  assign n12459 = ~n12455 ^ n12458;
  assign po107 = n12402 ^ ~n12459;
  assign n12461 = n12455 & ~n12458;
  assign n12462 = n12401 & ~n12461;
  assign n12463 = ~n12398 & n12462;
  assign n12464 = ~n12455 & n12458;
  assign n12465 = ~n12463 & ~n12464;
  assign n12466 = n12435 & n12454;
  assign n12467 = ~n12438 & ~n12453;
  assign n12468 = ~n12466 & ~n12467;
  assign n12469 = n12421 & n12434;
  assign n12470 = n12405 & ~n12420;
  assign n12471 = ~n12469 & ~n12470;
  assign n12472 = n12445 & ~n12452;
  assign n12473 = ~n12441 & ~n12444;
  assign n12474 = ~n12472 & ~n12473;
  assign n12475 = n12411 & ~n12412;
  assign n12476 = ~n12409 & ~n12410;
  assign n12477 = ~n12475 & ~n12476;
  assign n12478 = pi46 & pi61;
  assign n12479 = pi47 & pi60;
  assign n12480 = ~n12478 ^ ~n12479;
  assign n12481 = ~n12477 ^ ~n12480;
  assign n12482 = pi52 & pi55;
  assign n12483 = pi51 & pi56;
  assign n12484 = ~n12482 ^ ~n12483;
  assign n12485 = pi50 & pi57;
  assign n12486 = ~n12484 ^ n12485;
  assign n12487 = ~n12481 ^ n12486;
  assign n12488 = pi45 & pi62;
  assign n12489 = ~pi53 & pi54;
  assign n12490 = ~n12488 ^ ~n12489;
  assign n12491 = ~n12487 ^ ~n12490;
  assign n12492 = n12427 & ~n12428;
  assign n12493 = ~n12425 & ~n12426;
  assign n12494 = ~n12492 & ~n12493;
  assign n12495 = n12416 & ~n12417;
  assign n12496 = ~n12414 & ~n12415;
  assign n12497 = ~n12495 & ~n12496;
  assign n12498 = ~n12494 ^ ~n12497;
  assign n12499 = pi49 & pi58;
  assign n12500 = pi48 & pi59;
  assign n12501 = ~n12499 ^ ~n12500;
  assign n12502 = pi44 & pi63;
  assign n12503 = ~n12501 ^ n12502;
  assign n12504 = ~n12498 ^ n12503;
  assign n12505 = ~n12491 ^ ~n12504;
  assign n12506 = ~n12474 ^ n12505;
  assign n12507 = n12408 & n12419;
  assign n12508 = n12413 & n12418;
  assign n12509 = ~n12507 & ~n12508;
  assign n12510 = n12448 & n12450;
  assign n12511 = ~n12510 & ~n10650;
  assign n12512 = pi52 & pi53;
  assign n12513 = pi53 & pi62;
  assign n12514 = ~n12512 & ~n12513;
  assign n12515 = ~n12448 & n12514;
  assign n12516 = ~n12511 & ~n12515;
  assign n12517 = n12430 & n12433;
  assign n12518 = n12424 & ~n12429;
  assign n12519 = ~n12517 & ~n12518;
  assign n12520 = ~n12516 ^ n12519;
  assign n12521 = ~n12509 ^ ~n12520;
  assign n12522 = ~n12506 ^ n12521;
  assign n12523 = ~n12471 ^ n12522;
  assign n12524 = ~n12468 ^ ~n12523;
  assign po108 = ~n12465 ^ n12524;
  assign n12526 = n12506 & ~n12521;
  assign n12527 = ~n12468 & ~n12471;
  assign n12528 = ~n12506 & n12521;
  assign n12529 = ~n12527 & ~n12528;
  assign n12530 = n12468 & n12471;
  assign n12531 = ~n12529 & ~n12530;
  assign n12532 = ~n12526 & n12531;
  assign n12533 = n12465 & ~n12532;
  assign n12534 = ~n12530 & ~n12526;
  assign n12535 = ~n12534 & n12529;
  assign n12536 = ~n12465 & ~n12535;
  assign n12537 = ~n12533 & ~n12536;
  assign n12538 = n12530 & n12526;
  assign n12539 = n12527 & n12528;
  assign n12540 = ~n12538 & ~n12539;
  assign n12541 = ~n12537 & n12540;
  assign n12542 = ~n12474 & n12505;
  assign n12543 = ~n12491 & ~n12504;
  assign n12544 = ~n12542 & ~n12543;
  assign n12545 = n12509 & n12520;
  assign n12546 = n12516 & ~n12519;
  assign n12547 = ~n12545 & ~n12546;
  assign n12548 = n12501 & ~n12502;
  assign n12549 = ~n12499 & ~n12500;
  assign n12550 = ~n12548 & ~n12549;
  assign n12551 = n12484 & ~n12485;
  assign n12552 = ~n12482 & ~n12483;
  assign n12553 = ~n12551 & ~n12552;
  assign n12554 = ~n12550 ^ ~n12553;
  assign n12555 = ~n12488 & ~pi53;
  assign n12556 = ~n12555 & pi54;
  assign n12557 = ~n12554 ^ n12556;
  assign n12558 = ~n12547 ^ ~n12557;
  assign n12559 = n12477 & n12480;
  assign n12560 = n12478 & n12479;
  assign n12561 = ~n12559 & ~n12560;
  assign n12562 = pi47 & pi61;
  assign n12563 = ~n11209 ^ ~n12562;
  assign n12564 = pi45 & pi63;
  assign n12565 = ~n12563 ^ n12564;
  assign n12566 = pi50 & pi58;
  assign n12567 = pi49 & pi59;
  assign n12568 = ~n12566 ^ ~n12567;
  assign n12569 = pi48 & pi60;
  assign n12570 = ~n12568 ^ n12569;
  assign n12571 = ~n12565 ^ ~n12570;
  assign n12572 = ~n12561 ^ ~n12571;
  assign n12573 = ~n12558 ^ n12572;
  assign n12574 = ~n12544 ^ ~n12573;
  assign n12575 = n12487 & n12490;
  assign n12576 = n12481 & ~n12486;
  assign n12577 = ~n12575 & ~n12576;
  assign n12578 = n12498 & ~n12503;
  assign n12579 = n12494 & n12497;
  assign n12580 = ~n12578 & ~n12579;
  assign n12581 = pi53 & pi55;
  assign n12582 = pi52 & pi56;
  assign n12583 = ~n12581 ^ ~n12582;
  assign n12584 = pi51 & pi57;
  assign n12585 = ~n12583 ^ n12584;
  assign n12586 = ~n12580 ^ ~n12585;
  assign n12587 = ~n12577 ^ n12586;
  assign n12588 = ~n12574 ^ n12587;
  assign po109 = ~n12541 ^ n12588;
  assign n12590 = ~n12530 & ~n12588;
  assign n12591 = ~n12590 & ~n12528;
  assign n12592 = ~n12588 & ~n12526;
  assign n12593 = ~n12527 & ~n12592;
  assign n12594 = ~n12591 & ~n12593;
  assign n12595 = ~n12465 & ~n12594;
  assign n12596 = ~n12531 & n12588;
  assign n12597 = ~n12590 & n12526;
  assign n12598 = ~n12596 & ~n12597;
  assign n12599 = ~n12595 & n12598;
  assign n12600 = n12574 & ~n12587;
  assign n12601 = ~n12544 & ~n12573;
  assign n12602 = ~n12600 & ~n12601;
  assign n12603 = n12558 & ~n12572;
  assign n12604 = ~n12547 & ~n12557;
  assign n12605 = ~n12603 & ~n12604;
  assign n12606 = ~n12602 ^ n12605;
  assign n12607 = ~n12577 & n12586;
  assign n12608 = ~n12580 & ~n12585;
  assign n12609 = ~n12607 & ~n12608;
  assign n12610 = n12568 & ~n12569;
  assign n12611 = ~n12566 & ~n12567;
  assign n12612 = ~n12610 & ~n12611;
  assign n12613 = ~n12612 ^ ~n11372;
  assign n12614 = n12583 & ~n12584;
  assign n12615 = ~n12581 & ~n12582;
  assign n12616 = ~n12614 & ~n12615;
  assign n12617 = ~n12613 ^ ~n12616;
  assign n12618 = n12563 & ~n12564;
  assign n12619 = ~n11209 & ~n12562;
  assign n12620 = ~n12618 & ~n12619;
  assign n12621 = pi53 & pi56;
  assign n12622 = pi52 & pi57;
  assign n12623 = ~n12621 ^ ~n12622;
  assign n12624 = pi51 & pi58;
  assign n12625 = ~n12623 ^ n12624;
  assign n12626 = pi50 & pi59;
  assign n12627 = pi49 & pi60;
  assign n12628 = ~n12626 ^ ~n12627;
  assign n12629 = pi48 & pi61;
  assign n12630 = ~n12628 ^ n12629;
  assign n12631 = ~n12625 ^ ~n12630;
  assign n12632 = ~n12620 ^ ~n12631;
  assign n12633 = ~n12617 ^ ~n12632;
  assign n12634 = ~n12609 ^ n12633;
  assign n12635 = n12561 & n12571;
  assign n12636 = n12565 & n12570;
  assign n12637 = ~n12635 & ~n12636;
  assign n12638 = n12554 & ~n12556;
  assign n12639 = ~n12550 & ~n12553;
  assign n12640 = ~n12638 & ~n12639;
  assign n12641 = ~pi54 & pi55;
  assign n12642 = ~n11367 ^ n12641;
  assign n12643 = ~n12640 ^ n12642;
  assign n12644 = ~n12637 ^ n12643;
  assign n12645 = ~n12634 ^ n12644;
  assign n12646 = ~n12606 ^ n12645;
  assign po110 = n12599 ^ ~n12646;
  assign n12648 = ~n12634 & n12644;
  assign n12649 = n12605 & n12648;
  assign n12650 = n12602 & ~n12649;
  assign n12651 = n12634 & ~n12644;
  assign n12652 = n12605 & ~n12651;
  assign n12653 = ~n12652 & ~n12648;
  assign n12654 = ~n12650 & ~n12653;
  assign n12655 = ~n12599 & n12654;
  assign n12656 = ~n12605 & n12651;
  assign n12657 = ~n12656 & ~n12649;
  assign n12658 = ~n12606 & ~n12657;
  assign n12659 = ~n12655 & ~n12658;
  assign n12660 = n12602 & n12653;
  assign n12661 = ~n12660 & ~n12656;
  assign n12662 = n12599 & ~n12661;
  assign n12663 = n12659 & ~n12662;
  assign n12664 = n12644 & ~n12642;
  assign n12665 = n12637 & n12640;
  assign n12666 = ~n12664 & ~n12665;
  assign n12667 = n12623 & ~n12624;
  assign n12668 = ~n12621 & ~n12622;
  assign n12669 = ~n12667 & ~n12668;
  assign n12670 = pi51 & pi59;
  assign n12671 = pi50 & pi60;
  assign n12672 = ~n12670 ^ ~n12671;
  assign n12673 = pi49 & pi61;
  assign n12674 = ~n12672 ^ n12673;
  assign n12675 = ~n12669 ^ n12674;
  assign n12676 = n12628 & ~n12629;
  assign n12677 = ~n12626 & ~n12627;
  assign n12678 = ~n12676 & ~n12677;
  assign n12679 = ~n12675 ^ n12678;
  assign n12680 = ~n12666 ^ ~n12679;
  assign n12681 = n12620 & n12631;
  assign n12682 = ~n12625 & ~n12630;
  assign n12683 = ~n12681 & ~n12682;
  assign n12684 = ~n12680 ^ n12683;
  assign n12685 = ~n12609 & n12633;
  assign n12686 = n12617 & n12632;
  assign n12687 = ~n12685 & ~n12686;
  assign n12688 = ~n12684 ^ n12687;
  assign n12689 = n12613 & n12616;
  assign n12690 = n12612 & n11372;
  assign n12691 = ~n12689 & ~n12690;
  assign n12692 = pi48 & pi63;
  assign n12693 = ~n12692 & ~pi55;
  assign n12694 = ~n12693 & n11367;
  assign n12695 = pi48 & pi62;
  assign n12696 = pi47 & pi63;
  assign n12697 = ~n12695 & ~n12696;
  assign n12698 = pi54 & pi55;
  assign n12699 = ~n12697 & ~n12698;
  assign n12700 = ~n12694 & n12699;
  assign n12701 = n12697 & n12698;
  assign n12702 = ~pi48 ^ ~pi63;
  assign n12703 = pi55 & pi62;
  assign n12704 = ~n12702 & n12703;
  assign n12705 = n12704 & pi47;
  assign n12706 = ~n12701 & ~n12705;
  assign n12707 = ~n12700 & n12706;
  assign n12708 = pi54 & pi56;
  assign n12709 = pi53 & pi57;
  assign n12710 = ~n12708 ^ ~n12709;
  assign n12711 = pi52 & pi58;
  assign n12712 = ~n12710 ^ n12711;
  assign n12713 = ~n12707 ^ ~n12712;
  assign n12714 = ~n12691 ^ ~n12713;
  assign n12715 = ~n12688 ^ ~n12714;
  assign po111 = n12663 ^ ~n12715;
  assign n12717 = n12602 & ~n12605;
  assign n12718 = ~n12599 & ~n12717;
  assign n12719 = ~n12602 & n12605;
  assign n12720 = n12715 & ~n12651;
  assign n12721 = ~n12719 & ~n12720;
  assign n12722 = ~n12718 & n12721;
  assign n12723 = ~n12602 & n12652;
  assign n12724 = ~n12723 & ~n12715;
  assign n12725 = ~n12599 & ~n12724;
  assign n12726 = ~n12717 & n12715;
  assign n12727 = ~n12726 & ~n12648;
  assign n12728 = ~n12725 & n12727;
  assign n12729 = ~n12722 & ~n12728;
  assign n12730 = n12688 & n12714;
  assign n12731 = ~n12684 & n12687;
  assign n12732 = ~n12730 & ~n12731;
  assign n12733 = n12680 & ~n12683;
  assign n12734 = ~n12666 & ~n12679;
  assign n12735 = ~n12733 & ~n12734;
  assign n12736 = n12691 & n12713;
  assign n12737 = n12707 & n12712;
  assign n12738 = ~n12736 & ~n12737;
  assign n12739 = n12710 & ~n12711;
  assign n12740 = ~n12708 & ~n12709;
  assign n12741 = ~n12739 & ~n12740;
  assign n12742 = n12672 & ~n12673;
  assign n12743 = ~n12670 & ~n12671;
  assign n12744 = ~n12742 & ~n12743;
  assign n12745 = ~n12741 ^ ~n12744;
  assign n12746 = ~n12695 & ~n12698;
  assign n12747 = ~n12746 & n12696;
  assign n12748 = ~n12135 & ~pi47;
  assign n12749 = ~pi48 & ~pi63;
  assign n12750 = ~n12749 & n12703;
  assign n12751 = ~n12748 & n12750;
  assign n12752 = ~n12747 & ~n12751;
  assign n12753 = ~n12745 ^ n12752;
  assign n12754 = ~n12738 ^ ~n12753;
  assign n12755 = n12675 & ~n12678;
  assign n12756 = ~n12669 & n12674;
  assign n12757 = ~n12755 & ~n12756;
  assign n12758 = ~n12754 ^ n12757;
  assign n12759 = pi54 & pi57;
  assign n12760 = pi53 & pi58;
  assign n12761 = ~n12759 ^ ~n12760;
  assign n12762 = pi52 & pi59;
  assign n12763 = ~n12761 ^ n12762;
  assign n12764 = pi51 & pi60;
  assign n12765 = pi50 & pi61;
  assign n12766 = ~n12764 ^ ~n12765;
  assign n12767 = ~n12766 ^ n12692;
  assign n12768 = ~n12763 ^ ~n12767;
  assign n12769 = ~pi55 & pi56;
  assign n12770 = ~n11818 ^ ~n12769;
  assign n12771 = ~n12768 ^ ~n12770;
  assign n12772 = ~n12758 ^ n12771;
  assign n12773 = ~n12735 ^ ~n12772;
  assign n12774 = ~n12732 ^ ~n12773;
  assign po112 = ~n12729 ^ ~n12774;
  assign n12776 = n12758 & ~n12771;
  assign n12777 = n12735 & n12776;
  assign n12778 = n12732 & ~n12777;
  assign n12779 = ~n12735 & ~n12776;
  assign n12780 = ~n12758 & n12771;
  assign n12781 = ~n12779 & ~n12780;
  assign n12782 = ~n12778 & n12781;
  assign n12783 = n12729 & n12782;
  assign n12784 = n12732 & ~n12781;
  assign n12785 = ~n12735 & n12780;
  assign n12786 = ~n12784 & ~n12785;
  assign n12787 = ~n12729 & ~n12786;
  assign n12788 = ~n12783 & ~n12787;
  assign n12789 = n12732 & n12785;
  assign n12790 = ~n12732 & n12777;
  assign n12791 = ~n12789 & ~n12790;
  assign n12792 = n12788 & n12791;
  assign n12793 = n12754 & ~n12757;
  assign n12794 = ~n12738 & ~n12753;
  assign n12795 = ~n12793 & ~n12794;
  assign n12796 = n12766 & ~n12692;
  assign n12797 = ~n12764 & ~n12765;
  assign n12798 = ~n12796 & ~n12797;
  assign n12799 = pi52 & pi60;
  assign n12800 = pi51 & pi61;
  assign n12801 = ~n12799 ^ ~n12800;
  assign n12802 = ~n12801 ^ n11940;
  assign n12803 = ~n12798 ^ n12802;
  assign n12804 = pi55 & pi57;
  assign n12805 = pi54 & pi58;
  assign n12806 = ~n12804 ^ ~n12805;
  assign n12807 = pi53 & pi59;
  assign n12808 = ~n12806 ^ n12807;
  assign n12809 = ~n12803 ^ n12808;
  assign n12810 = ~n12795 ^ ~n12809;
  assign n12811 = n12745 & ~n12752;
  assign n12812 = n12741 & n12744;
  assign n12813 = ~n12811 & ~n12812;
  assign n12814 = n12768 & n12770;
  assign n12815 = ~n12763 & ~n12767;
  assign n12816 = ~n12814 & ~n12815;
  assign n12817 = n12761 & ~n12762;
  assign n12818 = ~n12759 & ~n12760;
  assign n12819 = ~n12817 & ~n12818;
  assign n12820 = ~n11818 & ~pi55;
  assign n12821 = ~n12820 & pi56;
  assign n12822 = pi50 & pi62;
  assign n12823 = ~n12821 ^ ~n12822;
  assign n12824 = ~n12819 ^ n12823;
  assign n12825 = ~n12816 ^ ~n12824;
  assign n12826 = ~n12813 ^ n12825;
  assign n12827 = ~n12810 ^ n12826;
  assign po113 = ~n12792 ^ n12827;
  assign n12829 = ~n12732 & n12735;
  assign n12830 = ~n12729 & ~n12829;
  assign n12831 = n12732 & ~n12735;
  assign n12832 = ~n12827 & ~n12776;
  assign n12833 = ~n12831 & ~n12832;
  assign n12834 = ~n12830 & n12833;
  assign n12835 = n12732 & n12779;
  assign n12836 = ~n12835 & n12827;
  assign n12837 = ~n12729 & ~n12836;
  assign n12838 = ~n12829 & ~n12827;
  assign n12839 = ~n12838 & ~n12780;
  assign n12840 = ~n12837 & n12839;
  assign n12841 = ~n12834 & ~n12840;
  assign n12842 = n12810 & ~n12826;
  assign n12843 = ~n12795 & ~n12809;
  assign n12844 = ~n12842 & ~n12843;
  assign n12845 = n12803 & ~n12808;
  assign n12846 = n12798 & ~n12802;
  assign n12847 = ~n12845 & ~n12846;
  assign n12848 = ~n12819 & n12823;
  assign n12849 = ~n12821 & ~n12822;
  assign n12850 = ~n12848 & ~n12849;
  assign n12851 = n12806 & ~n12807;
  assign n12852 = ~n12804 & ~n12805;
  assign n12853 = ~n12851 & ~n12852;
  assign n12854 = pi52 & pi61;
  assign n12855 = pi53 & pi60;
  assign n12856 = ~n12854 ^ ~n12855;
  assign n12857 = ~n12853 ^ ~n12856;
  assign n12858 = ~n12850 ^ ~n12857;
  assign n12859 = ~n12847 ^ ~n12858;
  assign n12860 = n12801 & ~n11940;
  assign n12861 = ~n12799 & ~n12800;
  assign n12862 = ~n12860 & ~n12861;
  assign n12863 = pi55 & pi58;
  assign n12864 = pi54 & pi59;
  assign n12865 = ~n12863 ^ ~n12864;
  assign n12866 = pi50 & pi63;
  assign n12867 = ~n12865 ^ n12866;
  assign n12868 = ~n12862 ^ n12867;
  assign n12869 = pi51 & pi62;
  assign n12870 = ~pi56 & pi57;
  assign n12871 = ~n12869 ^ ~n12870;
  assign n12872 = ~n12868 ^ ~n12871;
  assign n12873 = ~n12859 ^ n12872;
  assign n12874 = ~n12813 & n12825;
  assign n12875 = ~n12816 & ~n12824;
  assign n12876 = ~n12874 & ~n12875;
  assign n12877 = ~n12873 ^ ~n12876;
  assign n12878 = ~n12844 ^ n12877;
  assign po114 = n12841 ^ n12878;
  assign n12880 = ~n12844 & n12876;
  assign n12881 = n12859 & ~n12872;
  assign n12882 = ~n12880 & ~n12881;
  assign n12883 = n12844 & ~n12876;
  assign n12884 = ~n12859 & n12872;
  assign n12885 = ~n12883 & ~n12884;
  assign n12886 = ~n12882 & n12885;
  assign n12887 = ~n12841 & n12886;
  assign n12888 = n12883 & n12884;
  assign n12889 = n12880 & n12881;
  assign n12890 = ~n12888 & ~n12889;
  assign n12891 = ~n12887 & n12890;
  assign n12892 = n12883 & ~n12881;
  assign n12893 = ~n12880 & n12884;
  assign n12894 = ~n12892 & ~n12893;
  assign n12895 = n12841 & ~n12894;
  assign n12896 = n12891 & ~n12895;
  assign n12897 = n12847 & n12858;
  assign n12898 = ~n12850 & ~n12857;
  assign n12899 = ~n12897 & ~n12898;
  assign n12900 = n12868 & n12871;
  assign n12901 = n12862 & ~n12867;
  assign n12902 = ~n12900 & ~n12901;
  assign n12903 = pi53 & pi61;
  assign n12904 = ~n12269 ^ ~n12903;
  assign n12905 = pi51 & pi63;
  assign n12906 = ~n12904 ^ n12905;
  assign n12907 = pi56 & pi58;
  assign n12908 = pi55 & pi59;
  assign n12909 = ~n12907 ^ ~n12908;
  assign n12910 = pi54 & pi60;
  assign n12911 = ~n12909 ^ n12910;
  assign n12912 = ~n12906 ^ ~n12911;
  assign n12913 = ~n12902 ^ ~n12912;
  assign n12914 = ~n12899 ^ n12913;
  assign n12915 = n12853 & n12856;
  assign n12916 = n7772 & n12512;
  assign n12917 = ~n12915 & ~n12916;
  assign n12918 = n12865 & ~n12866;
  assign n12919 = ~n12863 & ~n12864;
  assign n12920 = ~n12918 & ~n12919;
  assign n12921 = ~n12917 ^ n12920;
  assign n12922 = ~n12869 & ~pi56;
  assign n12923 = ~n12922 & pi57;
  assign n12924 = ~n12921 ^ n12923;
  assign n12925 = ~n12914 ^ n12924;
  assign po115 = ~n12896 ^ ~n12925;
  assign n12927 = ~n12844 & n12859;
  assign n12928 = n12841 & ~n12927;
  assign n12929 = n12844 & ~n12859;
  assign n12930 = n12876 & ~n12872;
  assign n12931 = n12925 & ~n12930;
  assign n12932 = ~n12929 & ~n12931;
  assign n12933 = ~n12928 & n12932;
  assign n12934 = n12929 & ~n12930;
  assign n12935 = ~n12934 & ~n12925;
  assign n12936 = n12841 & ~n12935;
  assign n12937 = ~n12927 & n12925;
  assign n12938 = ~n12876 & n12872;
  assign n12939 = ~n12937 & ~n12938;
  assign n12940 = ~n12936 & n12939;
  assign n12941 = ~n12933 & ~n12940;
  assign n12942 = n12914 & ~n12924;
  assign n12943 = n12899 & ~n12913;
  assign n12944 = ~n12942 & ~n12943;
  assign n12945 = n12921 & ~n12923;
  assign n12946 = n12917 & ~n12920;
  assign n12947 = ~n12945 & ~n12946;
  assign n12948 = pi56 & pi59;
  assign n12949 = pi55 & pi60;
  assign n12950 = ~n12948 ^ ~n12949;
  assign n12951 = pi54 & pi61;
  assign n12952 = ~n12950 ^ n12951;
  assign n12953 = ~n12947 ^ n12952;
  assign n12954 = ~pi57 & pi58;
  assign n12955 = ~n12513 ^ n12954;
  assign n12956 = ~n12953 ^ n12955;
  assign n12957 = n12902 & n12912;
  assign n12958 = n12906 & n12911;
  assign n12959 = ~n12957 & ~n12958;
  assign n12960 = n12904 & ~n12905;
  assign n12961 = ~n12269 & ~n12903;
  assign n12962 = ~n12960 & ~n12961;
  assign n12963 = ~n12962 ^ ~n12359;
  assign n12964 = n12909 & ~n12910;
  assign n12965 = ~n12907 & ~n12908;
  assign n12966 = ~n12964 & ~n12965;
  assign n12967 = ~n12963 ^ ~n12966;
  assign n12968 = ~n12959 ^ n12967;
  assign n12969 = ~n12956 ^ ~n12968;
  assign n12970 = ~n12944 ^ ~n12969;
  assign po116 = ~n12941 ^ ~n12970;
  assign n12972 = n12959 & n12967;
  assign n12973 = ~n12956 & ~n12972;
  assign n12974 = ~n12959 & ~n12967;
  assign n12975 = ~n12973 & ~n12974;
  assign n12976 = n12956 & n12972;
  assign n12977 = n12944 & ~n12976;
  assign n12978 = n12975 & ~n12977;
  assign n12979 = n12941 & n12978;
  assign n12980 = ~n12944 & n12976;
  assign n12981 = ~n12979 & ~n12980;
  assign n12982 = ~n12956 & n12974;
  assign n12983 = ~n12944 & ~n12982;
  assign n12984 = ~n12975 & ~n12983;
  assign n12985 = ~n12941 & n12984;
  assign n12986 = n12944 & n12982;
  assign n12987 = ~n12985 & ~n12986;
  assign n12988 = n12981 & n12987;
  assign n12989 = n12953 & ~n12955;
  assign n12990 = n12947 & ~n12952;
  assign n12991 = ~n12989 & ~n12990;
  assign n12992 = ~n12265 & pi53;
  assign n12993 = pi57 & pi58;
  assign n12994 = ~n12992 & ~n12993;
  assign n12995 = pi54 & pi62;
  assign n12996 = ~n12995 & ~pi53;
  assign n12997 = n12994 & ~n12996;
  assign n12998 = ~pi54 ^ ~pi63;
  assign n12999 = n12513 & ~n12998;
  assign n13000 = n12999 & pi58;
  assign n13001 = ~n12997 & ~n13000;
  assign n13002 = ~n12996 & ~n12257;
  assign n13003 = n12998 & ~pi58;
  assign n13004 = n13002 & n13003;
  assign n13005 = ~n13002 & n12993;
  assign n13006 = ~n13004 & ~n13005;
  assign n13007 = n13001 & n13006;
  assign n13008 = n12950 & ~n12951;
  assign n13009 = ~n12948 & ~n12949;
  assign n13010 = ~n13008 & ~n13009;
  assign n13011 = ~n13007 ^ n13010;
  assign n13012 = pi57 & pi59;
  assign n13013 = pi56 & pi60;
  assign n13014 = ~n13012 ^ ~n13013;
  assign n13015 = pi55 & pi61;
  assign n13016 = ~n13014 ^ n13015;
  assign n13017 = ~n13011 ^ n13016;
  assign n13018 = n12963 & n12966;
  assign n13019 = n12962 & n12359;
  assign n13020 = ~n13018 & ~n13019;
  assign n13021 = ~n13017 ^ n13020;
  assign n13022 = ~n12991 ^ n13021;
  assign po117 = n12988 ^ n13022;
  assign n13024 = n12987 & ~n12991;
  assign n13025 = n13011 & ~n13016;
  assign n13026 = ~n13007 & n13010;
  assign n13027 = ~n13025 & ~n13026;
  assign n13028 = ~pi58 & pi59;
  assign n13029 = ~n12703 ^ ~n13028;
  assign n13030 = ~n13027 ^ n13029;
  assign n13031 = n13014 & ~n13015;
  assign n13032 = ~n13012 & ~n13013;
  assign n13033 = ~n13031 & ~n13032;
  assign n13034 = pi57 & pi60;
  assign n13035 = pi56 & pi61;
  assign n13036 = ~n13034 ^ ~n13035;
  assign n13037 = pi54 & pi63;
  assign n13038 = ~n13036 ^ n13037;
  assign n13039 = ~n13033 ^ n13038;
  assign n13040 = ~n12759 & ~pi53;
  assign n13041 = ~pi54 & ~pi63;
  assign n13042 = pi58 & pi62;
  assign n13043 = ~n13041 & n13042;
  assign n13044 = ~n13040 & n13043;
  assign n13045 = pi58 & pi63;
  assign n13046 = n12709 & n13045;
  assign n13047 = n12513 & n13037;
  assign n13048 = ~n13046 & ~n13047;
  assign n13049 = ~n13044 & n13048;
  assign n13050 = ~n13039 ^ n13049;
  assign n13051 = ~n13030 ^ n13050;
  assign n13052 = n13024 & n13051;
  assign n13053 = n12981 & ~n13051;
  assign n13054 = ~n13052 & ~n13053;
  assign n13055 = ~n12988 & n12991;
  assign n13056 = ~n13017 & n13020;
  assign n13057 = ~n13055 & ~n13056;
  assign n13058 = n13054 & n13057;
  assign n13059 = n12981 & n12991;
  assign n13060 = ~n13051 & n13056;
  assign n13061 = n13059 & n13060;
  assign n13062 = n13017 & ~n13020;
  assign n13063 = ~n13051 & n13062;
  assign n13064 = n13051 & n13056;
  assign n13065 = ~n13063 & ~n13064;
  assign n13066 = ~n12981 & ~n13065;
  assign n13067 = ~n13061 & ~n13066;
  assign n13068 = ~n13058 & n13067;
  assign n13069 = n12981 & n13051;
  assign n13070 = ~n12986 & ~n13051;
  assign n13071 = ~n12985 & n13070;
  assign n13072 = ~n13071 & n12991;
  assign n13073 = ~n13069 & ~n13072;
  assign n13074 = ~n13073 & ~n13062;
  assign n13075 = n13069 & ~n13024;
  assign n13076 = n13074 & ~n13075;
  assign n13077 = n13024 & n13063;
  assign n13078 = ~n13051 & ~n13056;
  assign n13079 = n13051 & ~n13062;
  assign n13080 = ~n13078 & ~n13079;
  assign n13081 = ~n12987 & n13080;
  assign n13082 = ~n13077 & ~n13081;
  assign n13083 = ~n13076 & n13082;
  assign po118 = ~n13068 | ~n13083;
  assign n13085 = ~n13059 & n12987;
  assign n13086 = ~n13085 & ~n13078;
  assign n13087 = ~n13086 & ~n13064;
  assign n13088 = n13087 & ~n13074;
  assign n13089 = n13030 & ~n13050;
  assign n13090 = n13027 & ~n13029;
  assign n13091 = ~n13089 & ~n13090;
  assign n13092 = n13039 & ~n13049;
  assign n13093 = n13033 & ~n13038;
  assign n13094 = ~n13092 & ~n13093;
  assign n13095 = ~n13091 ^ n13094;
  assign n13096 = n13036 & ~n13037;
  assign n13097 = ~n13034 & ~n13035;
  assign n13098 = ~n13096 & ~n13097;
  assign n13099 = n12703 & pi59;
  assign n13100 = pi58 & pi59;
  assign n13101 = pi55 & pi63;
  assign n13102 = ~n13100 & ~n13101;
  assign n13103 = ~n13099 & n13102;
  assign n13104 = pi59 & pi63;
  assign n13105 = n12863 & n13104;
  assign n13106 = pi59 & pi62;
  assign n13107 = n13101 & n13106;
  assign n13108 = ~n13105 & ~n13107;
  assign n13109 = ~n13103 & n13108;
  assign n13110 = ~n13098 ^ ~n13109;
  assign n13111 = pi57 & pi61;
  assign n13112 = pi58 & pi60;
  assign n13113 = ~n13111 ^ ~n13112;
  assign n13114 = pi56 & pi62;
  assign n13115 = ~n13113 ^ ~n13114;
  assign n13116 = ~n13110 ^ ~n13115;
  assign n13117 = ~n13095 ^ n13116;
  assign po119 = n13088 ^ ~n13117;
  assign n13119 = n13110 & n13115;
  assign n13120 = n13094 & ~n13119;
  assign n13121 = ~n13110 & ~n13115;
  assign n13122 = ~n13120 & ~n13121;
  assign n13123 = n13091 & n13122;
  assign n13124 = ~n13094 & n13119;
  assign n13125 = ~n13123 & ~n13124;
  assign n13126 = n13088 & ~n13125;
  assign n13127 = n13094 & n13121;
  assign n13128 = ~n13127 & ~n13124;
  assign n13129 = ~n13095 & ~n13128;
  assign n13130 = ~n13126 & ~n13129;
  assign n13131 = n13091 & ~n13127;
  assign n13132 = ~n13131 & ~n13122;
  assign n13133 = ~n13088 & n13132;
  assign n13134 = n13130 & ~n13133;
  assign n13135 = ~n13098 & ~pi63;
  assign n13136 = ~n13135 & n13099;
  assign n13137 = ~n13098 & ~n13105;
  assign n13138 = ~n13137 & ~n13102;
  assign n13139 = ~n13136 & ~n13138;
  assign n13140 = n13113 & n13114;
  assign n13141 = n7772 & n12993;
  assign n13142 = ~n13140 & ~n13141;
  assign n13143 = pi56 & pi63;
  assign n13144 = pi58 & pi61;
  assign n13145 = ~n13143 ^ ~n13144;
  assign n13146 = ~n13142 ^ n13145;
  assign n13147 = ~n13139 ^ n13146;
  assign n13148 = pi57 & pi62;
  assign n13149 = ~pi59 & pi60;
  assign n13150 = ~n13148 ^ ~n13149;
  assign n13151 = ~n13147 ^ ~n13150;
  assign po120 = n13134 ^ n13151;
  assign n13153 = ~n13091 & n13094;
  assign n13154 = ~n13153 & n13151;
  assign n13155 = ~n13154 & ~n13119;
  assign n13156 = n13091 & ~n13094;
  assign n13157 = n13151 & ~n13121;
  assign n13158 = ~n13156 & ~n13157;
  assign n13159 = ~n13155 & ~n13158;
  assign n13160 = ~n13088 & ~n13159;
  assign n13161 = ~n13154 & n13121;
  assign n13162 = ~n13151 & ~n13124;
  assign n13163 = n13162 & ~n13123;
  assign n13164 = ~n13161 & ~n13163;
  assign n13165 = ~n13160 & n13164;
  assign n13166 = n13147 & n13150;
  assign n13167 = ~n13139 & n13146;
  assign n13168 = ~n13166 & ~n13167;
  assign n13169 = ~n13142 & n13145;
  assign n13170 = n13045 & n13035;
  assign n13171 = ~n13169 & ~n13170;
  assign n13172 = pi59 & pi61;
  assign n13173 = ~n13042 ^ ~n13172;
  assign n13174 = pi57 & pi63;
  assign n13175 = ~n13173 ^ n13174;
  assign n13176 = ~n13171 ^ ~n13175;
  assign n13177 = ~n13148 & ~pi59;
  assign n13178 = ~n13177 & pi60;
  assign n13179 = ~n13176 ^ n13178;
  assign n13180 = ~n13168 ^ ~n13179;
  assign po121 = ~n13165 ^ ~n13180;
  assign n13182 = n13168 & n13179;
  assign n13183 = n13165 & ~n13182;
  assign n13184 = ~n13168 & ~n13179;
  assign n13185 = ~n13183 & ~n13184;
  assign n13186 = n13176 & ~n13178;
  assign n13187 = n13171 & n13175;
  assign n13188 = ~n13186 & ~n13187;
  assign n13189 = n13173 & ~n13174;
  assign n13190 = ~n13042 & ~n13172;
  assign n13191 = ~n13189 & ~n13190;
  assign n13192 = ~pi60 & pi61;
  assign n13193 = ~n13106 ^ ~n13192;
  assign n13194 = ~n13193 ^ ~n13045;
  assign n13195 = ~n13191 ^ n13194;
  assign n13196 = ~n13188 ^ n13195;
  assign po122 = n13185 ^ ~n13196;
  assign n13198 = ~n13184 & ~n13188;
  assign n13199 = ~n13183 & n13198;
  assign n13200 = ~n13188 & ~n13045;
  assign n13201 = ~n13199 & ~n13200;
  assign n13202 = ~n13191 & ~n13193;
  assign n13203 = ~n13201 & n13202;
  assign n13204 = n13188 & ~n13202;
  assign n13205 = n13191 & n13193;
  assign n13206 = ~n13204 & ~n13205;
  assign n13207 = n13206 & ~n13045;
  assign n13208 = n13185 & n13207;
  assign n13209 = n13188 & n13205;
  assign n13210 = ~n13185 & n13209;
  assign n13211 = ~n13208 & ~n13210;
  assign n13212 = ~n13203 & n13211;
  assign n13213 = n13185 & ~n13209;
  assign n13214 = ~n13206 & n13045;
  assign n13215 = ~n13213 & n13214;
  assign n13216 = n13212 & ~n13215;
  assign n13217 = ~pi61 & ~pi62;
  assign n13218 = ~n13217 & pi60;
  assign n13219 = ~n13218 & pi59;
  assign n13220 = ~n8820 ^ ~n13104;
  assign n13221 = ~n13219 & n13220;
  assign n13222 = ~n13220 & ~n13218;
  assign n13223 = ~n13221 & ~n13222;
  assign po123 = ~n13216 ^ ~n13223;
  assign n13225 = ~n13199 & n13045;
  assign n13226 = ~n13202 & n13223;
  assign n13227 = ~n13225 & ~n13226;
  assign n13228 = ~n13200 & n13223;
  assign n13229 = ~n13228 & ~n13205;
  assign n13230 = n13185 & n13229;
  assign n13231 = n13206 & ~n13223;
  assign n13232 = ~n13230 & ~n13231;
  assign n13233 = ~n13227 & n13232;
  assign n13234 = n7772 & pi59;
  assign n13235 = ~n13104 & pi62;
  assign n13236 = ~n13234 & ~n13235;
  assign n13237 = pi60 & pi63;
  assign n13238 = ~n13192 & ~n13237;
  assign n13239 = ~n13236 & ~n13238;
  assign n13240 = ~n13237 & ~pi62;
  assign n13241 = ~n13239 & ~n13240;
  assign po124 = n13233 ^ n13241;
  assign n13243 = ~pi59 & pi61;
  assign n13244 = n13233 & ~n13243;
  assign n13245 = ~n13244 & n10649;
  assign n13246 = ~n13245 & ~n13217;
  assign n13247 = ~n13246 & ~pi60;
  assign n13248 = ~n10649 & ~pi61;
  assign n13249 = ~n13233 & n13248;
  assign n13250 = ~n13234 & pi63;
  assign n13251 = ~n13250 & ~pi62;
  assign n13252 = ~n13249 & ~n13251;
  assign n13253 = ~n13248 & pi60;
  assign n13254 = pi59 & ~pi61;
  assign n13255 = n10649 & ~n13254;
  assign n13256 = n13253 & ~n13255;
  assign n13257 = n13233 & n13256;
  assign n13258 = n13252 & ~n13257;
  assign po125 = ~n13247 & n13258;
  assign n13260 = n13233 & n9224;
  assign n13261 = ~n13260 & ~pi61;
  assign n13262 = ~n13261 & n10649;
  assign n13263 = n13233 & n7772;
  assign n13264 = ~n13234 & ~pi62;
  assign n13265 = ~n13263 & n13264;
  assign n13266 = n13265 & pi63;
  assign po126 = n13262 | n13266;
  assign po127 = ~n13265 & pi63;
  assign po001 = 1'b0;
  assign po000 = pi00;
endmodule


