// Benchmark "mem_ctrl" written by ABC on Mon Nov 19 13:00:42 2018

module mem_ctrl ( 
    pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008,
    pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017,
    pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026,
    pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035,
    pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044,
    pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053,
    pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062,
    pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071,
    pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080,
    pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089,
    pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098,
    pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107,
    pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116,
    pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125,
    pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134,
    pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143,
    pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152,
    pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161,
    pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170,
    pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179,
    pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188,
    pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197,
    pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206,
    pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215,
    pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224,
    pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233,
    pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242,
    pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251,
    pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260,
    pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269,
    pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278,
    pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287,
    pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296,
    pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305,
    pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314,
    pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323,
    pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332,
    pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341,
    pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350,
    pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359,
    pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368,
    pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377,
    pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386,
    pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395,
    pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404,
    pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413,
    pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422,
    pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431,
    pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440,
    pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449,
    pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458,
    pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467,
    pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476,
    pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485,
    pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494,
    pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503,
    pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512,
    pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521,
    pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530,
    pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539,
    pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548,
    pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557,
    pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566,
    pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575,
    pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584,
    pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593,
    pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602,
    pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611,
    pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620,
    pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629,
    pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638,
    pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647,
    pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656,
    pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665,
    pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674,
    pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683,
    pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692,
    pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701,
    pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710,
    pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719,
    pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728,
    pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737,
    pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746,
    pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755,
    pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764,
    pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773,
    pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782,
    pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791,
    pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800,
    pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809,
    pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818,
    pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827,
    pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836,
    pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845,
    pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854,
    pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863,
    pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872,
    pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881,
    pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890,
    pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899,
    pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908,
    pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917,
    pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926,
    pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935,
    pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944,
    pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953,
    pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962,
    pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971,
    pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980,
    pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989,
    pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998,
    pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007,
    pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016,
    pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025,
    pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034,
    pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043,
    pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052,
    pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061,
    pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070,
    pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079,
    pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088,
    pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097,
    pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106,
    pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115,
    pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124,
    pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133,
    pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142,
    pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151,
    pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160,
    pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169,
    pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178,
    pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187,
    pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196,
    pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203,
    po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008,
    po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017,
    po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026,
    po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035,
    po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044,
    po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053,
    po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062,
    po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071,
    po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080,
    po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089,
    po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098,
    po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107,
    po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116,
    po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125,
    po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134,
    po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143,
    po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152,
    po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161,
    po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170,
    po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179,
    po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188,
    po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197,
    po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206,
    po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215,
    po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224,
    po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233,
    po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242,
    po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251,
    po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260,
    po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269,
    po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278,
    po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287,
    po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296,
    po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305,
    po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314,
    po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323,
    po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332,
    po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341,
    po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350,
    po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359,
    po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368,
    po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377,
    po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386,
    po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395,
    po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404,
    po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413,
    po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422,
    po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431,
    po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440,
    po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449,
    po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458,
    po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467,
    po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476,
    po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485,
    po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494,
    po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503,
    po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512,
    po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521,
    po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530,
    po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539,
    po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548,
    po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557,
    po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566,
    po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575,
    po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584,
    po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593,
    po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602,
    po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611,
    po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620,
    po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629,
    po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638,
    po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647,
    po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656,
    po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665,
    po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674,
    po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683,
    po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692,
    po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701,
    po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710,
    po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719,
    po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728,
    po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737,
    po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746,
    po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755,
    po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764,
    po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773,
    po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782,
    po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791,
    po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800,
    po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809,
    po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818,
    po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827,
    po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836,
    po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845,
    po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854,
    po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863,
    po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872,
    po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881,
    po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890,
    po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899,
    po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908,
    po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917,
    po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926,
    po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935,
    po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944,
    po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953,
    po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962,
    po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971,
    po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980,
    po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989,
    po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998,
    po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007,
    po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016,
    po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025,
    po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034,
    po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043,
    po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052,
    po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061,
    po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070,
    po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079,
    po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088,
    po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097,
    po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106,
    po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115,
    po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124,
    po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133,
    po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142,
    po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151,
    po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160,
    po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169,
    po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178,
    po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187,
    po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196,
    po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205,
    po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214,
    po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223,
    po1224, po1225, po1226, po1227, po1228, po1229, po1230  );
  input  pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007,
    pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016,
    pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025,
    pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034,
    pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043,
    pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052,
    pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061,
    pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070,
    pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079,
    pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088,
    pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097,
    pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106,
    pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115,
    pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124,
    pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133,
    pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142,
    pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151,
    pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160,
    pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169,
    pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178,
    pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187,
    pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196,
    pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205,
    pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214,
    pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223,
    pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232,
    pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241,
    pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250,
    pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259,
    pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268,
    pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277,
    pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286,
    pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295,
    pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304,
    pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313,
    pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322,
    pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331,
    pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340,
    pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349,
    pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358,
    pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367,
    pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376,
    pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385,
    pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394,
    pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403,
    pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412,
    pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421,
    pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430,
    pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439,
    pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448,
    pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457,
    pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466,
    pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475,
    pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484,
    pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493,
    pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502,
    pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511,
    pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520,
    pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529,
    pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538,
    pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547,
    pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556,
    pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565,
    pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574,
    pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583,
    pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592,
    pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601,
    pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610,
    pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619,
    pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628,
    pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637,
    pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646,
    pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655,
    pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664,
    pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673,
    pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682,
    pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691,
    pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700,
    pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709,
    pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718,
    pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727,
    pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736,
    pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745,
    pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754,
    pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763,
    pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772,
    pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781,
    pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790,
    pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799,
    pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808,
    pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817,
    pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826,
    pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835,
    pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844,
    pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853,
    pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862,
    pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871,
    pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880,
    pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889,
    pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898,
    pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907,
    pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916,
    pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925,
    pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934,
    pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943,
    pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952,
    pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961,
    pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970,
    pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979,
    pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988,
    pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997,
    pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006,
    pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015,
    pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024,
    pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033,
    pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042,
    pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051,
    pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060,
    pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069,
    pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078,
    pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087,
    pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096,
    pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105,
    pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114,
    pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123,
    pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132,
    pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141,
    pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150,
    pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159,
    pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168,
    pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177,
    pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186,
    pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195,
    pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203;
  output po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007,
    po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016,
    po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025,
    po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034,
    po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043,
    po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052,
    po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061,
    po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070,
    po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079,
    po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088,
    po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097,
    po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106,
    po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115,
    po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124,
    po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133,
    po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142,
    po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151,
    po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160,
    po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169,
    po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178,
    po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187,
    po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196,
    po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205,
    po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214,
    po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223,
    po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232,
    po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241,
    po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250,
    po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259,
    po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268,
    po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277,
    po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286,
    po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295,
    po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304,
    po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313,
    po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322,
    po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331,
    po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340,
    po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349,
    po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358,
    po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367,
    po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376,
    po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385,
    po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394,
    po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403,
    po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412,
    po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421,
    po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430,
    po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439,
    po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448,
    po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457,
    po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466,
    po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475,
    po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484,
    po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493,
    po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502,
    po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511,
    po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520,
    po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529,
    po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538,
    po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547,
    po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556,
    po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565,
    po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574,
    po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583,
    po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592,
    po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601,
    po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610,
    po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619,
    po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628,
    po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637,
    po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646,
    po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655,
    po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664,
    po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673,
    po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682,
    po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691,
    po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700,
    po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709,
    po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718,
    po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727,
    po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736,
    po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745,
    po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754,
    po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763,
    po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772,
    po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781,
    po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790,
    po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799,
    po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808,
    po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817,
    po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826,
    po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835,
    po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844,
    po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853,
    po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862,
    po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871,
    po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880,
    po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889,
    po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898,
    po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907,
    po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916,
    po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925,
    po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934,
    po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943,
    po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952,
    po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961,
    po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970,
    po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979,
    po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988,
    po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997,
    po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006,
    po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015,
    po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024,
    po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033,
    po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042,
    po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051,
    po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060,
    po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069,
    po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078,
    po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087,
    po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096,
    po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105,
    po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114,
    po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123,
    po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132,
    po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141,
    po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150,
    po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159,
    po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168,
    po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177,
    po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186,
    po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195,
    po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204,
    po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213,
    po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222,
    po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230;
  wire n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
    n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
    n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
    n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
    n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
    n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
    n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
    n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
    n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
    n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
    n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
    n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
    n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
    n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
    n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
    n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
    n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
    n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
    n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
    n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
    n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
    n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
    n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
    n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
    n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
    n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
    n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
    n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
    n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
    n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
    n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2748,
    n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
    n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
    n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
    n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
    n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
    n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
    n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
    n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
    n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
    n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
    n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
    n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
    n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
    n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
    n2889, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
    n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
    n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
    n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2938, n2939, n2940,
    n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
    n2951, n2952, n2953, n2954, n2955, n2956, n2958, n2959, n2960, n2961,
    n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
    n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
    n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
    n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3002,
    n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
    n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
    n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
    n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
    n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3052, n3053,
    n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
    n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
    n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
    n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3093, n3094,
    n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
    n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
    n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
    n3125, n3126, n3127, n3128, n3129, n3131, n3132, n3133, n3134, n3135,
    n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
    n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
    n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
    n3166, n3167, n3168, n3169, n3170, n3172, n3173, n3174, n3175, n3176,
    n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
    n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
    n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
    n3207, n3208, n3209, n3210, n3211, n3212, n3214, n3215, n3216, n3217,
    n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
    n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
    n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
    n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
    n3258, n3259, n3260, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
    n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
    n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
    n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
    n3299, n3300, n3301, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
    n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
    n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
    n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3338, n3339, n3340,
    n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
    n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
    n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
    n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
    n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
    n3392, n3393, n3394, n3395, n3396, n3398, n3399, n3400, n3401, n3402,
    n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
    n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
    n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
    n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3444,
    n3445, n3446, n3447, n3448, n3449, n3450, n3452, n3453, n3454, n3455,
    n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
    n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
    n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
    n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
    n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
    n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
    n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
    n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
    n3537, n3538, n3539, n3540, n3541, n3542, n3544, n3545, n3546, n3547,
    n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
    n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
    n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
    n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3587, n3588, n3589,
    n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
    n3601, n3602, n3603, n3605, n3606, n3608, n3609, n3611, n3612, n3614,
    n3615, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
    n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
    n3636, n3637, n3638, n3639, n3640, n3642, n3643, n3645, n3646, n3648,
    n3650, n3651, n3652, n3653, n3654, n3656, n3658, n3660, n3662, n3663,
    n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
    n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
    n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
    n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
    n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
    n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
    n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
    n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
    n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
    n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
    n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
    n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
    n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
    n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
    n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
    n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
    n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
    n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
    n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
    n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
    n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
    n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
    n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
    n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
    n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
    n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
    n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
    n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
    n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
    n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
    n3964, n3965, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
    n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
    n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
    n3995, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
    n4006, n4007, n4008, n4009, n4010, n4012, n4013, n4014, n4015, n4016,
    n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
    n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
    n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
    n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
    n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
    n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
    n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
    n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
    n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
    n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
    n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
    n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4136, n4137,
    n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
    n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
    n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
    n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
    n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
    n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
    n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
    n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
    n4218, n4219, n4220, n4221, n4222, n4224, n4225, n4226, n4227, n4228,
    n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
    n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
    n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
    n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
    n4269, n4270, n4271, n4272, n4274, n4275, n4276, n4277, n4278, n4280,
    n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
    n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
    n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
    n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4320, n4321, n4322,
    n4323, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
    n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
    n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
    n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
    n4364, n4365, n4366, n4367, n4369, n4370, n4371, n4372, n4373, n4374,
    n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
    n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4393, n4394, n4395,
    n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
    n4406, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4417, n4418,
    n4419, n4420, n4421, n4422, n4424, n4425, n4426, n4427, n4428, n4429,
    n4430, n4431, n4433, n4435, n4436, n4437, n4439, n4440, n4441, n4442,
    n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
    n4453, n4454, n4455, n4457, n4458, n4459, n4460, n4462, n4463, n4464,
    n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
    n4475, n4476, n4477, n4478, n4480, n4481, n4482, n4483, n4484, n4485,
    n4486, n4488, n4489, n4490, n4492, n4493, n4495, n4496, n4497, n4498,
    n4499, n4500, n4502, n4503, n4504, n4505, n4507, n4509, n4510, n4511,
    n4512, n4514, n4515, n4516, n4517, n4518, n4520, n4521, n4523, n4524,
    n4525, n4526, n4528, n4529, n4530, n4532, n4533, n4536, n4537, n4538,
    n4539, n4540, n4541, n4542, n4544, n4545, n4546, n4547, n4549, n4550,
    n4551, n4552, n4553, n4555, n4556, n4558, n4559, n4560, n4561, n4562,
    n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4573,
    n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4583, n4584,
    n4585, n4586, n4587, n4588, n4589, n4590, n4592, n4593, n4594, n4595,
    n4596, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
    n4607, n4609, n4610, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
    n4619, n4620, n4621, n4623, n4624, n4627, n4628, n4629, n4630, n4631,
    n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
    n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
    n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
    n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
    n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
    n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
    n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
    n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
    n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
    n4722, n4723, n4724, n4725, n4726, n4728, n4729, n4730, n4731, n4732,
    n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
    n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4753,
    n4754, n4756, n4757, n4759, n4760, n4761, n4762, n4763, n4765, n4766,
    n4768, n4769, n4773, n4774, n4775, n4776, n4777, n4779, n4780, n4781,
    n4783, n4784, n4786, n4787, n4788, n4789, n4790, n4791, n4793, n4794,
    n4795, n4797, n4798, n4799, n4801, n4802, n4803, n4805, n4806, n4807,
    n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4817, n4818,
    n4819, n4820, n4821, n4822, n4824, n4825, n4826, n4827, n4829, n4830,
    n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4842,
    n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4852, n4853,
    n4854, n4855, n4856, n4857, n4861, n4862, n4863, n4865, n4866, n4869,
    n4870, n4871, n4872, n4875, n4876, n4877, n4879, n4880, n4881, n4884,
    n4885, n4887, n4889, n4890, n4892, n4894, n4895, n4896, n4897, n4898,
    n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
    n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
    n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
    n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
    n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
    n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
    n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
    n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
    n4979, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
    n4990, n4992, n4993, n4995, n4996, n4998, n4999, n5000, n5001, n5002,
    n5003, n5004, n5005, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
    n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
    n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
    n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
    n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
    n5054, n5055, n5056, n5057, n5058, n5060, n5061, n5062, n5063, n5064,
    n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5073, n5074, n5075,
    n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
    n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
    n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
    n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
    n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
    n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
    n5136, n5137, n5138, n5139, n5140, n5142, n5143, n5144, n5145, n5146,
    n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
    n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
    n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
    n5177, n5178, n5180, n5181, n5182, n5183, n5184, n5185, n5187, n5188,
    n5189, n5190, n5191, n5192, n5193, n5195, n5196, n5197, n5198, n5199,
    n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
    n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
    n5220, n5221, n5222, n5223, n5224, n5225, n5227, n5228, n5229, n5230,
    n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
    n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
    n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
    n5261, n5262, n5263, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
    n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
    n5282, n5283, n5284, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
    n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
    n5303, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
    n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5322, n5323, n5324,
    n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
    n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
    n5345, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5355, n5356,
    n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
    n5367, n5368, n5369, n5371, n5372, n5373, n5374, n5376, n5377, n5378,
    n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
    n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
    n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
    n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
    n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
    n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
    n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
    n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5459,
    n5460, n5461, n5462, n5463, n5465, n5466, n5467, n5468, n5469, n5471,
    n5472, n5473, n5474, n5475, n5477, n5478, n5479, n5480, n5481, n5483,
    n5484, n5485, n5486, n5487, n5489, n5490, n5491, n5492, n5493, n5494,
    n5496, n5497, n5498, n5499, n5500, n5502, n5503, n5504, n5505, n5506,
    n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
    n5518, n5519, n5520, n5521, n5523, n5524, n5525, n5526, n5527, n5529,
    n5530, n5531, n5532, n5533, n5535, n5536, n5537, n5538, n5539, n5541,
    n5542, n5543, n5544, n5545, n5547, n5548, n5549, n5550, n5551, n5553,
    n5554, n5555, n5556, n5557, n5559, n5560, n5561, n5562, n5563, n5565,
    n5566, n5567, n5568, n5569, n5571, n5572, n5573, n5574, n5575, n5577,
    n5578, n5579, n5580, n5581, n5583, n5584, n5585, n5586, n5587, n5589,
    n5590, n5591, n5592, n5593, n5595, n5596, n5597, n5598, n5599, n5601,
    n5602, n5603, n5604, n5605, n5607, n5608, n5609, n5610, n5611, n5613,
    n5614, n5615, n5616, n5617, n5619, n5620, n5621, n5622, n5623, n5625,
    n5626, n5627, n5628, n5629, n5631, n5632, n5633, n5634, n5635, n5637,
    n5638, n5639, n5640, n5641, n5643, n5644, n5645, n5646, n5647, n5649,
    n5650, n5651, n5652, n5653, n5655, n5656, n5657, n5658, n5659, n5661,
    n5662, n5663, n5664, n5665, n5667, n5668, n5669, n5670, n5671, n5673,
    n5674, n5675, n5676, n5677, n5679, n5680, n5681, n5682, n5683, n5685,
    n5686, n5687, n5688, n5689, n5691, n5692, n5693, n5694, n5695, n5697,
    n5698, n5699, n5700, n5701, n5703, n5704, n5705, n5706, n5707, n5709,
    n5710, n5711, n5712, n5713, n5715, n5716, n5717, n5718, n5719, n5721,
    n5722, n5723, n5724, n5725, n5727, n5728, n5729, n5730, n5731, n5733,
    n5734, n5735, n5736, n5737, n5739, n5740, n5741, n5742, n5743, n5745,
    n5746, n5747, n5748, n5749, n5751, n5752, n5753, n5754, n5755, n5757,
    n5758, n5759, n5760, n5761, n5763, n5764, n5765, n5766, n5767, n5769,
    n5770, n5771, n5772, n5773, n5775, n5776, n5777, n5778, n5779, n5781,
    n5782, n5783, n5784, n5785, n5787, n5788, n5789, n5790, n5791, n5793,
    n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5802, n5803, n5804,
    n5805, n5806, n5807, n5808, n5809, n5810, n5812, n5813, n5814, n5815,
    n5816, n5818, n5819, n5820, n5821, n5822, n5824, n5825, n5826, n5827,
    n5828, n5830, n5831, n5832, n5833, n5834, n5836, n5837, n5838, n5839,
    n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
    n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
    n5860, n5861, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5871,
    n5872, n5873, n5874, n5875, n5876, n5878, n5879, n5880, n5881, n5882,
    n5883, n5884, n5885, n5886, n5887, n5889, n5890, n5891, n5893, n5894,
    n5895, n5896, n5897, n5898, n5900, n5901, n5902, n5903, n5904, n5906,
    n5907, n5908, n5909, n5910, n5912, n5913, n5914, n5915, n5916, n5918,
    n5919, n5920, n5921, n5922, n5924, n5925, n5926, n5927, n5928, n5930,
    n5931, n5932, n5933, n5934, n5936, n5937, n5938, n5939, n5940, n5942,
    n5943, n5944, n5945, n5946, n5948, n5949, n5950, n5951, n5952, n5954,
    n5955, n5956, n5957, n5958, n5960, n5961, n5962, n5963, n5964, n5966,
    n5967, n5968, n5970, n5971, n5972, n5973, n5974, n5976, n5977, n5978,
    n5980, n5981, n5982, n5983, n5984, n5986, n5987, n5988, n5989, n5990,
    n5992, n5993, n5994, n5995, n5996, n5998, n5999, n6000, n6001, n6002,
    n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6014,
    n6015, n6016, n6017, n6018, n6020, n6021, n6023, n6024, n6025, n6026,
    n6027, n6028, n6029, n6030, n6031, n6033, n6034, n6035, n6036, n6037,
    n6038, n6039, n6041, n6042, n6043, n6046, n6047, n6048, n6049, n6050,
    n6051, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
    n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
    n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
    n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
    n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
    n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
    n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
    n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
    n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
    n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
    n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
    n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6172, n6173,
    n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
    n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
    n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
    n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
    n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
    n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
    n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
    n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
    n6255, n6256, n6257, n6258, n6259, n6260, n6262, n6263, n6264, n6265,
    n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
    n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
    n6286, n6287, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
    n6297, n6298, n6299, n6300, n6301, n6303, n6304, n6305, n6306, n6307,
    n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
    n6318, n6319, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
    n6329, n6330, n6331, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
    n6340, n6341, n6342, n6343, n6344, n6345, n6347, n6348, n6349, n6350,
    n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
    n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
    n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6381,
    n6382, n6383, n6384, n6385, n6386, n6387, n6389, n6390, n6391, n6392,
    n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6401, n6402, n6403,
    n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6413, n6414,
    n6415, n6416, n6417, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
    n6426, n6427, n6428, n6429, n6431, n6432, n6433, n6434, n6435, n6437,
    n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6448, n6449,
    n6450, n6451, n6452, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
    n6461, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6472,
    n6473, n6474, n6475, n6476, n6478, n6479, n6480, n6481, n6482, n6484,
    n6485, n6486, n6487, n6488, n6490, n6491, n6492, n6493, n6494, n6496,
    n6497, n6498, n6499, n6500, n6502, n6503, n6504, n6505, n6506, n6508,
    n6509, n6510, n6511, n6512, n6514, n6515, n6516, n6517, n6518, n6519,
    n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6530, n6531,
    n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6541, n6542,
    n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6552, n6553,
    n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6563, n6564,
    n6565, n6566, n6567, n6568, n6569, n6570, n6572, n6573, n6574, n6575,
    n6576, n6577, n6578, n6579, n6581, n6582, n6583, n6584, n6585, n6586,
    n6587, n6588, n6589, n6590, n6592, n6593, n6594, n6595, n6596, n6597,
    n6598, n6599, n6600, n6601, n6603, n6604, n6605, n6606, n6607, n6608,
    n6609, n6610, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
    n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6630, n6631,
    n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6641, n6642,
    n6643, n6644, n6645, n6646, n6647, n6648, n6650, n6651, n6652, n6653,
    n6654, n6655, n6656, n6657, n6659, n6660, n6661, n6662, n6663, n6664,
    n6665, n6666, n6667, n6668, n6670, n6671, n6672, n6673, n6674, n6675,
    n6676, n6677, n6678, n6679, n6681, n6682, n6683, n6684, n6685, n6686,
    n6687, n6688, n6689, n6690, n6692, n6693, n6694, n6695, n6696, n6697,
    n6698, n6699, n6700, n6701, n6703, n6704, n6705, n6706, n6707, n6708,
    n6709, n6710, n6711, n6712, n6714, n6715, n6716, n6717, n6718, n6719,
    n6720, n6721, n6722, n6723, n6725, n6726, n6727, n6728, n6729, n6730,
    n6731, n6732, n6734, n6735, n6736, n6739, n6740, n6741, n6742, n6743,
    n6744, n6745, n6746, n6747, n6748, n6750, n6751, n6752, n6753, n6754,
    n6755, n6756, n6758, n6760, n6761, n6763, n6764, n6765, n6766, n6767,
    n6768, n6769, n6771, n6772, n6774, n6775, n6777, n6778, n6780, n6781,
    n6783, n6784, n6786, n6787, n6789, n6790, n6792, n6793, n6795, n6796,
    n6798, n6799, n6800, n6801, n6802, n6803, n6805, n6806, n6807, n6809,
    n6810, n6811, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
    n6821, n6822, n6823, n6824, n6825, n6826, n6828, n6829, n6831, n6832,
    n6834, n6835, n6837, n6838, n6840, n6841, n6843, n6844, n6846, n6847,
    n6849, n6850, n6851, n6852, n6853, n6854, n6856, n6857, n6858, n6860,
    n6862, n6863, n6865, n6866, n6868, n6870, n6871, n6872, n6874, n6875,
    n6877, n6878, n6879, n6881, n6882, n6883, n6885, n6886, n6888, n6889,
    n6891, n6892, n6894, n6895, n6897, n6898, n6900, n6901, n6903, n6904,
    n6906, n6907, n6909, n6910, n6912, n6913, n6915, n6916, n6918, n6919,
    n6920, n6922, n6923, n6925, n6926, n6927, n6929, n6930, n6932, n6933,
    n6935, n6936, n6938, n6939, n6941, n6942, n6944, n6945, n6947, n6948,
    n6950, n6951, n6952, n6954, n6955, n6957, n6958, n6960, n6961, n6963,
    n6964, n6966, n6967, n6969, n6970, n6972, n6973, n6975, n6976, n6978,
    n6979, n6981, n6982, n6984, n6985, n6987, n6988, n6990, n6991, n6993,
    n6994, n6996, n6997, n6999, n7000, n7002, n7003, n7005, n7006, n7008,
    n7009, n7011, n7012, n7014, n7015, n7017, n7018, n7020, n7021, n7023,
    n7024, n7026, n7027, n7029, n7030, n7032, n7033, n7035, n7036, n7038,
    n7039, n7041, n7042, n7044, n7045, n7047, n7048, n7050, n7051, n7053,
    n7054, n7056, n7057, n7059, n7060, n7062, n7063, n7065, n7066, n7068,
    n7069, n7071, n7072, n7074, n7075, n7077, n7078, n7080, n7081, n7083,
    n7084, n7086, n7087, n7089, n7090, n7092, n7093, n7095, n7096, n7098,
    n7099, n7101, n7102, n7104, n7105, n7107, n7108, n7110, n7111, n7113,
    n7114, n7116, n7117, n7119, n7120, n7122, n7123, n7125, n7126, n7128,
    n7129, n7131, n7132, n7134, n7135, n7137, n7138, n7140, n7141, n7143,
    n7144, n7146, n7147, n7149, n7150, n7152, n7153, n7155, n7156, n7158,
    n7159, n7161, n7162, n7164, n7165, n7167, n7168, n7170, n7171, n7173,
    n7174, n7176, n7177, n7179, n7180, n7182, n7183, n7185, n7186, n7188,
    n7189, n7191, n7192, n7194, n7195, n7197, n7198, n7200, n7201, n7203,
    n7204, n7206, n7207, n7209, n7210, n7212, n7213, n7215, n7216, n7218,
    n7219, n7221, n7222, n7224, n7225, n7227, n7228, n7230, n7231, n7233,
    n7234, n7236, n7237, n7239, n7240, n7242, n7243, n7245, n7246, n7248,
    n7249, n7251, n7252, n7254, n7255, n7257, n7258, n7260, n7261, n7263,
    n7264, n7266, n7267, n7269, n7270, n7272, n7273, n7275, n7276, n7278,
    n7279, n7281, n7282, n7284, n7285, n7287, n7288, n7290, n7291, n7293,
    n7294, n7296, n7297, n7299, n7300, n7302, n7303, n7304, n7305, n7306,
    n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
    n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7325, n7326, n7328,
    n7329, n7331, n7332, n7334, n7335, n7337, n7338, n7340, n7341, n7343,
    n7344, n7346, n7347, n7348, n7349, n7351, n7352, n7353, n7354, n7356,
    n7357, n7358, n7359, n7361, n7362, n7364, n7365, n7366, n7367, n7369,
    n7370, n7371, n7372, n7374, n7375, n7376, n7377, n7379, n7380, n7381,
    n7382, n7384, n7385, n7386, n7387, n7389, n7390, n7391, n7392, n7394,
    n7395, n7396, n7397, n7399, n7402, n7403, n7405, n7406, n7408, n7409,
    n7411, n7412, n7414, n7415, n7417, n7418, n7420, n7421, n7423, n7424,
    n7426, n7427, n7429, n7430, n7432, n7433, n7435, n7436, n7438, n7439,
    n7441, n7442, n7444, n7445, n7447, n7448, n7450, n7451, n7453, n7454,
    n7456, n7457, n7459, n7460, n7462, n7463, n7465, n7466, n7468, n7469,
    n7471, n7472, n7474, n7475, n7477, n7478, n7480, n7481, n7483, n7484,
    n7486, n7487, n7489, n7490, n7492, n7493, n7495, n7496, n7498, n7499,
    n7501, n7502, n7504, n7505, n7507, n7508, n7510, n7511, n7513, n7514,
    n7516, n7517, n7519, n7520, n7522, n7523, n7525, n7526, n7528, n7529,
    n7531, n7532, n7534, n7535, n7537, n7538, n7540, n7541, n7543, n7544,
    n7546, n7547, n7549, n7550, n7552, n7553, n7555, n7556, n7558, n7559,
    n7561, n7562, n7564, n7565, n7567, n7568, n7570, n7571, n7573, n7574,
    n7576, n7577, n7579, n7580, n7582, n7583, n7585, n7586, n7588, n7589,
    n7591, n7592, n7594, n7595, n7597, n7598, n7600, n7601, n7603, n7604,
    n7606, n7607, n7609, n7610, n7612, n7613, n7615, n7616, n7618, n7619,
    n7621, n7622, n7624, n7625, n7627, n7628, n7630, n7631, n7633, n7634,
    n7636, n7637, n7639, n7640, n7642, n7643, n7645, n7646, n7648, n7649,
    n7651, n7652, n7654, n7655, n7657, n7658, n7660, n7661, n7662, n7663,
    n7664, n7665, n7666, n7667, n7669, n7670, n7672, n7673, n7675, n7676,
    n7678, n7679, n7681, n7682, n7684, n7685, n7687, n7688, n7690, n7691,
    n7693, n7694, n7696, n7697, n7699, n7700, n7702, n7703, n7705, n7706,
    n7708, n7709, n7711, n7712, n7714, n7715, n7717, n7718, n7720, n7721,
    n7723, n7724, n7726, n7727, n7728, n7729, n7730, n7732, n7733, n7734,
    n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
    n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7753, n7754, n7755,
    n7757, n7758, n7759, n7761, n7762, n7763, n7765, n7766, n7767, n7768,
    n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
    n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
    n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
    n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
    n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
    n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
    n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
    n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
    n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
    n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
    n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
    n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
    n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
    n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
    n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
    n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
    n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
    n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
    n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
    n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
    n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
    n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
    n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
    n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
    n8009, n8010, n8012, n8013, n8014, n8016, n8017, n8018, n8020, n8021,
    n8022, n8023, n8025, n8027, n8028, n8029, n8030, n8031, n8033, n8034,
    n8036, n8038, n8039, n8040, n8042, n8043, n8045, n8046, n8047, n8048,
    n8050, n8051, n8052, n8053, n8054, n8055, n8057, n8058, n8059, n8060,
    n8061, n8062, n8064, n8066, n8067, n8068, n8069, n8070, n8072, n8073,
    n8074, n8076, n8077, n8078, n8080, n8081, n8082, n8084, n8085, n8086,
    n8088, n8089, n8090, n8092, n8093, n8094, n8096, n8097, n8098, n8100,
    n8101, n8102, n8103, n8105, n8106, n8107, n8108, n8110, n8111, n8112,
    n8113, n8114, n8116, n8117, n8118, n8119, n8120, n8122, n8123, n8124,
    n8126, n8127, n8128, n8130, n8131, n8132, n8134, n8135, n8136, n8138,
    n8139, n8140, n8142, n8143, n8144, n8146, n8147, n8148, n8149, n8150,
    n8152, n8153, n8154, n8155, n8157, n8158, n8159, n8161, n8162, n8163,
    n8165, n8166, n8167, n8169, n8170, n8171, n8173, n8174, n8175, n8177,
    n8178, n8179, n8181, n8182, n8183, n8185, n8186, n8187, n8189, n8190,
    n8191, n8193, n8194, n8195, n8197, n8198, n8199, n8201, n8202, n8203,
    n8205, n8206, n8207, n8209, n8210, n8211, n8213, n8214, n8215, n8217,
    n8218, n8219, n8221, n8222, n8223, n8225, n8226, n8227, n8229, n8230,
    n8231, n8233, n8234, n8235, n8237, n8238, n8239, n8241, n8242, n8243,
    n8245, n8246, n8247, n8249, n8250, n8251, n8253, n8254, n8255, n8257,
    n8258, n8259, n8261, n8262, n8263, n8265, n8266, n8267, n8269, n8270,
    n8271, n8273, n8274, n8275, n8277, n8278, n8279, n8281, n8282, n8283,
    n8285, n8286, n8287, n8289, n8290, n8291, n8293, n8294, n8295, n8296,
    n8297, n8298, n8299, n8300, n8301, n8303, n8304, n8305, n8307, n8308,
    n8309, n8311, n8312, n8313, n8315, n8316, n8317, n8318, n8319, n8320,
    n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
    n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
    n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
    n8351, n8352, n8353, n8354, n8355, n8356, n8358, n8359, n8360, n8361,
    n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
    n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
    n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
    n8393, n8394, n8395, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
    n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
    n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
    n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8432, n8433, n8434,
    n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
    n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
    n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
    n8465, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
    n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
    n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
    n8496, n8497, n8498, n8499, n8500, n8502, n8503, n8504, n8506, n8507,
    n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
    n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
    n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8538,
    n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
    n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
    n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8567, n8568, n8569,
    n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
    n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
    n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
    n8600, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
    n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
    n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
    n8631, n8632, n8633, n8634, n8635, n8637, n8638, n8639, n8640, n8641,
    n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
    n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
    n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8672,
    n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
    n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
    n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
    n8703, n8704, n8705, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
    n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
    n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
    n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8742, n8743, n8744,
    n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
    n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
    n8765, n8766, n8767, n8768, n8769, n8771, n8772, n8773, n8774, n8775,
    n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
    n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
    n8796, n8797, n8798, n8799, n8801, n8802, n8803, n8804, n8805, n8806,
    n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
    n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
    n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8836, n8837,
    n8838, n8840, n8841, n8842, n8844, n8845, n8846, n8847, n8848, n8849,
    n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
    n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
    n8870, n8871, n8874, n8875, n8876, n8878, n8879, n8880, n8881, n8882,
    n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
    n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
    n8903, n8904, n8905, n8906, n8907, n8908, n8910, n8911, n8912, n8914,
    n8915, n8916, n8918, n8919, n8920, n8922, n8923, n8924, n8925, n8926,
    n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
    n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
    n8947, n8948, n8949, n8950, n8951, n8952, n8954, n8955, n8956, n8958,
    n8959, n8960, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
    n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
    n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
    n8990, n8991, n8992, n8994, n8995, n8996, n8998, n8999, n9000, n9002,
    n9003, n9004, n9006, n9007, n9008, n9010, n9011, n9012, n9014, n9015,
    n9016, n9018, n9019, n9020, n9022, n9023, n9024, n9026, n9027, n9028,
    n9030, n9031, n9032, n9034, n9035, n9036, n9038, n9039, n9040, n9042,
    n9043, n9044, n9046, n9047, n9048, n9050, n9051, n9052, n9053, n9054,
    n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
    n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
    n9075, n9076, n9077, n9078, n9079, n9081, n9082, n9083, n9084, n9085,
    n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
    n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
    n9106, n9107, n9108, n9109, n9110, n9112, n9113, n9114, n9116, n9117,
    n9118, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
    n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
    n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
    n9149, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
    n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
    n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
    n9180, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
    n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
    n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
    n9211, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
    n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
    n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
    n9242, n9243, n9245, n9246, n9247, n9249, n9250, n9251, n9252, n9253,
    n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
    n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
    n9274, n9275, n9276, n9277, n9278, n9280, n9281, n9282, n9283, n9284,
    n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
    n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
    n9305, n9306, n9307, n9308, n9309, n9310, n9312, n9313, n9314, n9315,
    n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
    n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
    n9336, n9337, n9338, n9339, n9340, n9341, n9343, n9344, n9345, n9346,
    n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
    n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
    n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9375, n9376, n9377,
    n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
    n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
    n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9407, n9408,
    n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
    n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9430,
    n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
    n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
    n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
    n9462, n9463, n9464, n9466, n9467, n9468, n9470, n9471, n9472, n9474,
    n9475, n9476, n9478, n9479, n9480, n9482, n9483, n9484, n9486, n9487,
    n9488, n9490, n9491, n9492, n9494, n9495, n9496, n9498, n9499, n9500,
    n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
    n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
    n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
    n9533, n9534, n9535, n9537, n9538, n9539, n9541, n9542, n9543, n9545,
    n9546, n9547, n9549, n9550, n9551, n9554, n9555, n9556, n9558, n9559,
    n9560, n9562, n9563, n9564, n9566, n9567, n9568, n9570, n9571, n9572,
    n9574, n9575, n9576, n9578, n9579, n9580, n9582, n9583, n9585, n9586,
    n9587, n9589, n9590, n9591, n9593, n9594, n9595, n9597, n9598, n9599,
    n9601, n9602, n9603, n9605, n9606, n9607, n9609, n9610, n9611, n9613,
    n9614, n9615, n9617, n9618, n9619, n9621, n9622, n9623, n9625, n9626,
    n9627, n9629, n9630, n9631, n9633, n9634, n9635, n9637, n9638, n9639,
    n9641, n9642, n9643, n9645, n9646, n9647, n9649, n9650, n9651, n9653,
    n9654, n9655, n9656, n9657, n9658, n9659, n9661, n9663, n9664, n9665,
    n9667, n9668, n9669, n9671, n9672, n9673, n9675, n9677, n9678, n9679,
    n9681, n9682, n9683, n9685, n9686, n9687, n9689, n9691, n9692, n9693,
    n9695, n9696, n9697, n9699, n9700, n9701, n9703, n9704, n9705, n9707,
    n9708, n9709, n9710, n9711, n9712, n9713, n9717, n9718, n9720, n9722,
    n9723, n9725, n9726, n9728, n9729, n9731, n9732, n9734, n9735, n9737,
    n9738, n9740, n9741, n9743, n9744, n9746, n9747, n9749, n9750, n9752,
    n9753, n9754, n9756, n9757, n9759, n9760, n9761, n9762, n9763, n9764,
    n9766, n9767, n9769, n9770, n9772, n9773, n9775, n9776, n9779, n9780,
    n9782, n9783, n9786, n9787, n9789, n9790, n9792, n9793, n9795, n9796,
    n9798, n9799, n9801, n9802, n9804, n9805, n9807, n9808, n9810, n9811,
    n9813, n9814, n9819, n9822, n9823, n9824, n9826, n9827, n9828, n9829,
    n9830, n9831, n9832, n9833, n9834, n9835, n9837, n9838, n9839, n9840,
    n9841, n9842, n9843, n9844, n9845, n9847, n9848, n9849, n9850, n9851,
    n9852, n9853, n9854, n9855, n9857, n9858, n9859, n9860, n9861, n9862,
    n9863, n9864, n9865, n9867, n9868, n9869, n9872, n9873, n9875, n9878,
    n9880, n9881, n9883, n9884, n9886, n9887, n9889, n9890, n9892, n9893,
    n9895, n9896, n9898, n9899, n9901, n9902, n9904, n9905, n9907, n9908,
    n9910, n9911, n9913, n9914, n9916, n9917, n9919, n9920, n9922, n9923,
    n9925, n9926, n9928, n9929, n9931, n9932, n9934, n9935, n9937, n9938,
    n9940, n9941, n9943, n9944, n9946, n9947, n9949, n9950, n9952, n9953,
    n9955, n9956, n9958, n9959, n9961, n9962, n9964, n9965, n9967, n9968,
    n9970, n9971, n9973, n9974, n9976, n9977, n9979, n9980, n9982, n9983,
    n9985, n9986, n9988, n9989, n9991, n9992, n9994, n9995, n9997, n9998,
    n10000, n10001, n10003, n10004, n10006, n10007, n10009, n10010, n10012,
    n10013, n10015, n10016, n10018, n10019, n10021, n10022, n10024, n10025,
    n10027, n10028, n10030, n10031, n10033, n10034, n10036, n10037, n10039,
    n10040, n10042, n10043, n10045, n10046, n10048, n10049, n10051, n10052,
    n10054, n10055, n10057, n10058, n10060, n10061, n10063, n10064, n10066,
    n10067, n10069, n10070, n10072, n10073, n10075, n10076, n10077, n10078,
    n10079, n10080, n10081, n10083, n10084, n10086, n10087, n10089, n10090,
    n10092, n10093, n10095, n10096, n10098, n10099, n10102, n10103, n10105,
    n10106, n10108, n10109, n10111, n10112, n10114, n10115, n10117, n10118,
    n10120, n10121, n10123, n10124, n10126, n10127, n10130, n10131, n10133,
    n10134, n10136, n10137, n10139, n10140, n10142, n10143, n10145, n10146,
    n10148, n10149, n10151, n10152, n10154, n10155, n10157, n10158, n10160,
    n10161, n10163, n10164, n10166, n10167, n10169, n10170, n10172, n10173,
    n10175, n10176, n10178, n10179, n10181, n10182, n10184, n10185, n10187,
    n10188, n10191, n10192, n10193, n10196, n10197, n10200;
  assign n2437 = ~pi0085 & ~pi0106;
  assign n2438 = n2437 & ~pi0076;
  assign n2439 = ~pi0048 & ~pi0061;
  assign n2440 = n2438 & n2439;
  assign n2441 = n2440 & ~pi0104;
  assign n2442 = n2441 & ~pi0089;
  assign n2443 = n2442 & ~pi0049;
  assign n2444 = n2443 & ~pi0045;
  assign n2445 = ~pi0073 & ~pi0084;
  assign n2446 = n2445 & ~pi0068;
  assign n2447 = n2446 & ~pi0066;
  assign n2448 = n2444 & n2447;
  assign n2449 = ~pi0069 & ~pi0083;
  assign n2450 = n2449 & ~pi0103;
  assign n2451 = n2448 & n2450;
  assign n2452 = ~pi0036 & ~pi0067;
  assign n2453 = pi0082 & pi0111;
  assign n2454 = n2452 & ~n2453;
  assign n2455 = ~pi0082 & ~pi0111;
  assign n2456 = pi0036 & pi0067;
  assign n2457 = n2455 & ~n2456;
  assign n2458 = ~n2454 & ~n2457;
  assign n2459 = n2451 & ~n2458;
  assign n2460 = n2455 & n2452;
  assign n2461 = n2450 & n2460;
  assign n2462 = ~n2459 & ~n2461;
  assign n2463 = ~n2440 & pi0104;
  assign n2464 = ~n2463 & ~pi0049;
  assign n2465 = ~n2442 & ~n2464;
  assign n2466 = ~n2441 & pi0089;
  assign n2467 = ~n2466 & ~pi0045;
  assign n2468 = ~n2465 & n2467;
  assign n2469 = ~n2468 & ~n2443;
  assign n2470 = ~n2437 & pi0076;
  assign n2471 = pi0085 & pi0106;
  assign n2472 = n2439 & ~n2471;
  assign n2473 = ~n2470 & n2472;
  assign n2474 = ~pi0048 ^ ~pi0061;
  assign n2475 = n2438 & n2474;
  assign n2476 = ~n2473 & ~n2475;
  assign n2477 = ~n2476 & n2447;
  assign n2478 = ~n2469 & n2477;
  assign n2479 = ~n2445 & pi0068;
  assign n2480 = ~n2447 & ~n2479;
  assign n2481 = pi0073 & pi0084;
  assign n2482 = ~n2481 & ~pi0066;
  assign n2483 = ~n2446 & ~n2482;
  assign n2484 = n2480 & ~n2483;
  assign n2485 = n2444 & n2484;
  assign n2486 = ~n2478 & ~n2485;
  assign n2487 = ~n2462 & ~n2486;
  assign n2488 = n2448 & n2460;
  assign n2489 = pi0069 ^ ~pi0083;
  assign n2490 = ~n2489 & ~pi0103;
  assign n2491 = ~n2490 & ~n2449;
  assign n2492 = n2488 & ~n2491;
  assign n2493 = ~n2487 & ~n2492;
  assign n2494 = n2455 & ~pi0036;
  assign n2495 = n2494 & ~pi0066;
  assign n2496 = n2495 & n2450;
  assign n2497 = n2444 & n2496;
  assign n2498 = n2497 & ~pi0073;
  assign n2499 = ~pi0088 & ~pi0098;
  assign n2500 = ~pi0102 & ~pi0107;
  assign n2501 = n2499 & n2500;
  assign n2502 = ~pi0064 & ~pi0065;
  assign n2503 = n2502 & ~pi0063;
  assign n2504 = n2501 & n2503;
  assign n2505 = n2504 & ~pi0081;
  assign n2506 = n2498 & n2505;
  assign n2507 = n2506 & n2488;
  assign n2508 = ~pi0071 & ~pi0081;
  assign n2509 = n2504 & n2508;
  assign n2510 = ~n2507 & ~n2509;
  assign n2511 = ~n2493 & ~n2510;
  assign n2512 = ~pi0067 & ~pi0068;
  assign n2513 = ~pi0071 & ~pi0084;
  assign n2514 = n2512 & n2513;
  assign n2515 = n2498 & n2514;
  assign n2516 = ~pi0102 ^ ~pi0107;
  assign n2517 = ~pi0088 ^ ~pi0098;
  assign n2518 = ~n2516 & ~n2517;
  assign n2519 = ~n2499 & ~n2500;
  assign n2520 = ~n2518 & ~n2519;
  assign n2521 = n2520 & ~pi0081;
  assign n2522 = n2501 & pi0081;
  assign n2523 = ~n2521 & ~n2522;
  assign n2524 = n2514 & ~pi0102;
  assign n2525 = n2499 & ~pi0081;
  assign n2526 = n2524 & n2525;
  assign n2527 = n2523 & n2526;
  assign n2528 = pi0064 & pi0065;
  assign n2529 = n2527 & ~n2528;
  assign n2530 = ~n2523 & n2502;
  assign n2531 = ~n2529 & ~n2530;
  assign n2532 = ~n2531 & ~pi0063;
  assign n2533 = n2527 & n2502;
  assign n2534 = ~n2532 & ~n2533;
  assign n2535 = n2515 & ~n2534;
  assign n2536 = ~n2511 & ~n2535;
  assign n2537 = ~pi0053 & ~pi0060;
  assign n2538 = n2537 & ~pi0050;
  assign n2539 = n2538 & ~pi0077;
  assign n2540 = ~pi0097 & ~pi0108;
  assign n2541 = n2539 & n2540;
  assign n2542 = ~pi0086 & ~pi0094;
  assign n2543 = n2541 & n2542;
  assign n2544 = ~n2536 & n2543;
  assign n2545 = n2506 & n2514;
  assign n2546 = pi0097 & pi0108;
  assign n2547 = n2542 & ~n2546;
  assign n2548 = ~n2541 & ~n2547;
  assign n2549 = ~n2539 & ~n2540;
  assign n2550 = ~n2548 & ~n2549;
  assign n2551 = n2545 & n2550;
  assign n2552 = ~n2544 & ~n2551;
  assign n2553 = pi0053 & pi0060;
  assign n2554 = ~n2553 & ~pi0077;
  assign n2555 = ~n2538 & ~n2554;
  assign n2556 = ~n2537 & pi0050;
  assign n2557 = ~pi0046 & ~pi0109;
  assign n2558 = ~n2556 & n2557;
  assign n2559 = ~n2555 & n2558;
  assign n2560 = ~n2552 & n2559;
  assign n2561 = pi0086 & pi0094;
  assign n2562 = n2560 & ~n2561;
  assign n2563 = n2545 & n2543;
  assign n2564 = n2562 & ~n2563;
  assign n2565 = ~pi0091 & ~pi0109;
  assign n2566 = ~n2565 & ~pi0046;
  assign n2567 = n2563 & n2566;
  assign n2568 = ~pi0058 & ~pi0090;
  assign n2569 = ~pi0047 & ~pi0110;
  assign n2570 = n2568 & n2569;
  assign n2571 = ~n2567 & n2570;
  assign n2572 = ~n2564 & n2571;
  assign n2573 = n2563 & n2559;
  assign n2574 = ~pi0091 & ~pi0093;
  assign n2575 = n2570 & n2574;
  assign n2576 = ~n2573 & ~n2575;
  assign n2577 = ~pi0047 ^ ~pi0091;
  assign n2578 = ~n2568 & n2577;
  assign n2579 = ~pi0035 & ~pi0093;
  assign n2580 = ~n2578 & n2579;
  assign n2581 = ~n2569 & pi0091;
  assign n2582 = n2580 & ~n2581;
  assign n2583 = n2568 & ~pi0047;
  assign n2584 = pi0058 & pi0090;
  assign n2585 = ~n2584 & ~pi0110;
  assign n2586 = ~n2583 & ~n2585;
  assign n2587 = n2582 & ~n2586;
  assign n2588 = ~n2576 & n2587;
  assign n2589 = ~n2572 & n2588;
  assign n2590 = ~pi0046 & ~pi0047;
  assign n2591 = n2565 & n2590;
  assign n2592 = ~pi0077 & ~pi0086;
  assign n2593 = ~pi0050 & ~pi0110;
  assign n2594 = n2592 & n2593;
  assign n2595 = n2591 & n2594;
  assign n2596 = n2537 & ~pi0058;
  assign n2597 = n2540 & ~pi0094;
  assign n2598 = n2596 & n2597;
  assign n2599 = n2595 & n2598;
  assign n2600 = n2545 & n2599;
  assign n2601 = n2600 & ~pi0090;
  assign n2602 = pi0035 ^ ~pi0093;
  assign n2603 = n2601 & ~n2602;
  assign n2604 = ~n2589 & ~n2603;
  assign n2605 = ~pi0072 & ~pi0096;
  assign n2606 = ~pi0051 & ~pi0070;
  assign n2607 = n2605 & n2606;
  assign n2608 = ~pi0032 & ~pi0095;
  assign n2609 = n2608 & ~pi0040;
  assign n2610 = n2607 & n2609;
  assign n2611 = ~n2604 & n2610;
  assign n2612 = n2579 & ~pi0090;
  assign n2613 = n2600 & n2612;
  assign n2614 = pi0051 & pi0070;
  assign n2615 = pi0072 & pi0096;
  assign n2616 = ~n2614 & ~n2615;
  assign n2617 = n2609 & n2616;
  assign n2618 = ~n2605 & ~n2606;
  assign n2619 = n2617 & ~n2618;
  assign n2620 = n2613 & n2619;
  assign n2621 = ~n2611 & ~n2620;
  assign n2622 = n2612 & n2607;
  assign n2623 = n2600 & n2622;
  assign n2624 = n2621 & ~n2623;
  assign n2625 = pi0040 ^ ~pi0095;
  assign n2626 = ~n2625 & ~pi0032;
  assign n2627 = pi0032 & ~pi0095;
  assign n2628 = n2627 & ~pi0040;
  assign n2629 = ~n2626 & ~n2628;
  assign n2630 = n2623 & n2629;
  assign n2631 = ~n2624 & ~n2630;
  assign n2632 = ~n2631 & ~n2610;
  assign n2633 = n2575 & pi0097;
  assign n2634 = n2560 & n2633;
  assign n2635 = n2610 & n2575;
  assign n2636 = n2635 & ~pi0035;
  assign n2637 = n2634 & n2636;
  assign n2638 = n2620 & pi0096;
  assign n2639 = ~n2637 & ~n2638;
  assign n2640 = pi1091 & pi1093;
  assign n2641 = ~pi0833 & pi0957;
  assign n2642 = n2640 & n2641;
  assign n2643 = ~pi1091 & pi1093;
  assign n2644 = ~n2642 & ~n2643;
  assign n2645 = pi0950 & pi1092;
  assign n2646 = n2645 & pi0829;
  assign po0840 = n2644 & n2646;
  assign n2648 = po0840 & ~pi0841;
  assign n2649 = n2600 & n2648;
  assign n2650 = po0840 & pi1093;
  assign n2651 = ~pi0046 & ~pi0094;
  assign n2652 = ~pi0036 ^ ~pi0097;
  assign n2653 = n2651 & n2652;
  assign n2654 = n2650 & n2653;
  assign n2655 = ~n2649 & ~n2654;
  assign n2656 = ~n2639 & ~n2655;
  assign n2657 = ~pi0174 & ~pi0189;
  assign n2658 = n2657 & ~pi0144;
  assign n2659 = ~pi0142 & ~pi0299;
  assign n2660 = ~n2658 & n2659;
  assign n2661 = ~pi0152 & ~pi0166;
  assign n2662 = n2661 & ~pi0161;
  assign n2663 = ~pi0146 & pi0299;
  assign n2664 = ~n2662 & n2663;
  assign n2665 = ~n2660 & ~n2664;
  assign n2666 = ~pi0198 & ~pi0299;
  assign n2667 = ~pi0210 & pi0299;
  assign n2668 = ~n2666 & ~n2667;
  assign n2669 = n2665 & ~n2668;
  assign n2670 = n2656 & n2669;
  assign n2671 = n2537 & ~pi0035;
  assign n2672 = ~n2671 & ~pi0097;
  assign n2673 = ~n2672 & ~pi0137;
  assign n2674 = ~n2670 & n2673;
  assign n2675 = n2573 & n2569;
  assign n2676 = ~pi0109 & ~pi0110;
  assign n2677 = ~n2590 & ~n2676;
  assign n2678 = n2563 & ~n2677;
  assign n2679 = ~n2675 & n2678;
  assign n2680 = ~n2679 & n2568;
  assign n2681 = ~n2680 & n2588;
  assign n2682 = ~pi0040 & ~pi0051;
  assign n2683 = n2605 & n2682;
  assign n2684 = n2683 & n2579;
  assign n2685 = ~pi0093 & pi0225;
  assign n2686 = ~n2685 & pi0035;
  assign n2687 = ~n2684 & ~n2686;
  assign n2688 = n2601 & n2687;
  assign n2689 = ~n2688 & ~pi0095;
  assign n2690 = ~n2681 & n2689;
  assign n2691 = ~n2589 & n2690;
  assign n2692 = ~n2674 & ~n2691;
  assign n2693 = ~n2632 & n2692;
  assign n2694 = pi0095 & ~pi0479;
  assign n2695 = ~n2638 & ~n2694;
  assign n2696 = ~n2693 & n2695;
  assign n2697 = ~n2695 & ~pi0234;
  assign n2698 = ~n2696 & ~n2697;
  assign n2699 = n2623 & ~pi0040;
  assign n2700 = n2699 & n2627;
  assign n2701 = ~n2668 & ~pi0841;
  assign n2702 = ~n2701 & pi0225;
  assign n2703 = n2700 & n2702;
  assign n2704 = ~n2698 & ~n2703;
  assign n2705 = n2631 & ~pi0228;
  assign n2706 = pi0105 & pi0228;
  assign n2707 = ~n2705 & ~n2706;
  assign n2708 = ~pi0216 & ~pi0221;
  assign n2709 = ~pi0215 & pi0299;
  assign n2710 = n2708 & n2709;
  assign n2711 = ~n2707 & n2710;
  assign n2712 = ~pi0223 & ~pi0224;
  assign n2713 = n2712 & ~pi0222;
  assign n2714 = n2713 & ~pi0299;
  assign n2715 = ~n2711 & ~n2714;
  assign n2716 = n2704 & ~n2715;
  assign n2717 = n2708 & ~pi0215;
  assign n2718 = ~n2707 & n2717;
  assign n2719 = ~pi0216 & pi0833;
  assign n2720 = n2719 & ~pi0929;
  assign n2721 = ~pi0221 & pi0265;
  assign n2722 = ~n2720 & ~n2721;
  assign n2723 = ~n2722 & ~pi0215;
  assign n2724 = ~n2719 & pi0221;
  assign n2725 = ~n2724 & ~pi0215;
  assign n2726 = ~n2725 & ~pi1144;
  assign n2727 = ~n2723 & ~n2726;
  assign n2728 = ~n2727 & ~pi0332;
  assign n2729 = ~n2728 & ~n2717;
  assign n2730 = ~n2729 & pi0299;
  assign n2731 = ~n2706 & pi0153;
  assign n2732 = n2731 & ~pi0332;
  assign n2733 = ~n2732 & n2717;
  assign n2734 = n2730 & ~n2733;
  assign n2735 = ~n2718 & n2734;
  assign n2736 = ~n2716 & ~n2735;
  assign n2737 = ~pi0075 & ~pi0100;
  assign n2738 = n2737 & ~pi0074;
  assign n2739 = ~pi0038 & ~pi0054;
  assign n2740 = n2738 & n2739;
  assign n2741 = ~pi0087 & ~pi0092;
  assign n2742 = n2741 & ~pi0039;
  assign n2743 = n2740 & n2742;
  assign n2744 = ~pi0056 & ~pi0062;
  assign n2745 = n2744 & ~pi0055;
  assign n2746 = ~pi0057 & ~pi0059;
  assign po1038 = ~n2745 | ~n2746;
  assign n2748 = n2743 & ~po1038;
  assign n2749 = ~n2736 & n2748;
  assign n2750 = n2623 & n2609;
  assign n2751 = n2750 & n2743;
  assign n2752 = pi0057 & ~pi0059;
  assign n2753 = n2744 & n2752;
  assign n2754 = n2751 & n2753;
  assign n2755 = ~pi0055 & n2754;
  assign n2756 = n2750 & ~po1038;
  assign n2757 = ~pi0074 & ~pi0092;
  assign n2758 = n2757 & ~pi0054;
  assign n2759 = n2737 & ~pi0087;
  assign n2760 = n2758 & n2759;
  assign n2761 = pi0038 & ~pi0039;
  assign n2762 = n2760 & n2761;
  assign n2763 = n2756 & n2762;
  assign n2764 = ~pi0039 & ~pi0087;
  assign n2765 = n2764 & ~pi0038;
  assign n2766 = n2737 & ~pi0092;
  assign n2767 = n2765 & n2766;
  assign n2768 = n2767 & ~pi0074;
  assign n2769 = n2744 & ~pi0057;
  assign n2770 = pi0054 & pi0059;
  assign n2771 = n2769 & ~n2770;
  assign n2772 = ~pi0054 & ~pi0059;
  assign n2773 = ~n2772 ^ ~pi0055;
  assign n2774 = n2771 & ~n2773;
  assign n2775 = n2768 & n2774;
  assign n2776 = n2750 & n2775;
  assign n2777 = ~n2763 & ~n2776;
  assign n2778 = ~n2755 & n2777;
  assign n2779 = n2756 & n2765;
  assign n2780 = ~pi0054 & ~pi0075;
  assign n2781 = ~pi0074 ^ ~pi0092;
  assign n2782 = n2780 & n2781;
  assign n2783 = pi0054 ^ ~pi0075;
  assign n2784 = n2757 & ~n2783;
  assign n2785 = ~n2782 & ~n2784;
  assign n2786 = n2779 & ~n2785;
  assign n2787 = n2786 & ~pi0100;
  assign n2788 = n2778 & ~n2787;
  assign n2789 = n2751 & n2746;
  assign n2790 = ~pi0056 ^ ~pi0062;
  assign n2791 = n2790 & ~pi0055;
  assign n2792 = n2789 & n2791;
  assign n2793 = ~pi0087 ^ ~pi0092;
  assign n2794 = ~pi0039 ^ ~pi0100;
  assign n2795 = ~n2793 & ~n2794;
  assign n2796 = ~pi0039 & ~pi0100;
  assign n2797 = ~n2741 & ~n2796;
  assign n2798 = ~n2795 & ~n2797;
  assign n2799 = ~pi0074 & ~pi0075;
  assign n2800 = n2799 & n2739;
  assign n2801 = n2798 & n2800;
  assign n2802 = n2756 & n2801;
  assign n2803 = ~n2792 & ~n2802;
  assign n2804 = n2788 & n2803;
  assign n2805 = ~n2804 & n2789;
  assign n2806 = n2805 & ~pi0228;
  assign n2807 = n2806 & n2717;
  assign n2808 = n2717 & ~n2731;
  assign n2809 = ~n2807 & ~n2808;
  assign n2810 = n2694 & pi0234;
  assign n2811 = ~n2810 & n2706;
  assign n2812 = ~n2805 & n2811;
  assign n2813 = ~n2812 & ~n2792;
  assign n2814 = ~n2809 & n2813;
  assign n2815 = ~pi0105 & pi0228;
  assign n2816 = ~n2815 & ~pi0137;
  assign n2817 = n2717 & ~n2816;
  assign n2818 = n2746 & ~pi0228;
  assign n2819 = n2731 & ~n2818;
  assign n2820 = n2817 & ~n2819;
  assign n2821 = ~n2804 & n2820;
  assign n2822 = ~n2729 & po1038;
  assign n2823 = ~n2821 & n2822;
  assign n2824 = ~n2814 & n2823;
  assign n2825 = n2740 & n2793;
  assign n2826 = ~pi0039 & pi0252;
  assign n2827 = ~n2825 & n2826;
  assign n2828 = ~n2662 & ~pi0146;
  assign n2829 = n2827 & ~n2828;
  assign n2830 = n2801 & ~pi0228;
  assign n2831 = ~n2829 & n2830;
  assign n2832 = n2750 & n2831;
  assign n2833 = n2832 & n2717;
  assign n2834 = n2710 & n2706;
  assign n2835 = ~n2714 & ~n2834;
  assign n2836 = ~n2810 & ~pi0332;
  assign n2837 = ~n2835 & n2836;
  assign n2838 = ~n2833 & ~n2837;
  assign n2839 = ~n2828 & ~pi0210;
  assign n2840 = ~pi0137 & ~pi0332;
  assign n2841 = ~n2839 & n2840;
  assign n2842 = n2730 & n2841;
  assign n2843 = n2714 & n2840;
  assign n2844 = ~n2658 & ~pi0142;
  assign n2845 = ~n2844 & ~pi0198;
  assign n2846 = n2843 & ~n2845;
  assign n2847 = pi0075 ^ ~pi0100;
  assign n2848 = n2758 & ~n2847;
  assign n2849 = ~n2846 & n2848;
  assign n2850 = n2737 & pi0137;
  assign n2851 = ~n2785 & n2850;
  assign n2852 = ~n2849 & ~n2851;
  assign n2853 = ~n2842 & ~n2852;
  assign n2854 = n2750 & n2853;
  assign n2855 = n2854 & n2765;
  assign n2856 = ~n2838 & ~n2855;
  assign n2857 = ~n2833 & n2734;
  assign n2858 = ~n2856 & ~n2857;
  assign n2859 = ~n2734 & n2760;
  assign n2860 = ~n2859 & ~n2825;
  assign n2861 = ~n2860 & ~pi0039;
  assign n2862 = n2739 & n2757;
  assign n2863 = n2759 & n2862;
  assign n2864 = ~n2861 & ~n2863;
  assign n2865 = n2815 & pi0153;
  assign n2866 = n2817 & ~n2865;
  assign n2867 = ~n2866 & ~pi0332;
  assign n2868 = n2730 & n2867;
  assign n2869 = ~n2868 & ~n2843;
  assign n2870 = ~n2864 & n2869;
  assign n2871 = n2750 & n2870;
  assign n2872 = ~n2743 & ~po1038;
  assign n2873 = ~n2871 & n2872;
  assign n2874 = ~n2858 & n2873;
  assign n2875 = ~pi0224 & pi0833;
  assign n2876 = ~n2875 & pi0222;
  assign n2877 = ~n2876 & ~pi0223;
  assign n2878 = ~n2877 & pi1144;
  assign n2879 = n2875 & pi0929;
  assign n2880 = pi0224 & pi0265;
  assign n2881 = ~n2880 & ~pi0222;
  assign n2882 = ~n2879 & ~n2881;
  assign n2883 = ~n2882 & ~pi0223;
  assign n2884 = ~n2878 & ~n2883;
  assign n2885 = ~po1038 & ~pi0299;
  assign n2886 = n2884 & n2885;
  assign n2887 = ~n2874 & ~n2886;
  assign n2888 = ~n2824 & n2887;
  assign n2889 = ~n2749 & n2888;
  assign po0153 = n2889 | pi0332;
  assign n2891 = n2631 & n2748;
  assign n2892 = ~n2891 & ~n2805;
  assign n2893 = ~n2892 & ~pi0228;
  assign n2894 = n2832 & ~po1038;
  assign n2895 = ~n2893 & ~n2894;
  assign n2896 = ~n2895 & n2717;
  assign n2897 = ~n2896 & ~n2885;
  assign n2898 = n2717 & ~n2706;
  assign n2899 = n2898 & ~pi0154;
  assign n2900 = ~pi0215 & pi0221;
  assign n2901 = n2719 & n2900;
  assign n2902 = n2901 & pi0939;
  assign n2903 = pi0216 & ~pi0221;
  assign n2904 = n2903 & ~pi0215;
  assign n2905 = n2904 & pi0276;
  assign n2906 = ~n2902 & ~n2905;
  assign n2907 = ~n2899 & n2906;
  assign n2908 = ~n2725 & pi1146;
  assign n2909 = n2907 & ~n2908;
  assign n2910 = n2717 & n2706;
  assign n2911 = n2910 & n2694;
  assign n2912 = n2911 & pi0239;
  assign n2913 = n2909 & ~n2912;
  assign n2914 = n2897 & ~n2913;
  assign n2915 = n2743 & n2717;
  assign n2916 = n2915 & pi0299;
  assign n2917 = ~n2695 & n2916;
  assign n2918 = n2705 & n2917;
  assign n2919 = ~n2743 & ~n2694;
  assign n2920 = ~n2695 & ~n2919;
  assign n2921 = n2920 & ~n2835;
  assign n2922 = ~n2918 & ~n2921;
  assign n2923 = ~n2922 & pi0239;
  assign n2924 = ~n2877 & ~pi0299;
  assign n2925 = n2924 & pi1146;
  assign n2926 = ~pi0223 & ~pi0299;
  assign n2927 = n2926 & pi0222;
  assign n2928 = n2927 & n2875;
  assign n2929 = n2928 & pi0939;
  assign n2930 = n2926 & pi0224;
  assign n2931 = n2930 & ~pi0222;
  assign n2932 = n2931 & pi0276;
  assign n2933 = ~n2929 & ~n2932;
  assign n2934 = ~n2925 & n2933;
  assign n2935 = ~n2923 & n2934;
  assign n2936 = ~n2935 & ~po1038;
  assign po0154 = n2914 | n2936;
  assign n2938 = ~n2706 & ~pi0151;
  assign n2939 = n2717 & ~n2938;
  assign n2940 = n2904 & pi0274;
  assign n2941 = ~n2939 & ~n2940;
  assign n2942 = n2901 & ~pi0927;
  assign n2943 = n2941 & ~n2942;
  assign n2944 = ~n2725 & ~pi1145;
  assign n2945 = n2943 & ~n2944;
  assign n2946 = n2911 & pi0235;
  assign n2947 = ~n2945 & ~n2946;
  assign n2948 = n2897 & ~n2947;
  assign n2949 = ~n2922 & pi0235;
  assign n2950 = n2924 & pi1145;
  assign n2951 = n2931 & ~pi0274;
  assign n2952 = n2928 & pi0927;
  assign n2953 = ~n2951 & ~n2952;
  assign n2954 = ~n2950 & n2953;
  assign n2955 = ~n2949 & n2954;
  assign n2956 = ~n2955 & ~po1038;
  assign po0155 = n2948 | n2956;
  assign n2958 = n2707 & pi0146;
  assign n2959 = n2695 & pi0284;
  assign n2960 = ~n2707 & ~n2959;
  assign n2961 = ~n2958 & ~n2960;
  assign n2962 = ~n2961 & n2915;
  assign n2963 = n2910 & ~n2694;
  assign n2964 = n2963 & ~pi0284;
  assign n2965 = n2904 & ~pi0264;
  assign n2966 = n2901 & pi0944;
  assign n2967 = ~n2965 & ~n2966;
  assign n2968 = ~n2964 & n2967;
  assign n2969 = n2898 & pi0146;
  assign n2970 = ~n2725 & pi1143;
  assign n2971 = ~n2969 & ~n2970;
  assign n2972 = n2968 & n2971;
  assign n2973 = ~n2833 & ~n2972;
  assign n2974 = ~n2973 & pi0299;
  assign n2975 = ~n2832 & ~n2706;
  assign n2976 = ~n2694 & pi0284;
  assign n2977 = n2717 & ~n2976;
  assign n2978 = n2977 & ~n2815;
  assign n2979 = ~n2975 & n2978;
  assign n2980 = n2974 & ~n2979;
  assign n2981 = ~n2980 & ~n2916;
  assign n2982 = ~n2962 & ~n2981;
  assign n2983 = ~n2922 & ~pi0238;
  assign n2984 = n2714 & pi0284;
  assign n2985 = ~n2920 & n2984;
  assign n2986 = n2931 & pi0264;
  assign n2987 = ~n2986 & ~po1038;
  assign n2988 = n2928 & ~pi0944;
  assign n2989 = n2987 & ~n2988;
  assign n2990 = n2924 & ~pi1143;
  assign n2991 = n2989 & ~n2990;
  assign n2992 = ~n2985 & n2991;
  assign n2993 = ~n2983 & n2992;
  assign n2994 = ~n2982 & n2993;
  assign n2995 = pi0228 & pi0238;
  assign n2996 = ~n2807 & ~n2995;
  assign n2997 = ~n2996 & n2978;
  assign n2998 = ~n2807 & ~n2972;
  assign n2999 = ~n2997 & ~n2998;
  assign n3000 = ~n2999 & po1038;
  assign po0156 = n2994 | n3000;
  assign n3002 = ~n2806 & ~n2706;
  assign n3003 = n3002 & ~n2894;
  assign n3004 = ~n3003 & ~pi0262;
  assign n3005 = n3002 & ~pi0172;
  assign n3006 = n2706 & n2694;
  assign n3007 = ~n3005 & ~n3006;
  assign n3008 = ~n3004 & n3007;
  assign n3009 = ~n3008 & n2717;
  assign n3010 = ~n2719 & ~pi1142;
  assign n3011 = ~n3010 & pi0221;
  assign n3012 = n2719 & ~pi0932;
  assign n3013 = n3011 & ~n3012;
  assign n3014 = n2903 & ~pi0277;
  assign n3015 = ~n3013 & ~n3014;
  assign n3016 = ~n3015 & ~pi0215;
  assign n3017 = pi0215 & pi1142;
  assign n3018 = ~n3016 & ~n3017;
  assign n3019 = ~n3009 & n3018;
  assign n3020 = ~po1038 & pi0262;
  assign n3021 = n2833 & n3020;
  assign n3022 = n2694 & ~pi0249;
  assign n3023 = n2910 & n3022;
  assign n3024 = ~n2885 & ~n3023;
  assign n3025 = ~n3021 & n3024;
  assign n3026 = ~n3019 & n3025;
  assign n3027 = ~n2920 & pi0262;
  assign n3028 = n2714 & ~n3022;
  assign n3029 = ~n3027 & n3028;
  assign n3030 = n2924 & pi1142;
  assign n3031 = n2931 & ~pi0277;
  assign n3032 = n2928 & pi0932;
  assign n3033 = ~n3031 & ~n3032;
  assign n3034 = ~n3030 & n3033;
  assign n3035 = ~n3029 & n3034;
  assign n3036 = ~n3035 & ~po1038;
  assign n3037 = ~n3026 & ~n3036;
  assign n3038 = ~n2695 & ~pi0249;
  assign n3039 = n3038 & n2714;
  assign n3040 = n3015 & n2709;
  assign n3041 = ~n3039 & ~n3040;
  assign n3042 = ~n3041 & n2748;
  assign n3043 = ~n3037 & ~n3042;
  assign n3044 = n2707 & pi0172;
  assign n3045 = n3042 & n2710;
  assign n3046 = ~n3044 & n3045;
  assign n3047 = n2695 & pi0262;
  assign n3048 = ~n3038 & ~n3047;
  assign n3049 = ~n2707 & ~n3048;
  assign n3050 = n3046 & ~n3049;
  assign po0157 = n3043 | n3050;
  assign n3052 = n2898 & pi0171;
  assign n3053 = ~n2694 & pi0861;
  assign n3054 = n2910 & ~n3053;
  assign n3055 = ~n3052 & ~n3054;
  assign n3056 = n2901 & ~pi0935;
  assign n3057 = n2904 & pi0270;
  assign n3058 = ~n3056 & ~n3057;
  assign n3059 = ~n2725 & ~pi1141;
  assign n3060 = n3058 & ~n3059;
  assign n3061 = n3055 & n3060;
  assign n3062 = ~n2718 & ~n3061;
  assign n3063 = ~n3062 & n2743;
  assign n3064 = ~n3063 & pi0299;
  assign n3065 = ~n2638 & n3053;
  assign n3066 = ~n2715 & ~n3065;
  assign n3067 = ~n3064 & ~n3066;
  assign n3068 = n2833 & pi0861;
  assign n3069 = ~n2833 & n3061;
  assign n3070 = ~n3068 & ~n3069;
  assign n3071 = n3070 & pi0299;
  assign n3072 = ~n3053 & ~pi0299;
  assign n3073 = ~n2743 & ~n3072;
  assign n3074 = ~n3071 & n3073;
  assign n3075 = ~n3067 & ~n3074;
  assign n3076 = n2924 & ~pi1141;
  assign n3077 = n2928 & ~pi0935;
  assign n3078 = n2931 & pi0270;
  assign n3079 = ~n3077 & ~n3078;
  assign n3080 = ~n3076 & n3079;
  assign n3081 = ~n3075 & n3080;
  assign n3082 = ~n2922 & pi0241;
  assign n3083 = ~n3082 & ~po1038;
  assign n3084 = ~n3081 & n3083;
  assign n3085 = ~n2807 & n3061;
  assign n3086 = ~n2911 & po1038;
  assign n3087 = po1038 & ~pi0241;
  assign n3088 = ~n3086 & ~n3087;
  assign n3089 = ~n3085 & ~n3088;
  assign n3090 = n2807 & pi0861;
  assign n3091 = n3089 & ~n3090;
  assign po0158 = ~n3084 & ~n3091;
  assign n3093 = n2705 & n2743;
  assign n3094 = ~n3093 & n2975;
  assign n3095 = ~n3094 & pi0869;
  assign n3096 = ~n3095 & n2717;
  assign n3097 = n3094 & ~pi0170;
  assign n3098 = n3096 & ~n3097;
  assign n3099 = ~n2725 & pi1140;
  assign n3100 = n2719 & pi0921;
  assign n3101 = pi0216 & pi0282;
  assign n3102 = ~n3101 & ~pi0221;
  assign n3103 = ~n3100 & ~n3102;
  assign n3104 = ~n3103 & ~pi0215;
  assign n3105 = ~n3099 & ~n3104;
  assign n3106 = ~n3105 & pi0299;
  assign n3107 = ~n3098 & n3106;
  assign n3108 = n2924 & pi1140;
  assign n3109 = ~n2694 & pi0869;
  assign n3110 = n2714 & n3109;
  assign n3111 = ~n3108 & ~n3110;
  assign n3112 = n2928 & pi0921;
  assign n3113 = n2931 & ~pi0282;
  assign n3114 = ~n3112 & ~n3113;
  assign n3115 = n3111 & n3114;
  assign n3116 = ~n3107 & n3115;
  assign n3117 = n2922 & ~po1038;
  assign n3118 = ~n3116 & n3117;
  assign n3119 = ~n3086 & pi0248;
  assign n3120 = ~n3117 & n3119;
  assign n3121 = ~n2807 & ~n2963;
  assign n3122 = ~n3121 & pi0869;
  assign n3123 = ~n2706 & ~pi0170;
  assign n3124 = n2717 & ~n3123;
  assign n3125 = ~n3105 & ~n3124;
  assign n3126 = ~n2807 & n3125;
  assign n3127 = ~n3122 & ~n3126;
  assign n3128 = ~n3127 & po1038;
  assign n3129 = ~n3120 & ~n3128;
  assign po0159 = n3118 | ~n3129;
  assign n3131 = n2707 & ~pi0148;
  assign n3132 = ~n3131 & n2916;
  assign n3133 = n2695 & pi0862;
  assign n3134 = ~n2695 & pi0247;
  assign n3135 = ~n3133 & ~n3134;
  assign n3136 = ~n2707 & ~n3135;
  assign n3137 = n3132 & ~n3136;
  assign n3138 = n2920 & pi0247;
  assign n3139 = ~n2920 & pi0862;
  assign n3140 = ~n3138 & ~n3139;
  assign n3141 = n3140 & n2714;
  assign n3142 = n2898 & pi0148;
  assign n3143 = n2901 & ~pi0920;
  assign n3144 = ~n3142 & ~n3143;
  assign n3145 = ~n2725 & ~pi1139;
  assign n3146 = n2904 & pi0281;
  assign n3147 = ~n3145 & ~n3146;
  assign n3148 = n3144 & n3147;
  assign n3149 = n2963 & ~pi0862;
  assign n3150 = n2911 & ~pi0247;
  assign n3151 = ~n3149 & ~n3150;
  assign n3152 = n3148 & n3151;
  assign n3153 = ~n3152 & ~n2915;
  assign n3154 = ~n2833 & n3153;
  assign n3155 = n2833 & ~pi0862;
  assign n3156 = ~n3154 & ~n3155;
  assign n3157 = ~n3156 & pi0299;
  assign n3158 = n2931 & pi0281;
  assign n3159 = ~n3158 & ~po1038;
  assign n3160 = n2928 & ~pi0920;
  assign n3161 = n3159 & ~n3160;
  assign n3162 = n2924 & ~pi1139;
  assign n3163 = n3161 & ~n3162;
  assign n3164 = ~n3157 & n3163;
  assign n3165 = ~n3141 & n3164;
  assign n3166 = ~n3137 & n3165;
  assign n3167 = ~n2807 & ~n3152;
  assign n3168 = ~n3167 & po1038;
  assign n3169 = n2807 & ~pi0862;
  assign n3170 = n3168 & ~n3169;
  assign po0160 = n3166 | n3170;
  assign n3172 = n2695 & ~pi0877;
  assign n3173 = ~n2695 & ~pi0246;
  assign n3174 = ~n3172 & ~n3173;
  assign n3175 = ~n2707 & ~n3174;
  assign n3176 = n2707 & pi0169;
  assign n3177 = ~n3175 & ~n3176;
  assign n3178 = n3177 & n2743;
  assign n3179 = n2975 & ~pi0169;
  assign n3180 = ~n2694 & pi0877;
  assign n3181 = ~n2975 & n3180;
  assign n3182 = ~n3179 & ~n3181;
  assign n3183 = n3182 & n2717;
  assign n3184 = ~n3183 & ~n2915;
  assign n3185 = ~n3178 & ~n3184;
  assign n3186 = ~n2725 & ~pi1138;
  assign n3187 = n2904 & pi0269;
  assign n3188 = n2901 & ~pi0940;
  assign n3189 = ~n3187 & ~n3188;
  assign n3190 = ~n3186 & n3189;
  assign n3191 = n3190 & pi0299;
  assign n3192 = ~n3185 & n3191;
  assign n3193 = n2921 & ~pi0246;
  assign n3194 = n2924 & pi1138;
  assign n3195 = n2931 & ~pi0269;
  assign n3196 = n2714 & pi0877;
  assign n3197 = ~n3195 & ~n3196;
  assign n3198 = ~n3194 & n3197;
  assign n3199 = n2928 & pi0940;
  assign n3200 = n3198 & ~n3199;
  assign n3201 = ~n2921 & n3200;
  assign n3202 = ~n3193 & ~n3201;
  assign n3203 = ~n3202 & ~po1038;
  assign n3204 = ~n3192 & n3203;
  assign n3205 = ~n3002 & n3180;
  assign n3206 = ~n3205 & n2717;
  assign n3207 = n3002 & ~pi0169;
  assign n3208 = n3206 & ~n3207;
  assign n3209 = ~n3208 & n3190;
  assign n3210 = n2911 & pi0246;
  assign n3211 = ~n3210 & po1038;
  assign n3212 = ~n3209 & n3211;
  assign po0161 = ~n3204 & ~n3212;
  assign n3214 = ~n2695 & ~pi0240;
  assign n3215 = n2695 & ~pi0878;
  assign n3216 = ~n3214 & ~n3215;
  assign n3217 = ~n2707 & ~n3216;
  assign n3218 = ~n2706 & pi0168;
  assign n3219 = ~n2705 & n3218;
  assign n3220 = ~n2921 & ~n2743;
  assign n3221 = ~n3220 & n2710;
  assign n3222 = ~n3219 & n3221;
  assign n3223 = ~n3217 & n3222;
  assign n3224 = ~n2694 & pi0878;
  assign n3225 = ~n3224 & n2706;
  assign n3226 = n2717 & ~n3218;
  assign n3227 = ~n3225 & n3226;
  assign n3228 = n2904 & ~pi0280;
  assign n3229 = ~n3227 & ~n3228;
  assign n3230 = ~n2833 & ~n3229;
  assign n3231 = ~n2725 & pi1137;
  assign n3232 = n2901 & pi0933;
  assign n3233 = ~n3231 & ~n3232;
  assign n3234 = n3233 & pi0299;
  assign n3235 = ~n3230 & n3234;
  assign n3236 = n2833 & pi0878;
  assign n3237 = n3235 & ~n3236;
  assign n3238 = n2921 & n2743;
  assign n3239 = ~n3237 & ~n3238;
  assign n3240 = n3239 & ~n2916;
  assign n3241 = ~n3223 & ~n3240;
  assign n3242 = n2924 & ~pi1137;
  assign n3243 = n2714 & ~n3224;
  assign n3244 = n2931 & pi0280;
  assign n3245 = ~n3243 & ~n3244;
  assign n3246 = ~n3242 & n3245;
  assign n3247 = n2928 & ~pi0933;
  assign n3248 = n3246 & ~n3247;
  assign n3249 = ~n3241 & n3248;
  assign n3250 = n2714 & pi0240;
  assign n3251 = n2920 & n3250;
  assign n3252 = ~n3251 & ~po1038;
  assign n3253 = ~n3249 & n3252;
  assign n3254 = n2911 & pi0240;
  assign n3255 = n3233 & ~n3254;
  assign n3256 = n3255 & n3229;
  assign n3257 = ~n2807 & ~n3256;
  assign n3258 = ~n3257 & po1038;
  assign n3259 = n2807 & pi0878;
  assign n3260 = n3258 & ~n3259;
  assign po0162 = ~n3253 & ~n3260;
  assign n3262 = n2707 & ~po1038;
  assign n3263 = n2975 & pi0166;
  assign n3264 = ~n2694 & pi0875;
  assign n3265 = ~n2975 & n3264;
  assign n3266 = ~n3263 & ~n3265;
  assign n3267 = n3262 & n3266;
  assign n3268 = ~n3267 & n2717;
  assign n3269 = n3002 & pi0166;
  assign n3270 = ~n2694 & ~pi0875;
  assign n3271 = ~n3002 & ~n3270;
  assign n3272 = ~n3269 & ~n3271;
  assign n3273 = n3272 & ~n2748;
  assign n3274 = ~n3262 & n3273;
  assign n3275 = ~n3266 & ~n2748;
  assign n3276 = ~n2695 & ~pi0245;
  assign n3277 = n2695 & ~pi0875;
  assign n3278 = ~n3276 & ~n3277;
  assign n3279 = ~n3275 & ~n3278;
  assign n3280 = ~n2707 & n3279;
  assign n3281 = ~n3274 & ~n3280;
  assign n3282 = n3268 & n3281;
  assign n3283 = ~n2725 & pi1136;
  assign n3284 = n2901 & pi0928;
  assign n3285 = n2904 & pi0266;
  assign n3286 = ~n3284 & ~n3285;
  assign n3287 = ~n3283 & n3286;
  assign n3288 = n3287 & ~n2885;
  assign n3289 = ~n3282 & n3288;
  assign n3290 = n2920 & pi0245;
  assign n3291 = ~po1038 & n2714;
  assign n3292 = ~n3290 & n3291;
  assign n3293 = ~n2920 & pi0875;
  assign n3294 = n3292 & ~n3293;
  assign n3295 = n2924 & ~pi1136;
  assign n3296 = n2931 & ~pi0266;
  assign n3297 = n2928 & ~pi0928;
  assign n3298 = ~n3296 & ~n3297;
  assign n3299 = ~n3295 & n3298;
  assign n3300 = ~n3299 & ~po1038;
  assign n3301 = ~n3294 & ~n3300;
  assign po0163 = ~n3289 & n3301;
  assign n3303 = n3094 & ~pi0161;
  assign n3304 = ~n3303 & n2717;
  assign n3305 = ~n2920 & pi0879;
  assign n3306 = ~n3094 & ~n3305;
  assign n3307 = n3304 & ~n3306;
  assign n3308 = ~n2922 & pi0244;
  assign n3309 = ~n2975 & n2710;
  assign n3310 = ~n3309 & ~n2714;
  assign n3311 = n3305 & ~n3310;
  assign n3312 = n2931 & pi0279;
  assign n3313 = ~n3312 & ~po1038;
  assign n3314 = n2928 & pi0938;
  assign n3315 = n3313 & ~n3314;
  assign n3316 = n2924 & pi1135;
  assign n3317 = n3315 & ~n3316;
  assign n3318 = ~n3311 & n3317;
  assign n3319 = ~n3308 & n3318;
  assign n3320 = ~n3307 & n3319;
  assign n3321 = n3002 & ~pi0161;
  assign n3322 = ~n2694 & pi0879;
  assign n3323 = n2694 & pi0244;
  assign n3324 = ~n3322 & ~n3323;
  assign n3325 = ~n3002 & n3324;
  assign n3326 = ~n3321 & ~n3325;
  assign n3327 = n3326 & n2717;
  assign n3328 = ~n3327 & po1038;
  assign n3329 = ~n3320 & ~n3328;
  assign n3330 = ~n2725 & pi1135;
  assign n3331 = n2901 & pi0938;
  assign n3332 = n2904 & pi0279;
  assign n3333 = ~n3331 & ~n3332;
  assign n3334 = ~n3330 & n3333;
  assign n3335 = ~n3329 & n3334;
  assign n3336 = n3319 & ~pi0299;
  assign po0164 = ~n3335 & ~n3336;
  assign n3338 = n3094 & pi0152;
  assign n3339 = ~n3338 & n2717;
  assign n3340 = ~n2920 & pi0846;
  assign n3341 = n2920 & pi0242;
  assign n3342 = ~n3340 & ~n3341;
  assign n3343 = ~n3094 & ~n3342;
  assign n3344 = n3339 & ~n3343;
  assign n3345 = n3342 & n2714;
  assign n3346 = n2928 & ~pi0930;
  assign n3347 = n2931 & ~pi0278;
  assign n3348 = ~n3346 & ~n3347;
  assign n3349 = n3348 & ~po1038;
  assign n3350 = ~n3345 & n3349;
  assign n3351 = ~n3344 & n3350;
  assign n3352 = ~n2694 & pi0846;
  assign n3353 = n2694 & pi0242;
  assign n3354 = ~n3352 & ~n3353;
  assign n3355 = ~n3002 & ~n3354;
  assign n3356 = ~n3355 & n2717;
  assign n3357 = n3002 & pi0152;
  assign n3358 = n3356 & ~n3357;
  assign n3359 = ~n3358 & po1038;
  assign n3360 = ~n3351 & ~n3359;
  assign n3361 = n2904 & ~pi0278;
  assign n3362 = n2901 & ~pi0930;
  assign n3363 = ~n3361 & ~n3362;
  assign n3364 = ~n3360 & n3363;
  assign n3365 = n3350 & ~pi0299;
  assign n3366 = ~n3364 & ~n3365;
  assign n3367 = n2885 & ~n2924;
  assign n3368 = ~n2885 & n2725;
  assign n3369 = ~n3367 & ~n3368;
  assign n3370 = n3369 & ~pi1134;
  assign po0165 = ~n3366 & ~n3370;
  assign n3372 = n2545 & n2597;
  assign n3373 = n2588 & ~n3372;
  assign n3374 = n2562 & n3373;
  assign n3375 = pi0093 & pi0841;
  assign n3376 = n2603 & ~n3375;
  assign n3377 = ~n3376 & n2683;
  assign n3378 = ~n2681 & n3377;
  assign n3379 = ~n3374 & n3378;
  assign n3380 = ~n2632 & ~n3379;
  assign n3381 = ~n3380 & ~n2699;
  assign n3382 = n2699 & ~n2701;
  assign n3383 = ~n3382 & pi0032;
  assign n3384 = ~pi0070 & ~pi0095;
  assign n3385 = n2537 & n3384;
  assign n3386 = ~n3383 & n3385;
  assign n3387 = ~n3386 & pi0032;
  assign n3388 = ~n2750 & n2748;
  assign n3389 = ~n3387 & n3388;
  assign n3390 = ~n3381 & n3389;
  assign n3391 = ~pi0614 & ~pi0616;
  assign n3392 = n3391 & ~pi0642;
  assign n3393 = n3392 & pi0603;
  assign n3394 = ~pi0661 & ~pi0662;
  assign n3395 = n3394 & ~pi0681;
  assign n3396 = n3395 & pi0680;
  assign po1101 = n3393 | n3396;
  assign n3398 = ~pi0332 & ~pi0468;
  assign n3399 = ~po1101 & ~n3398;
  assign n3400 = ~pi0969 & ~pi0971;
  assign n3401 = ~pi0974 & ~pi0977;
  assign n3402 = n3400 & n3401;
  assign n3403 = ~pi0587 & ~pi0602;
  assign n3404 = ~pi0961 & ~pi0967;
  assign n3405 = n3403 & n3404;
  assign n3406 = n3402 & n3405;
  assign n3407 = n3406 & n3398;
  assign n3408 = ~n3399 & ~n3407;
  assign n3409 = n3398 & pi0299;
  assign n3410 = ~n3408 & ~n3409;
  assign n3411 = n2645 & pi0824;
  assign n3412 = ~n2642 & n3411;
  assign po0950 = ~po0840 & ~n3412;
  assign n3414 = ~n3410 & ~po0950;
  assign n3415 = ~pi0979 & ~pi0984;
  assign n3416 = n3415 & ~pi0287;
  assign n3417 = ~pi0252 & ~pi1001;
  assign n3418 = ~n3417 & pi0835;
  assign n3419 = n3416 & n3418;
  assign n3420 = n3414 & n3419;
  assign n3421 = ~n2709 & ~n2926;
  assign n3422 = n3420 & n3421;
  assign n3423 = ~pi0970 & ~pi0972;
  assign n3424 = ~pi0975 & ~pi0978;
  assign n3425 = n3423 & n3424;
  assign n3426 = ~pi0907 & ~pi0947;
  assign n3427 = ~pi0960 & ~pi0963;
  assign n3428 = n3426 & n3427;
  assign n3429 = n3425 & n3428;
  assign n3430 = n3429 & n3398;
  assign n3431 = n3430 & pi0299;
  assign n3432 = n3422 & ~n3431;
  assign n3433 = n3432 & pi0039;
  assign n3434 = ~pi0041 & ~pi0101;
  assign n3435 = n3434 & ~pi0099;
  assign n3436 = n3435 & ~pi0113;
  assign n3437 = ~pi0043 & ~pi0044;
  assign n3438 = ~pi0042 & ~pi0114;
  assign n3439 = n3437 & n3438;
  assign n3440 = ~pi0115 & ~pi0116;
  assign n3441 = n3439 & n3440;
  assign n3442 = n3436 & n3441;
  assign po1057 = ~n3442 | pi0052;
  assign n3444 = ~pi0129 & pi0250;
  assign n3445 = ~n3444 & pi0683;
  assign n3446 = po1057 & n3445;
  assign n3447 = ~n3446 & ~n2665;
  assign n3448 = ~n2665 & ~pi0250;
  assign n3449 = n3411 & ~pi1093;
  assign n3450 = n2646 & ~pi1093;
  assign po0740 = n3449 | n3450;
  assign n3452 = n3448 & po0740;
  assign n3453 = n2665 & ~pi0252;
  assign n3454 = ~n3452 & ~n3453;
  assign n3455 = ~n3447 & n3454;
  assign n3456 = ~n3455 & pi0100;
  assign n3457 = ~pi0087 & pi0100;
  assign n3458 = ~n2765 & ~n3457;
  assign n3459 = ~n3458 & ~pi0074;
  assign n3460 = ~n3456 & n3459;
  assign n3461 = n2927 & pi0224;
  assign n3462 = n3408 & n3461;
  assign n3463 = ~n3399 & ~n3430;
  assign n3464 = n2900 & pi0299;
  assign n3465 = n3464 & pi0216;
  assign n3466 = n3463 & n3465;
  assign n3467 = ~n3462 & ~n3466;
  assign n3468 = n2650 & n3419;
  assign n3469 = ~n3467 & n3468;
  assign n3470 = n3469 & pi0039;
  assign n3471 = ~n3460 & ~n3470;
  assign n3472 = ~n3433 & n3471;
  assign n3473 = ~n2804 & n3472;
  assign n3474 = ~n2755 & ~n2792;
  assign n3475 = ~n3473 & n3474;
  assign po0167 = n3390 | ~n3475;
  assign n3477 = n2748 & n2610;
  assign n3478 = n2681 & n3477;
  assign n3479 = ~n2891 & ~n3478;
  assign n3480 = ~n2449 & pi0067;
  assign n3481 = n2494 & ~n3480;
  assign n3482 = n2489 & ~pi0067;
  assign n3483 = n3481 & ~n3482;
  assign n3484 = n2448 & n3483;
  assign n3485 = n2508 & ~pi0085;
  assign n3486 = ~n2485 & n3485;
  assign n3487 = ~n3484 & n3486;
  assign n3488 = n3487 & ~pi0082;
  assign n3489 = ~n3372 & n3488;
  assign n3490 = n2569 & ~pi0058;
  assign n3491 = ~n3489 & n3490;
  assign n3492 = n3377 & n3491;
  assign n3493 = pi0103 & ~pi0314;
  assign n3494 = ~n3493 & ~pi0109;
  assign n3495 = ~n3492 & n3494;
  assign n3496 = ~n3479 & ~n3495;
  assign n3497 = ~n3496 & ~pi0072;
  assign n3498 = ~n2621 & n2748;
  assign n3499 = n2700 & n2701;
  assign n3500 = n2526 & n2502;
  assign n3501 = n3500 & n2599;
  assign n3502 = n2497 & n3501;
  assign n3503 = n2622 & ~pi0073;
  assign n3504 = n3502 & n3503;
  assign n3505 = n2694 & ~pi0032;
  assign n3506 = n3504 & n3505;
  assign n3507 = n2607 & n2608;
  assign n3508 = ~pi0058 & pi0841;
  assign n3509 = ~pi0058 ^ ~pi0090;
  assign n3510 = ~n3508 & n3509;
  assign n3511 = n3507 & n3510;
  assign n3512 = ~n3506 & ~n3511;
  assign n3513 = ~n3499 & n3512;
  assign n3514 = n3513 & ~n2609;
  assign n3515 = n2748 & n2607;
  assign n3516 = n2588 & n3515;
  assign n3517 = ~n3514 & n3516;
  assign n3518 = ~n3498 & ~n3517;
  assign n3519 = ~n3497 & ~n3518;
  assign n3520 = pi0158 & pi0159;
  assign n3521 = n3520 & pi0197;
  assign n3522 = pi0160 & pi0232;
  assign n3523 = n3521 & n3522;
  assign n3524 = ~n3523 & pi0299;
  assign n3525 = ~n3524 & n3398;
  assign n3526 = pi0109 & pi0145;
  assign n3527 = pi0180 & pi0181;
  assign n3528 = n3526 & n3527;
  assign n3529 = pi0182 & pi0232;
  assign n3530 = n3528 & n3529;
  assign n3531 = pi0109 & pi0299;
  assign n3532 = ~n3530 & ~n3531;
  assign n3533 = n3525 & ~n3532;
  assign n3534 = n3519 & ~n3533;
  assign n3535 = n3534 & ~pi0228;
  assign n3536 = n2779 & n2758;
  assign n3537 = ~pi0075 & pi0100;
  assign n3538 = n3455 & n3537;
  assign n3539 = n3536 & n3538;
  assign n3540 = n2788 & ~n3539;
  assign n3541 = n3412 & pi1093;
  assign n3542 = pi0829 & pi1092;
  assign po1107 = n3542 & ~n2643;
  assign n3544 = n3541 & ~po1107;
  assign n3545 = n3544 & n3419;
  assign n3546 = ~n2927 & ~n3464;
  assign n3547 = n3545 & ~n3546;
  assign n3548 = ~n3461 & ~n3465;
  assign n3549 = n3468 & ~n3548;
  assign n3550 = ~n3547 & ~n3549;
  assign n3551 = n2863 & pi0039;
  assign n3552 = ~n3550 & n3551;
  assign n3553 = n2750 & n3552;
  assign n3554 = ~n3553 & ~pi0228;
  assign n3555 = n3540 & n3554;
  assign n3556 = ~pi0030 & pi0228;
  assign n3557 = ~po1038 & ~n3556;
  assign n3558 = ~n3555 & n3557;
  assign n3559 = ~n3535 & ~n3558;
  assign n3560 = n3398 & ~pi0299;
  assign n3561 = ~n3559 & n3560;
  assign n3562 = n3561 & pi0602;
  assign n3563 = n3519 & ~pi0228;
  assign n3564 = n2788 & ~pi0228;
  assign n3565 = po1038 & ~n3556;
  assign n3566 = ~n3564 & n3565;
  assign n3567 = ~n3558 & ~n3566;
  assign n3568 = ~n3563 & n3567;
  assign n3569 = ~n3565 & ~pi0299;
  assign n3570 = pi0109 & ~pi0228;
  assign n3571 = n3523 & n3570;
  assign n3572 = ~n3571 & n3398;
  assign n3573 = ~n3569 & n3572;
  assign n3574 = n3573 & pi0907;
  assign n3575 = n3396 & ~n3398;
  assign n3576 = ~n3574 & ~n3575;
  assign n3577 = ~n3568 & ~n3576;
  assign po0171 = ~n3562 & ~n3577;
  assign n3579 = ~n3559 & ~n3560;
  assign n3580 = ~n3579 & ~n3566;
  assign n3581 = n3393 & ~n3398;
  assign n3582 = n3398 & pi0947;
  assign n3583 = ~n3581 & ~n3582;
  assign n3584 = ~n3580 & ~n3583;
  assign n3585 = n3561 & pi0587;
  assign po0172 = ~n3584 & ~n3585;
  assign n3587 = n3561 & pi0967;
  assign n3588 = ~n3568 & n3573;
  assign n3589 = n3588 & pi0970;
  assign po0173 = ~n3587 & ~n3589;
  assign n3591 = pi0299 & pi0972;
  assign n3592 = n3591 & ~pi0109;
  assign n3593 = ~pi0299 & pi0961;
  assign n3594 = ~n3592 & ~n3593;
  assign n3595 = ~n3530 & ~n3594;
  assign n3596 = ~n3523 & n3591;
  assign n3597 = ~n3595 & ~n3596;
  assign n3598 = n3563 & ~n3597;
  assign n3599 = ~n3591 & ~n3593;
  assign n3600 = n3558 & ~n3599;
  assign n3601 = n3566 & pi0972;
  assign n3602 = ~n3600 & ~n3601;
  assign n3603 = ~n3598 & n3602;
  assign po0174 = n3603 | ~n3398;
  assign n3605 = n3561 & pi0977;
  assign n3606 = n3588 & pi0960;
  assign po0175 = ~n3605 & ~n3606;
  assign n3608 = n3561 & pi0969;
  assign n3609 = n3588 & pi0963;
  assign po0176 = ~n3608 & ~n3609;
  assign n3611 = n3561 & pi0971;
  assign n3612 = n3588 & pi0975;
  assign po0177 = ~n3611 & ~n3612;
  assign n3614 = n3561 & pi0974;
  assign n3615 = n3588 & pi0978;
  assign po0178 = ~n3614 & ~n3615;
  assign n3617 = n2609 & ~pi0096;
  assign n3618 = ~pi0090 & ~pi0093;
  assign n3619 = ~pi0035 & ~pi0070;
  assign n3620 = n3618 & n3619;
  assign n3621 = n3617 & n3620;
  assign n3622 = n2599 & n3621;
  assign n3623 = n2506 & n3622;
  assign n3624 = n2740 & ~pi0092;
  assign n3625 = n3624 & ~po1038;
  assign n3626 = n3623 & n3625;
  assign n3627 = pi0039 & ~pi0072;
  assign n3628 = n3626 & n3627;
  assign n3629 = ~pi0051 & ~pi0087;
  assign n3630 = n2514 & n3629;
  assign n3631 = n3628 & n3630;
  assign n3632 = ~n2885 & n2900;
  assign n3633 = n3463 & n3632;
  assign n3634 = ~po1038 & n2927;
  assign n3635 = n3408 & n3634;
  assign n3636 = ~n3633 & ~n3635;
  assign n3637 = ~n3636 & n3545;
  assign n3638 = ~n3469 & ~n3637;
  assign n3639 = n3631 & ~n3638;
  assign n3640 = n3540 & ~n3639;
  assign po0195 = n3534 | ~n3640;
  assign n3642 = po0195 & ~pi0954;
  assign n3643 = ~pi0024 & pi0954;
  assign po0182 = n3642 | n3643;
  assign n3645 = n2827 & n2665;
  assign n3646 = n2802 & ~n3645;
  assign po0275 = ~n2892 | n3646;
  assign n3648 = po0275 & ~pi0228;
  assign po0183 = n3648 | n2706;
  assign n3650 = ~pi0119 & ~pi0228;
  assign n3651 = pi0252 & ~pi0468;
  assign n3652 = n3650 & n3651;
  assign n3653 = pi0119 & ~pi0468;
  assign n3654 = n3653 & ~pi1056;
  assign po0184 = ~n3652 & ~n3654;
  assign n3656 = n3653 & ~pi1077;
  assign po0185 = ~n3652 & ~n3656;
  assign n3658 = n3653 & ~pi1073;
  assign po0186 = ~n3652 & ~n3658;
  assign n3660 = n3653 & ~pi1041;
  assign po0187 = ~n3652 & ~n3660;
  assign n3662 = n2589 & n2606;
  assign n3663 = n3662 & pi0098;
  assign n3664 = n3618 & pi0051;
  assign n3665 = ~pi0051 & ~pi0841;
  assign n3666 = ~pi0090 ^ ~pi0093;
  assign n3667 = n3665 & n3666;
  assign n3668 = ~n3664 & ~n3667;
  assign n3669 = ~n3668 & n3619;
  assign n3670 = n2600 & n3669;
  assign n3671 = ~n3663 & ~n3670;
  assign n3672 = n3671 & ~pi0096;
  assign n3673 = ~pi0098 & pi1091;
  assign n3674 = ~po0740 & ~n3673;
  assign n3675 = ~n3674 & ~pi0072;
  assign n3676 = n3675 & ~po0950;
  assign n3677 = ~n3672 & n3676;
  assign n3678 = n2675 & pi0091;
  assign n3679 = ~pi0024 & ~pi0058;
  assign n3680 = n3678 & n3679;
  assign n3681 = ~n2634 & ~n3680;
  assign n3682 = n2650 & ~pi0122;
  assign n3683 = n2606 & ~pi0072;
  assign n3684 = n2612 & n3683;
  assign n3685 = n3682 & n3684;
  assign n3686 = ~n3681 & n3685;
  assign n3687 = ~n3677 & ~n3686;
  assign n3688 = n2613 & n2606;
  assign n3689 = ~pi0122 & pi0829;
  assign n3690 = n3689 & ~pi0841;
  assign n3691 = n2609 & n3690;
  assign n3692 = n3688 & n3691;
  assign n3693 = ~n3692 & ~n3617;
  assign n3694 = ~n3687 & ~n3693;
  assign n3695 = ~pi0039 & ~pi0072;
  assign n3696 = n3617 & n3695;
  assign n3697 = ~n3671 & n3696;
  assign n3698 = ~n3697 & ~pi0087;
  assign n3699 = ~n3698 & ~po0950;
  assign n3700 = ~n2794 & ~pi0075;
  assign n3701 = ~n3699 & n3700;
  assign n3702 = ~n3694 & n3701;
  assign n3703 = ~n2662 & pi0299;
  assign n3704 = n3398 & pi0232;
  assign n3705 = ~n3703 & n3704;
  assign n3706 = ~n2658 & ~pi0299;
  assign n3707 = n3705 & ~n3706;
  assign n3708 = po1057 & ~n3707;
  assign n3709 = n3708 & pi0252;
  assign n3710 = ~pi0024 & ~pi0100;
  assign n3711 = n3710 & ~pi0087;
  assign n3712 = n3682 & n3711;
  assign n3713 = n3709 & n3712;
  assign n3714 = n2750 & n3713;
  assign n3715 = ~n3714 & pi0075;
  assign n3716 = n2862 & n2796;
  assign n3717 = n2750 & n3716;
  assign n3718 = ~n3715 & n3717;
  assign n3719 = ~n2927 & ~n2930;
  assign n3720 = n3408 & ~n3719;
  assign n3721 = ~n2708 & n2709;
  assign n3722 = n3463 & n3721;
  assign n3723 = ~n3720 & ~n3722;
  assign n3724 = n2927 & ~pi0224;
  assign n3725 = n3464 & ~pi0216;
  assign n3726 = ~n3724 & ~n3725;
  assign n3727 = ~n3723 & ~n3726;
  assign n3728 = n3727 & n3468;
  assign n3729 = ~n3728 & pi0039;
  assign n3730 = n3682 & n3708;
  assign n3731 = n3730 & pi0228;
  assign n3732 = ~n3731 & pi0100;
  assign n3733 = n2800 & n2741;
  assign n3734 = ~n3732 & n3733;
  assign n3735 = ~n3729 & n3734;
  assign n3736 = n2750 & n3735;
  assign n3737 = ~n3736 & ~n2743;
  assign n3738 = ~n3718 & n3737;
  assign n3739 = ~pi0373 ^ ~pi0374;
  assign n3740 = ~pi0375 ^ ~pi0384;
  assign n3741 = n3739 ^ ~n3740;
  assign n3742 = pi0440 ^ ~pi0442;
  assign n3743 = n3741 ^ ~n3742;
  assign n3744 = pi0370 ^ ~pi0371;
  assign n3745 = n3744 ^ ~pi0369;
  assign n3746 = n3743 ^ ~n3745;
  assign n3747 = n3746 & pi1198;
  assign n3748 = ~pi0380 ^ ~pi0386;
  assign n3749 = ~pi0363 ^ ~pi0372;
  assign n3750 = n3748 ^ ~n3749;
  assign n3751 = pi0387 ^ ~pi0388;
  assign n3752 = n3750 ^ ~n3751;
  assign n3753 = pi0338 ^ ~pi0339;
  assign n3754 = n3753 ^ ~pi0337;
  assign n3755 = n3752 ^ ~n3754;
  assign n3756 = n3755 & pi1196;
  assign n3757 = ~n3747 & ~n3756;
  assign n3758 = ~pi0366 ^ ~pi0367;
  assign n3759 = ~pi0368 ^ ~pi0383;
  assign n3760 = n3758 ^ ~n3759;
  assign n3761 = pi0389 ^ ~pi0447;
  assign n3762 = n3760 ^ ~n3761;
  assign n3763 = pi0364 ^ ~pi0365;
  assign n3764 = n3763 ^ ~pi0336;
  assign n3765 = n3762 ^ ~n3764;
  assign n3766 = n3765 & pi1197;
  assign n3767 = n3757 & ~n3766;
  assign n3768 = pi0378 ^ ~pi0379;
  assign n3769 = pi0385 ^ ~pi0439;
  assign n3770 = ~n3768 ^ ~n3769;
  assign n3771 = ~pi0381 ^ ~pi0382;
  assign n3772 = ~n3770 ^ ~n3771;
  assign n3773 = pi0376 ^ ~pi0377;
  assign n3774 = n3773 ^ ~pi0317;
  assign n3775 = ~n3772 ^ ~n3774;
  assign n3776 = n3775 & pi1199;
  assign n3777 = ~n3776 & ~pi0591;
  assign n3778 = n3767 & n3777;
  assign n3779 = ~n3778 & ~pi0590;
  assign n3780 = ~pi0354 ^ ~pi0356;
  assign n3781 = ~pi0357 ^ ~pi0360;
  assign n3782 = n3780 ^ ~n3781;
  assign n3783 = pi0461 ^ ~pi0462;
  assign n3784 = n3782 ^ ~n3783;
  assign n3785 = pi0352 ^ ~pi0353;
  assign n3786 = n3785 ^ ~pi0351;
  assign n3787 = n3784 ^ ~n3786;
  assign n3788 = n3787 & pi1199;
  assign n3789 = pi0361 ^ ~pi0441;
  assign n3790 = pi0458 ^ ~pi0460;
  assign n3791 = ~n3789 ^ ~n3790;
  assign n3792 = ~pi0452 ^ ~pi0455;
  assign n3793 = ~n3791 ^ ~n3792;
  assign n3794 = pi0342 ^ ~pi0355;
  assign n3795 = n3794 ^ ~pi0320;
  assign n3796 = ~n3793 ^ ~n3795;
  assign n3797 = n3796 & pi1196;
  assign n3798 = ~n3788 & ~n3797;
  assign n3799 = pi0322 ^ ~pi0347;
  assign n3800 = pi0350 ^ ~pi0359;
  assign n3801 = ~n3799 ^ ~n3800;
  assign n3802 = ~pi0348 ^ ~pi0349;
  assign n3803 = ~n3801 ^ ~n3802;
  assign n3804 = pi0316 ^ ~pi0321;
  assign n3805 = n3804 ^ ~pi0315;
  assign n3806 = ~n3803 ^ ~n3805;
  assign n3807 = n3806 & pi1198;
  assign n3808 = ~pi0344 ^ ~pi0345;
  assign n3809 = ~pi0346 ^ ~pi0358;
  assign n3810 = n3808 ^ ~n3809;
  assign n3811 = pi0362 ^ ~pi0450;
  assign n3812 = n3810 ^ ~n3811;
  assign n3813 = pi0327 ^ ~pi0343;
  assign n3814 = n3813 ^ ~pi0323;
  assign n3815 = n3812 ^ ~n3814;
  assign n3816 = n3815 & pi1197;
  assign n3817 = ~n3807 & ~n3816;
  assign n3818 = n3798 & n3817;
  assign n3819 = ~pi0591 & ~pi0592;
  assign n3820 = ~n3818 & n3819;
  assign n3821 = ~n3779 & ~n3820;
  assign n3822 = ~pi0590 & ~pi0592;
  assign n3823 = n3822 & ~pi0591;
  assign n3824 = ~n3821 & ~n3823;
  assign n3825 = n3824 & pi0588;
  assign n3826 = ~n3825 & ~pi0217;
  assign n3827 = ~pi0423 ^ ~pi0424;
  assign n3828 = ~pi0425 ^ ~pi0432;
  assign n3829 = n3827 ^ ~n3828;
  assign n3830 = pi0454 ^ ~pi0459;
  assign n3831 = n3829 ^ ~n3830;
  assign n3832 = pi0420 ^ ~pi0421;
  assign n3833 = n3832 ^ ~pi0419;
  assign n3834 = n3831 ^ ~n3833;
  assign n3835 = n3834 & pi1198;
  assign n3836 = ~pi0437 ^ ~pi0438;
  assign n3837 = ~pi0418 ^ ~pi0431;
  assign n3838 = n3836 ^ ~n3837;
  assign n3839 = pi0453 ^ ~pi0464;
  assign n3840 = n3838 ^ ~n3839;
  assign n3841 = pi0416 ^ ~pi0417;
  assign n3842 = n3841 ^ ~pi0415;
  assign n3843 = n3840 ^ ~n3842;
  assign n3844 = n3843 & pi1197;
  assign n3845 = ~n3835 & ~n3844;
  assign n3846 = ~pi0445 ^ ~pi0448;
  assign n3847 = ~pi0430 ^ ~pi0433;
  assign n3848 = n3846 ^ ~n3847;
  assign n3849 = pi0449 ^ ~pi0451;
  assign n3850 = n3848 ^ ~n3849;
  assign n3851 = pi0427 ^ ~pi0428;
  assign n3852 = n3851 ^ ~pi0426;
  assign n3853 = n3850 ^ ~n3852;
  assign n3854 = n3853 & pi1199;
  assign n3855 = pi0434 ^ ~pi0435;
  assign n3856 = pi0444 ^ ~pi0446;
  assign n3857 = ~n3855 ^ ~n3856;
  assign n3858 = ~pi0436 ^ ~pi0443;
  assign n3859 = ~n3857 ^ ~n3858;
  assign n3860 = pi0422 ^ ~pi0429;
  assign n3861 = n3860 ^ ~pi0414;
  assign n3862 = ~n3859 ^ ~n3861;
  assign n3863 = n3862 & pi1196;
  assign n3864 = ~n3854 & ~n3863;
  assign n3865 = n3845 & n3864;
  assign n3866 = n3822 & pi0588;
  assign n3867 = ~n3865 & n3866;
  assign n3868 = ~n3824 & ~n3867;
  assign n3869 = n3826 & ~n3868;
  assign n3870 = ~pi0391 ^ ~pi0392;
  assign n3871 = ~pi0393 ^ ~pi0407;
  assign n3872 = n3870 ^ ~n3871;
  assign n3873 = pi0413 ^ ~pi0463;
  assign n3874 = n3872 ^ ~n3873;
  assign n3875 = pi0334 ^ ~pi0335;
  assign n3876 = n3875 ^ ~pi0333;
  assign n3877 = n3874 ^ ~n3876;
  assign n3878 = n3877 & pi1197;
  assign n3879 = pi0395 ^ ~pi0396;
  assign n3880 = pi0400 ^ ~pi0408;
  assign n3881 = ~n3879 ^ ~n3880;
  assign n3882 = ~pi0398 ^ ~pi0399;
  assign n3883 = ~n3881 ^ ~n3882;
  assign n3884 = pi0329 ^ ~pi0394;
  assign n3885 = n3884 ^ ~pi0328;
  assign n3886 = ~n3883 ^ ~n3885;
  assign n3887 = n3886 & pi1198;
  assign n3888 = ~n3878 & ~n3887;
  assign n3889 = ~n3888 & ~pi0592;
  assign n3890 = ~n3889 & pi0591;
  assign n3891 = ~pi0410 ^ ~pi0411;
  assign n3892 = ~pi0397 ^ ~pi0404;
  assign n3893 = n3891 ^ ~n3892;
  assign n3894 = pi0412 ^ ~pi0456;
  assign n3895 = n3893 ^ ~n3894;
  assign n3896 = pi0324 ^ ~pi0390;
  assign n3897 = n3896 ^ ~pi0319;
  assign n3898 = n3895 ^ ~n3897;
  assign n3899 = n3898 & pi1196;
  assign n3900 = pi0401 ^ ~pi0402;
  assign n3901 = pi0406 ^ ~pi0409;
  assign n3902 = ~n3900 ^ ~n3901;
  assign n3903 = ~pi0403 ^ ~pi0405;
  assign n3904 = ~n3902 ^ ~n3903;
  assign n3905 = pi0325 ^ ~pi0326;
  assign n3906 = n3905 ^ ~pi0318;
  assign n3907 = ~n3904 ^ ~n3906;
  assign n3908 = n3907 & pi1199;
  assign n3909 = ~n3899 & ~n3908;
  assign n3910 = ~n3909 & n3822;
  assign n3911 = n3910 & pi0567;
  assign n3912 = n3890 & ~n3911;
  assign n3913 = n3869 & ~n3912;
  assign n3914 = n3913 & n2643;
  assign n3915 = ~n3738 & ~n3914;
  assign n3916 = ~n3702 & n3915;
  assign n3917 = n3869 & ~n3890;
  assign n3918 = ~pi0286 & ~pi0289;
  assign n3919 = ~pi0285 & ~pi0288;
  assign n3920 = n3918 & n3919;
  assign n3921 = ~n3917 & ~n3920;
  assign n3922 = ~n3916 & ~n3921;
  assign n3923 = pi1092 & pi1093;
  assign n3924 = ~pi0098 & pi0567;
  assign n3925 = n3923 & ~n3924;
  assign n3926 = ~pi1161 & ~pi1162;
  assign n3927 = n3926 & ~pi1163;
  assign n3928 = ~n3925 & n3927;
  assign n3929 = ~po1038 & n3928;
  assign n3930 = ~n3922 & n3929;
  assign n3931 = ~n3670 & ~n2794;
  assign n3932 = n3411 & n2643;
  assign n3933 = n3696 & n3932;
  assign n3934 = n3670 & ~n3933;
  assign n3935 = ~n3931 & ~n3934;
  assign n3936 = ~po0740 & pi0567;
  assign n3937 = ~n3936 & ~pi1199;
  assign n3938 = ~pi0217 & ~pi0588;
  assign n3939 = pi0591 & ~pi1091;
  assign n3940 = n3938 & n3939;
  assign n3941 = ~n3937 & n3940;
  assign n3942 = n3941 & n3888;
  assign n3943 = n3942 & n3910;
  assign n3944 = n3935 & ~n3943;
  assign n3945 = ~n3694 & ~n3944;
  assign n3946 = ~n3945 & ~n3737;
  assign n3947 = ~po0950 & ~n2759;
  assign n3948 = n3718 & n3947;
  assign n3949 = n3932 & ~pi0122;
  assign n3950 = n3949 & ~pi0098;
  assign n3951 = ~n3948 & ~n3950;
  assign n3952 = n3943 & n3936;
  assign n3953 = ~n3951 & ~n3952;
  assign n3954 = ~n3946 & ~n3953;
  assign n3955 = n3930 & ~n3954;
  assign n3956 = n3949 & ~n3920;
  assign n3957 = n3924 & n3926;
  assign n3958 = n3956 & n3957;
  assign n3959 = n3958 & po1038;
  assign n3960 = ~n3913 & n3959;
  assign n3961 = n3923 & ~pi0031;
  assign n3962 = pi1161 & pi1162;
  assign n3963 = n3961 & n3962;
  assign n3964 = ~n3960 & ~n3963;
  assign n3965 = ~n3964 & ~pi1163;
  assign po0189 = n3955 | n3965;
  assign n3967 = n2511 & pi0076;
  assign n3968 = ~po0840 & ~n3920;
  assign n3969 = ~n2668 & ~pi0137;
  assign n3970 = n3969 & ~pi0050;
  assign n3971 = ~n3968 & n3970;
  assign n3972 = n3967 & n3971;
  assign n3973 = n2545 & ~pi0024;
  assign n3974 = n3973 & pi0050;
  assign n3975 = n2668 & ~pi0841;
  assign n3976 = ~pi0024 & ~pi0841;
  assign n3977 = ~n3976 & pi0032;
  assign n3978 = ~n3975 & n3977;
  assign n3979 = ~n3974 & ~n3978;
  assign n3980 = ~n3972 & n3979;
  assign n3981 = n2891 & ~n3980;
  assign n3982 = ~n3448 & ~pi0129;
  assign n3983 = ~n3452 & ~n3982;
  assign n3984 = n3983 & n3537;
  assign n3985 = n3984 & ~n3453;
  assign n3986 = ~n3708 & pi0252;
  assign n3987 = n3710 & pi0075;
  assign n3988 = ~po0840 & n3987;
  assign n3989 = ~n3986 & n3988;
  assign n3990 = ~n3985 & ~n3989;
  assign n3991 = n3988 & n2665;
  assign n3992 = n3708 & ~n3991;
  assign n3993 = ~n3992 & ~pi0137;
  assign n3994 = ~n3990 & n3993;
  assign n3995 = n3536 & n3994;
  assign po0190 = n3981 | n3995;
  assign n3997 = n2538 & ~pi0070;
  assign n3998 = ~n2621 & ~n3997;
  assign n3999 = ~n3513 & n2588;
  assign n4000 = ~n3998 & ~n3999;
  assign n4001 = n3502 & pi0073;
  assign n4002 = n2622 & n2608;
  assign n4003 = n4001 & n4002;
  assign n4004 = n4000 & ~n4003;
  assign n4005 = ~pi0195 & ~pi0196;
  assign n4006 = ~pi0138 & ~pi0139;
  assign n4007 = n4005 & n4006;
  assign n4008 = ~pi0079 & ~pi0118;
  assign n4009 = ~pi0033 & ~pi0034;
  assign n4010 = n4008 & n4009;
  assign po0997 = n4007 & n4010;
  assign n4012 = ~pi0033 ^ ~pi0954;
  assign n4013 = ~po0997 & ~n4012;
  assign n4014 = ~pi0063 & ~pi0107;
  assign n4015 = n4014 & ~pi0040;
  assign n4016 = ~n4013 & n4015;
  assign n4017 = pi0164 & pi0299;
  assign n4018 = pi0186 & ~pi0299;
  assign n4019 = ~n4017 & ~n4018;
  assign n4020 = n3704 & ~n4019;
  assign n4021 = ~n4020 & ~n2739;
  assign n4022 = n2768 & ~n4021;
  assign n4023 = n4016 & n4022;
  assign n4024 = n4004 & n4023;
  assign n4025 = ~n3406 & n3461;
  assign n4026 = n4025 & ~pi0174;
  assign n4027 = ~n3429 & n3465;
  assign n4028 = n4027 & ~pi0152;
  assign n4029 = ~n4026 & ~n4028;
  assign n4030 = n3545 & ~n4029;
  assign n4031 = n4025 & pi0176;
  assign n4032 = n4027 & pi0154;
  assign n4033 = ~n4031 & ~n4032;
  assign n4034 = n3468 & ~n4033;
  assign n4035 = ~n4030 & ~n4034;
  assign n4036 = n2750 & ~n4035;
  assign n4037 = ~n4036 & pi0039;
  assign n4038 = ~n4037 & n3704;
  assign n4039 = n3504 & n2608;
  assign n4040 = ~n3468 & ~n3545;
  assign n4041 = ~n3467 & ~n4040;
  assign n4042 = n4039 & n4041;
  assign n4043 = n4042 & n2741;
  assign n4044 = ~n4038 & n4043;
  assign n4045 = n4039 & n2764;
  assign n4046 = n4045 & pi0092;
  assign n4047 = pi0176 & ~pi0299;
  assign n4048 = pi0154 & pi0299;
  assign n4049 = ~n4047 & ~n4048;
  assign n4050 = n3704 & ~n4049;
  assign n4051 = n4050 & n4015;
  assign n4052 = n4046 & n4051;
  assign n4053 = n4016 & ~n2742;
  assign n4054 = ~n4045 & n4053;
  assign n4055 = ~n4052 & ~n4054;
  assign n4056 = ~n4044 & ~n4055;
  assign n4057 = n3696 & n2741;
  assign n4058 = n3688 & n4057;
  assign n4059 = ~n4058 & pi0038;
  assign n4060 = ~n4059 & ~pi0054;
  assign n4061 = ~n4056 & n4060;
  assign n4062 = ~n4021 & ~pi0074;
  assign n4063 = ~n4061 & n4062;
  assign n4064 = pi0191 & ~pi0299;
  assign n4065 = pi0169 & pi0299;
  assign n4066 = ~n4064 & ~n4065;
  assign n4067 = n3704 & ~n4066;
  assign n4068 = n4067 & pi0074;
  assign n4069 = ~n4068 & n2737;
  assign n4070 = ~n4063 & n4069;
  assign n4071 = n3704 & ~n2737;
  assign n4072 = ~pi0149 ^ ~pi0157;
  assign n4073 = ~n4072 & pi0299;
  assign n4074 = ~pi0178 ^ ~pi0183;
  assign n4075 = ~n4074 & ~pi0299;
  assign n4076 = ~n4073 & ~n4075;
  assign n4077 = n4071 & n4076;
  assign n4078 = ~n4070 & ~n4077;
  assign n4079 = ~n4078 & ~po1038;
  assign n4080 = ~n4024 & n4079;
  assign n4081 = n2588 & n3511;
  assign n4082 = ~pi0172 & pi0299;
  assign n4083 = ~pi0193 & ~pi0299;
  assign n4084 = ~n4082 & ~n4083;
  assign n4085 = n4081 & n4084;
  assign n4086 = pi0158 & pi0299;
  assign n4087 = pi0180 & ~pi0299;
  assign n4088 = ~n4086 & ~n4087;
  assign n4089 = ~n4088 & n2694;
  assign n4090 = n2623 & n4089;
  assign n4091 = n2627 & ~pi0841;
  assign n4092 = n4091 & n2666;
  assign n4093 = n3504 & n4092;
  assign n4094 = ~n3997 & ~pi0299;
  assign n4095 = ~n4093 & ~n4094;
  assign n4096 = ~n4095 & pi0183;
  assign n4097 = pi0032 & ~pi0841;
  assign n4098 = n4097 & ~pi0210;
  assign n4099 = n3997 & ~n4098;
  assign n4100 = ~n4099 & pi0149;
  assign n4101 = ~n4100 & ~pi0073;
  assign n4102 = pi0073 & pi0152;
  assign n4103 = ~n4102 & pi0299;
  assign n4104 = pi0073 & ~pi0299;
  assign n4105 = n4104 & ~pi0174;
  assign n4106 = ~n4103 & ~n4105;
  assign n4107 = ~n4101 & ~n4106;
  assign n4108 = ~n4096 & ~n4107;
  assign n4109 = ~n4090 & n4108;
  assign n4110 = ~n4085 & n4109;
  assign n4111 = n2631 & ~n4110;
  assign n4112 = ~n4111 & ~pi0039;
  assign n4113 = n4038 & n2863;
  assign n4114 = ~n4112 & n4113;
  assign n4115 = n4080 & ~n4114;
  assign n4116 = n2751 & n2744;
  assign n4117 = ~n4116 & ~n4013;
  assign n4118 = n3704 & pi0149;
  assign n4119 = n4116 & n4118;
  assign n4120 = ~n4117 & ~n4119;
  assign n4121 = n2746 & n2739;
  assign n4122 = n2738 & n4121;
  assign n4123 = n4122 & n4015;
  assign n4124 = ~n4120 & n4123;
  assign n4125 = ~n4121 & ~pi0074;
  assign n4126 = n4125 & pi0164;
  assign n4127 = pi0074 & pi0169;
  assign n4128 = ~n4126 & ~n4127;
  assign n4129 = ~n4128 & n3704;
  assign n4130 = ~n4129 & n2737;
  assign n4131 = n4071 & n4072;
  assign n4132 = ~n4130 & ~n4131;
  assign n4133 = ~n4132 & po1038;
  assign n4134 = ~n4124 & n4133;
  assign po0191 = n4115 | n4134;
  assign n4136 = n4004 & n2748;
  assign n4137 = n2742 & n2744;
  assign n4138 = n4039 & n4137;
  assign n4139 = ~n4138 & ~n2745;
  assign n4140 = ~n4136 & ~n4139;
  assign n4141 = ~pi0033 & ~pi0954;
  assign n4142 = n4141 & ~pi0034;
  assign n4143 = ~po0997 & n4142;
  assign n4144 = ~n4141 & pi0034;
  assign n4145 = ~n4143 & ~n4144;
  assign n4146 = ~n4140 & n4145;
  assign n4147 = ~n4046 & n4145;
  assign n4148 = n4043 & pi0039;
  assign n4149 = ~n4147 & ~n4148;
  assign n4150 = pi0155 & pi0299;
  assign n4151 = pi0177 & ~pi0299;
  assign n4152 = ~n4150 & ~n4151;
  assign n4153 = n3704 & ~n4152;
  assign n4154 = n4046 & n4153;
  assign n4155 = n4149 & ~n4154;
  assign n4156 = n4025 & ~pi0144;
  assign n4157 = n4027 & ~pi0161;
  assign n4158 = ~n4156 & ~n4157;
  assign n4159 = ~n4158 & n3544;
  assign n4160 = n4025 & pi0177;
  assign n4161 = n4027 & pi0155;
  assign n4162 = ~n4160 & ~n4161;
  assign n4163 = ~n4162 & n2650;
  assign n4164 = ~n4159 & ~n4163;
  assign n4165 = ~n4164 & n3704;
  assign n4166 = n4043 & ~n4165;
  assign n4167 = ~n2743 & n2745;
  assign n4168 = ~n4166 & n4167;
  assign n4169 = ~n4155 & n4168;
  assign n4170 = ~n4146 & ~n4169;
  assign n4171 = ~n4170 & n4123;
  assign n4172 = ~n2659 & ~n2663;
  assign n4173 = n4081 & ~n4172;
  assign n4174 = ~n4095 & pi0140;
  assign n4175 = pi0162 & pi0299;
  assign n4176 = ~n4099 & n4175;
  assign n4177 = pi0161 & pi0299;
  assign n4178 = ~n4177 & pi0073;
  assign n4179 = pi0144 & ~pi0299;
  assign n4180 = n4178 & ~n4179;
  assign n4181 = pi0159 & pi0299;
  assign n4182 = pi0181 & ~pi0299;
  assign n4183 = ~n4181 & ~n4182;
  assign n4184 = n3505 & ~n4183;
  assign n4185 = ~n4180 & ~n4184;
  assign n4186 = ~n4176 & n4185;
  assign n4187 = ~n4174 & n4186;
  assign n4188 = ~n4173 & n4187;
  assign n4189 = n2891 & ~n4188;
  assign n4190 = ~pi0188 & ~pi0299;
  assign n4191 = ~pi0167 & pi0299;
  assign n4192 = ~n4190 & ~n4191;
  assign n4193 = n4192 & ~pi0074;
  assign n4194 = ~n4060 & n4193;
  assign n4195 = pi0148 & pi0299;
  assign n4196 = pi0141 & ~pi0299;
  assign n4197 = ~n4195 & ~n4196;
  assign n4198 = ~n4197 & pi0074;
  assign n4199 = ~po1038 & ~n4198;
  assign n4200 = ~n4194 & n4199;
  assign n4201 = n4125 & pi0167;
  assign n4202 = pi0074 & pi0148;
  assign n4203 = po1038 & ~n4202;
  assign n4204 = ~n4201 & n4203;
  assign n4205 = ~n4204 & n2737;
  assign n4206 = ~n4200 & n4205;
  assign n4207 = ~pi0149 & ~pi0157;
  assign n4208 = ~pi0162 ^ ~pi0197;
  assign n4209 = ~n4207 ^ ~n4208;
  assign n4210 = ~n2885 & n4209;
  assign n4211 = ~n4210 & ~n2737;
  assign n4212 = ~pi0178 & ~pi0183;
  assign n4213 = ~pi0140 ^ ~pi0145;
  assign n4214 = n4212 ^ ~n4213;
  assign n4215 = n2885 & ~n4214;
  assign n4216 = n4211 & ~n4215;
  assign n4217 = ~n4206 & ~n4216;
  assign n4218 = ~n4189 & n4217;
  assign n4219 = n2805 & n4138;
  assign n4220 = n4219 & pi0162;
  assign n4221 = n4218 & ~n4220;
  assign n4222 = ~n4221 & n3704;
  assign po0192 = ~n4171 & ~n4222;
  assign n4224 = pi0035 & ~pi0093;
  assign n4225 = n4224 & pi0841;
  assign n4226 = ~pi0035 & pi0093;
  assign n4227 = n4226 & ~pi0841;
  assign n4228 = ~n4225 & ~n4227;
  assign n4229 = n3491 & n4228;
  assign n4230 = ~po0740 & ~pi0122;
  assign n4231 = ~n3968 & n4230;
  assign n4232 = ~n3969 & pi0076;
  assign n4233 = n4231 & n4232;
  assign n4234 = ~n2675 & ~n4233;
  assign n4235 = ~n4229 & ~n4234;
  assign n4236 = pi0040 & pi1082;
  assign n4237 = ~n4235 & ~n4236;
  assign n4238 = n2631 & ~n4237;
  assign n4239 = ~n3499 & n2772;
  assign n4240 = pi0024 & ~pi0059;
  assign n4241 = ~n4239 & ~n4240;
  assign n4242 = ~n4238 & ~n4241;
  assign n4243 = ~n4058 & n4125;
  assign n4244 = ~n4243 & n2767;
  assign n4245 = ~n4242 & n4244;
  assign n4246 = ~po0840 & pi0137;
  assign n4247 = ~n3986 & ~n4246;
  assign n4248 = po1057 & ~n2665;
  assign n4249 = ~pi0038 & pi0075;
  assign n4250 = ~n4248 & n4249;
  assign n4251 = ~n4247 & n4250;
  assign n4252 = pi0038 & ~pi0075;
  assign n4253 = ~n4251 & ~n4252;
  assign n4254 = ~n4253 & n3710;
  assign n4255 = n3708 & n3412;
  assign n4256 = n4255 & pi0683;
  assign n4257 = ~n3708 & pi0137;
  assign n4258 = ~n4257 & pi0252;
  assign n4259 = ~n4256 & n4258;
  assign n4260 = ~n2665 & ~pi0137;
  assign n4261 = ~n4260 & n2739;
  assign n4262 = ~n4248 & n4261;
  assign n4263 = n3984 & n4262;
  assign n4264 = ~n4259 & n4263;
  assign n4265 = ~n4254 & ~n4264;
  assign n4266 = n4058 & ~n4265;
  assign n4267 = n4242 & n4266;
  assign n4268 = ~n4245 & ~n4267;
  assign n4269 = pi0024 & pi0059;
  assign n4270 = ~pi0055 & ~pi0074;
  assign n4271 = ~n4269 & n4270;
  assign n4272 = n2771 & n4271;
  assign po0193 = ~n4268 & n4272;
  assign n4274 = n2599 & pi0036;
  assign n4275 = n2511 & n4274;
  assign n4276 = ~n3680 & ~n4275;
  assign n4277 = n3477 & n2612;
  assign n4278 = ~n4276 & n4277;
  assign po0194 = n4278 & po0740;
  assign n4280 = n4277 & n2599;
  assign n4281 = n2511 & n4280;
  assign n4282 = n4281 & ~pi0841;
  assign n4283 = ~pi0070 & ~pi0089;
  assign n4284 = ~n4283 & pi0332;
  assign n4285 = n4282 & n4284;
  assign n4286 = n2535 & n4280;
  assign n4287 = n4286 & pi0064;
  assign n4288 = n4287 & ~pi0841;
  assign n4289 = ~n4285 & ~n4288;
  assign n4290 = n2763 & pi0024;
  assign po0196 = ~n4289 | n4290;
  assign n4292 = ~po0740 & ~pi0986;
  assign n4293 = ~n4292 & pi0252;
  assign n4294 = pi0108 & pi0314;
  assign n4295 = ~n4293 & n4294;
  assign n4296 = ~pi0035 & ~pi0048;
  assign n4297 = n4296 & ~pi0047;
  assign n4298 = ~n4295 & n4297;
  assign n4299 = ~n4296 & pi0841;
  assign n4300 = ~n4298 & ~n4299;
  assign n4301 = n3498 & n4300;
  assign n4302 = n2700 & n3975;
  assign n4303 = n4302 & n2748;
  assign n4304 = n3631 & ~pi0287;
  assign n4305 = ~n3422 & ~pi1093;
  assign n4306 = ~n3431 & pi0835;
  assign n4307 = n3414 & n4306;
  assign n4308 = ~n4305 & n4307;
  assign n4309 = pi0835 & pi0984;
  assign n4310 = ~n4309 & ~pi0979;
  assign n4311 = n4310 & ~n3417;
  assign n4312 = pi0786 & ~pi1082;
  assign n4313 = n4311 & n4312;
  assign n4314 = ~n4307 & n4313;
  assign n4315 = ~n4314 & n4311;
  assign n4316 = ~n4308 & n4315;
  assign n4317 = n4304 & n4316;
  assign n4318 = ~n4303 & ~n4317;
  assign po0197 = n4301 | ~n4318;
  assign n4320 = pi0040 & ~pi1082;
  assign n4321 = n4320 & ~pi0102;
  assign n4322 = ~pi0040 & pi0102;
  assign n4323 = ~n4321 & ~n4322;
  assign po0198 = n2891 & ~n4323;
  assign n4325 = ~po0840 & ~n2605;
  assign n4326 = ~n3672 & ~n4325;
  assign n4327 = ~n3730 & n3537;
  assign n4328 = ~n4327 & ~n2759;
  assign n4329 = ~n4328 & pi0228;
  assign n4330 = ~n3686 & n4329;
  assign n4331 = ~n4326 & n4330;
  assign n4332 = ~pi0250 & pi0252;
  assign n4333 = pi0901 & ~pi0959;
  assign n4334 = n4332 & n4333;
  assign n4335 = pi0094 & ~pi0110;
  assign n4336 = n4334 & n4335;
  assign n4337 = ~pi0094 & pi0110;
  assign n4338 = ~pi0480 & pi0949;
  assign n4339 = n4337 & n4338;
  assign n4340 = ~n4336 & ~n4339;
  assign n4341 = ~n3662 & ~n4340;
  assign n4342 = ~pi0087 & ~pi0100;
  assign n4343 = ~n2750 & ~n4342;
  assign n4344 = n4340 & ~pi0228;
  assign n4345 = pi0087 & pi0100;
  assign n4346 = n2862 & ~n4345;
  assign n4347 = ~po1038 & n4346;
  assign n4348 = ~n4344 & n4347;
  assign n4349 = ~n4343 & n4348;
  assign n4350 = ~n3715 & n4349;
  assign n4351 = n4350 & ~n3693;
  assign n4352 = ~n4341 & n4351;
  assign n4353 = ~n4331 & n4352;
  assign n4354 = n4353 & ~pi0044;
  assign n4355 = n4354 & ~pi0101;
  assign n4356 = n4355 ^ ~pi0041;
  assign n4357 = n4356 & n3695;
  assign n4358 = n3630 & pi0287;
  assign n4359 = n3626 & n4358;
  assign n4360 = ~n4359 & n3704;
  assign n4361 = ~n2885 & pi0161;
  assign n4362 = n4361 & n2661;
  assign n4363 = n2885 & pi0144;
  assign n4364 = n4363 & n2657;
  assign n4365 = ~n4362 & ~n4364;
  assign n4366 = n4360 & ~n4365;
  assign n4367 = ~n4366 & n3627;
  assign po0199 = ~n4357 & ~n4367;
  assign n4369 = n4354 & n3436;
  assign n4370 = n4369 & n3440;
  assign n4371 = n4370 & ~pi0114;
  assign n4372 = n4371 ^ ~pi0042;
  assign n4373 = ~n4372 & n3695;
  assign n4374 = n2885 & ~pi0189;
  assign n4375 = ~n2885 & ~pi0166;
  assign n4376 = ~n4374 & ~n4375;
  assign n4377 = n4360 & ~n4376;
  assign n4378 = ~n4377 & n3627;
  assign n4379 = ~pi0199 & ~pi0200;
  assign n4380 = ~n4379 & ~pi0299;
  assign n4381 = ~po1038 & n4380;
  assign n4382 = pi0207 & pi0208;
  assign n4383 = ~n4382 & ~pi0199;
  assign n4384 = n4381 & ~n4383;
  assign n4385 = pi0212 & pi0214;
  assign n4386 = n4385 & pi0211;
  assign n4387 = ~n2885 & n4386;
  assign n4388 = ~n4384 & ~n4387;
  assign n4389 = ~n2885 & pi0219;
  assign n4390 = n4388 & ~n4389;
  assign n4391 = n4378 & ~n4390;
  assign po0200 = n4373 | n4391;
  assign n4393 = n4371 & ~pi0042;
  assign n4394 = n4393 ^ ~pi0043;
  assign n4395 = ~n4394 & n3695;
  assign n4396 = ~n4382 & ~pi0200;
  assign n4397 = ~n4379 & n4382;
  assign n4398 = ~n4396 & ~n4397;
  assign n4399 = n2885 & ~n4398;
  assign n4400 = ~pi0211 & ~pi0219;
  assign n4401 = n4385 & n4400;
  assign n4402 = ~n4385 & pi0211;
  assign n4403 = ~n4401 & ~n4402;
  assign n4404 = ~n2885 & n4403;
  assign n4405 = ~n4399 & ~n4404;
  assign n4406 = n4378 & n4405;
  assign po0201 = n4395 | n4406;
  assign n4408 = n4353 ^ ~pi0044;
  assign n4409 = ~n4408 & n3695;
  assign n4410 = n4360 & n3627;
  assign n4411 = n2885 & n2658;
  assign n4412 = ~n2885 & n2662;
  assign n4413 = ~n4411 & ~n4412;
  assign n4414 = n4410 & ~n4413;
  assign po0202 = n4409 | n4414;
  assign po0203 = n4304 & pi0979;
  assign n4417 = pi0046 & ~pi0109;
  assign n4418 = n3477 & n4417;
  assign n4419 = n2563 & n4418;
  assign n4420 = n2588 & n4419;
  assign n4421 = n4420 & pi0024;
  assign n4422 = n4282 & pi0061;
  assign po0204 = n4421 | n4422;
  assign n4424 = ~po0840 & ~n3449;
  assign n4425 = n4278 & n4424;
  assign n4426 = ~n4281 & ~n4286;
  assign n4427 = ~pi0036 & ~pi0088;
  assign n4428 = n4427 & ~pi0104;
  assign n4429 = ~n3412 & ~n4428;
  assign n4430 = ~n4426 & n4429;
  assign n4431 = n4276 & n4430;
  assign po0205 = n4425 | n4431;
  assign n4433 = n4281 & pi0841;
  assign po0206 = n4433 & pi0048;
  assign n4435 = n3710 & pi0074;
  assign n4436 = n2786 & n4435;
  assign n4437 = n4433 & pi0049;
  assign po0207 = n4436 | n4437;
  assign n4439 = n2589 & n4277;
  assign n4440 = pi0024 & pi0050;
  assign n4441 = n4439 & n4440;
  assign n4442 = ~n3538 & ~n3988;
  assign n4443 = ~n4442 & n4248;
  assign n4444 = n3536 & n4443;
  assign n4445 = n4277 & ~pi0058;
  assign n4446 = n2591 & ~pi0086;
  assign n4447 = n2541 & n4446;
  assign n4448 = n4445 & n4447;
  assign n4449 = n2545 & n4448;
  assign n4450 = n4449 & n4335;
  assign n4451 = ~n3708 & ~pi0252;
  assign n4452 = ~po0840 & pi0252;
  assign n4453 = ~n4451 & ~n4452;
  assign n4454 = n4450 & n4453;
  assign n4455 = ~n4444 & ~n4454;
  assign po0208 = n4441 | ~n4455;
  assign n4457 = n2451 & n2452;
  assign n4458 = n4280 & n2509;
  assign n4459 = n4457 & n4458;
  assign n4460 = pi0082 & ~pi0111;
  assign po0209 = n4459 & n4460;
  assign n4462 = n4353 & n3442;
  assign n4463 = ~n4462 ^ ~pi0052;
  assign n4464 = n4463 & n3695;
  assign n4465 = ~pi0211 & pi0219;
  assign n4466 = ~n2885 & ~n4465;
  assign n4467 = ~n4403 & ~pi0219;
  assign n4468 = pi0211 & ~pi0219;
  assign n4469 = ~n4467 & ~n4468;
  assign n4470 = n4466 & n4469;
  assign n4471 = ~pi0199 & pi0200;
  assign n4472 = ~n4471 & ~pi0299;
  assign n4473 = ~po1038 & n4472;
  assign n4474 = ~n4383 & ~pi0200;
  assign n4475 = n4473 & ~n4474;
  assign n4476 = ~n4470 & ~n4475;
  assign n4477 = n4390 & ~n4476;
  assign n4478 = n4378 & n4477;
  assign po0210 = n4464 | n4478;
  assign n4480 = n4309 & ~pi0979;
  assign n4481 = n4304 & n4480;
  assign n4482 = n4445 & n2595;
  assign n4483 = n3372 & n4482;
  assign n4484 = pi0053 & ~pi0060;
  assign n4485 = n4483 & n4484;
  assign n4486 = n4485 & pi0024;
  assign po0211 = n4481 | n4486;
  assign n4488 = n2787 & pi0024;
  assign n4489 = n4488 & n2768;
  assign n4490 = n4282 & pi0106;
  assign po0212 = n4489 | n4490;
  assign n4492 = n4219 & pi0024;
  assign n4493 = n4281 & pi0045;
  assign po0213 = n4492 | n4493;
  assign n4495 = ~pi0062 & pi0841;
  assign n4496 = n4495 & n2791;
  assign n4497 = pi0055 & ~pi0056;
  assign n4498 = ~pi0024 & ~pi0062;
  assign n4499 = n4497 & n4498;
  assign n4500 = ~n4496 & ~n4499;
  assign po0214 = n2789 & ~n4500;
  assign n4502 = n2792 & ~pi0841;
  assign n4503 = pi0062 & pi0924;
  assign n4504 = n4502 & ~n4503;
  assign n4505 = n2755 & pi0024;
  assign po0215 = n4504 | n4505;
  assign n4507 = n3478 & n2600;
  assign po0216 = n4507 & ~pi0841;
  assign n4509 = n4502 & n4503;
  assign n4510 = n2745 & ~pi0057;
  assign n4511 = n4510 & n4269;
  assign n4512 = n2751 & n4511;
  assign po0217 = n4509 | n4512;
  assign n4514 = n4310 & n3417;
  assign n4515 = n4304 & n4514;
  assign n4516 = ~pi0053 & pi0060;
  assign n4517 = n4483 & n4516;
  assign n4518 = n4517 & pi0024;
  assign po0218 = n4515 | n4518;
  assign n4520 = n4433 & pi0061;
  assign n4521 = n4517 & ~pi0024;
  assign po0219 = n4520 | n4521;
  assign n4523 = ~n4498 & pi0057;
  assign n4524 = pi0062 & pi0841;
  assign n4525 = ~n4524 & ~pi0057;
  assign n4526 = ~n4523 & ~n4525;
  assign po0220 = ~n2804 & n4526;
  assign n4528 = n4420 & ~pi0024;
  assign n4529 = n4286 & pi0063;
  assign n4530 = n4529 & pi0999;
  assign po0221 = n4528 | n4530;
  assign n4532 = n4287 & pi0841;
  assign n4533 = n4286 & pi0107;
  assign po0222 = n4532 | n4533;
  assign po0223 = n4304 & n4314;
  assign n4536 = n2515 & n4280;
  assign n4537 = n2503 & pi0314;
  assign n4538 = n2522 & n4537;
  assign n4539 = n4536 & n4538;
  assign n4540 = pi0219 & pi0299;
  assign n4541 = pi0199 & ~pi0299;
  assign n4542 = ~n4540 & ~n4541;
  assign po0224 = n4539 & ~n4542;
  assign n4544 = n2488 & ~pi0069;
  assign n4545 = n4544 & n4458;
  assign n4546 = n4545 & pi0314;
  assign n4547 = pi0083 & ~pi0103;
  assign po0225 = n4546 & n4547;
  assign n4549 = n3631 & n3545;
  assign n4550 = n3408 & n2931;
  assign n4551 = n2904 & pi0299;
  assign n4552 = n3463 & n4551;
  assign n4553 = ~n4550 & ~n4552;
  assign po0226 = n4549 & ~n4553;
  assign n4555 = pi0069 & ~pi0314;
  assign n4556 = ~n4555 & ~pi0071;
  assign po0227 = n4281 & ~n4556;
  assign n4558 = pi0024 & pi0070;
  assign n4559 = n3498 & n4558;
  assign n4560 = n3631 & n3468;
  assign n4561 = ~n4549 & ~n4560;
  assign n4562 = n3463 & n2710;
  assign n4563 = n4562 & pi0210;
  assign n4564 = n3408 & n2714;
  assign n4565 = n4564 & pi0198;
  assign n4566 = ~n4563 & ~n4565;
  assign n4567 = ~n4566 & pi0589;
  assign n4568 = ~n4561 & n4567;
  assign n4569 = n4568 & ~pi0593;
  assign n4570 = n3628 & n4358;
  assign n4571 = ~n4569 & ~n4570;
  assign po0228 = n4559 | ~n4571;
  assign n4573 = ~n4468 & pi0299;
  assign n4574 = ~n4472 & ~n4573;
  assign n4575 = n4539 & n4574;
  assign n4576 = ~n2462 & n4458;
  assign n4577 = n2447 & pi0085;
  assign n4578 = n4577 & n2473;
  assign n4579 = ~n2469 & n4578;
  assign n4580 = n4579 & pi0314;
  assign n4581 = n4576 & n4580;
  assign po0229 = n4575 | n4581;
  assign n4583 = n3541 & pi0088;
  assign n4584 = ~n2621 & n4583;
  assign n4585 = ~n4584 & ~pi0038;
  assign n4586 = n2620 & pi0072;
  assign n4587 = n4586 & pi0024;
  assign n4588 = n4585 & ~n4587;
  assign n4589 = ~n4588 & n2748;
  assign n4590 = n4549 & n3727;
  assign po0230 = n4589 | n4590;
  assign n4592 = n2891 & pi0073;
  assign n4593 = n4549 & ~n3467;
  assign n4594 = ~n4592 & ~n4593;
  assign n4595 = ~pi0314 & pi1050;
  assign n4596 = ~n4595 & ~pi0039;
  assign po0231 = ~n4594 & ~n4596;
  assign n4598 = n2668 & pi0479;
  assign n4599 = ~po0740 & ~n4598;
  assign n4600 = ~n4599 & ~pi0096;
  assign n4601 = ~pi0479 & ~pi0841;
  assign n4602 = ~n4601 & pi0096;
  assign n4603 = ~po0840 & ~n4602;
  assign n4604 = n2748 & n4603;
  assign n4605 = ~n4600 & n4604;
  assign n4606 = ~n2639 & n4605;
  assign n4607 = n4488 & pi0074;
  assign po0232 = n4606 | n4607;
  assign n4609 = n2656 & n2748;
  assign n4610 = n4488 & pi0075;
  assign po0233 = n4609 | n4610;
  assign n4612 = n3969 & n3920;
  assign n4613 = ~n4231 & ~n4612;
  assign n4614 = n3967 & n4613;
  assign n4615 = ~n3708 & pi0094;
  assign n4616 = ~n4614 & ~n4615;
  assign n4617 = ~n3969 & ~pi0094;
  assign n4618 = po0840 & ~n4617;
  assign n4619 = pi0094 & ~pi0252;
  assign n4620 = n4618 & ~n4619;
  assign n4621 = ~n4616 & ~n4620;
  assign po0234 = n2891 & n4621;
  assign n4623 = pi0077 & pi0314;
  assign n4624 = ~n2592 & ~n4623;
  assign po0235 = n3498 & n4624;
  assign po0236 = n3653 & pi0232;
  assign n4627 = n4142 ^ ~pi0079;
  assign n4628 = ~po0997 & ~n4627;
  assign n4629 = n4004 & ~n4628;
  assign n4630 = n4014 & ~pi0166;
  assign n4631 = n4630 & n4001;
  assign n4632 = ~pi0163 & pi0299;
  assign n4633 = ~n4631 & n4632;
  assign n4634 = ~n4081 & ~n4633;
  assign n4635 = n2574 & pi0153;
  assign n4636 = n3510 & n4635;
  assign n4637 = ~pi0040 & pi0095;
  assign n4638 = ~n4636 & ~n4637;
  assign n4639 = ~n4638 & pi0299;
  assign n4640 = n2675 & n4639;
  assign n4641 = pi0175 & ~pi0299;
  assign n4642 = ~n4640 & ~n4641;
  assign n4643 = ~n4634 & n4642;
  assign n4644 = pi0166 & pi0299;
  assign n4645 = pi0189 & ~pi0299;
  assign n4646 = ~n4644 & ~n4645;
  assign n4647 = n4003 & ~n4646;
  assign n4648 = ~n4647 & n3704;
  assign n4649 = pi0160 & pi0299;
  assign n4650 = pi0182 & ~pi0299;
  assign n4651 = ~n4649 & ~n4650;
  assign n4652 = n3506 & n4651;
  assign n4653 = n4648 & ~n4652;
  assign n4654 = ~n4095 & ~pi0184;
  assign n4655 = n4653 & ~n4654;
  assign n4656 = ~n4643 & n4655;
  assign n4657 = ~n4004 & n4656;
  assign n4658 = ~n4629 & ~n4657;
  assign n4659 = n4658 & ~pi0039;
  assign n4660 = ~n4042 & ~n4628;
  assign n4661 = n4025 & ~pi0189;
  assign n4662 = n4027 & ~pi0166;
  assign n4663 = ~n4661 & ~n4662;
  assign n4664 = n3545 & ~n4663;
  assign n4665 = n4025 & pi0179;
  assign n4666 = n4027 & pi0156;
  assign n4667 = ~n4665 & ~n4666;
  assign n4668 = n3468 & ~n4667;
  assign n4669 = ~n4664 & ~n4668;
  assign n4670 = ~n4669 & n3704;
  assign n4671 = n4039 & n4670;
  assign n4672 = ~n4671 & pi0039;
  assign n4673 = ~n4660 & n4672;
  assign n4674 = n2741 & n4014;
  assign n4675 = n4674 & ~pi0038;
  assign n4676 = ~n4673 & n4675;
  assign n4677 = ~n4659 & n4676;
  assign n4678 = ~n4046 & n4628;
  assign n4679 = ~n4678 & n4014;
  assign n4680 = pi0179 & ~pi0299;
  assign n4681 = pi0156 & pi0299;
  assign n4682 = ~n4680 & ~n4681;
  assign n4683 = n3704 & ~n4682;
  assign n4684 = n4046 & ~n4683;
  assign n4685 = n4679 & ~n4684;
  assign n4686 = ~n4685 & n2740;
  assign n4687 = ~n4686 & ~n2760;
  assign n4688 = ~n4059 & ~pi0040;
  assign n4689 = ~n4687 & n4688;
  assign n4690 = ~n4677 & n4689;
  assign n4691 = n4207 & n4208;
  assign n4692 = ~pi0162 & ~pi0197;
  assign n4693 = ~n4691 & ~n4692;
  assign n4694 = ~n4693 ^ ~pi0163;
  assign n4695 = ~n4694 & pi0299;
  assign n4696 = ~n4212 & n4213;
  assign n4697 = pi0140 & pi0145;
  assign n4698 = ~n4696 & ~n4697;
  assign n4699 = n4698 ^ ~pi0184;
  assign n4700 = ~n4699 & ~pi0299;
  assign n4701 = ~n4695 & ~n4700;
  assign n4702 = n4701 & n4071;
  assign n4703 = n2738 & ~n2739;
  assign n4704 = pi0187 & ~pi0299;
  assign n4705 = pi0147 & pi0299;
  assign n4706 = ~n4704 & ~n4705;
  assign n4707 = n3704 & ~n4706;
  assign n4708 = n4703 & ~n4707;
  assign n4709 = ~n4702 & ~n4708;
  assign n4710 = ~n4690 & n4709;
  assign n4711 = ~n4710 & ~po1038;
  assign n4712 = n3704 & pi0163;
  assign n4713 = n4138 & ~n4712;
  assign n4714 = ~n4138 & n4628;
  assign n4715 = ~n4713 & ~n4714;
  assign n4716 = n4715 & n4014;
  assign n4717 = ~n2745 & ~pi0040;
  assign n4718 = n4122 & n4717;
  assign n4719 = ~n4716 & n4718;
  assign n4720 = n4694 & n4071;
  assign n4721 = n3704 & pi0147;
  assign n4722 = ~n4721 & n2738;
  assign n4723 = ~n4720 & ~n4722;
  assign n4724 = po1038 & ~n4122;
  assign n4725 = ~n4723 & n4724;
  assign n4726 = ~n4719 & ~n4725;
  assign po0237 = n4711 | ~n4726;
  assign n4728 = ~n3479 & ~pi0063;
  assign n4729 = ~n4728 & n2804;
  assign n4730 = ~n3909 & ~pi0592;
  assign n4731 = n3890 & ~n4730;
  assign n4732 = ~pi0588 & ~pi0590;
  assign n4733 = n3888 & ~n4732;
  assign n4734 = ~n3949 & ~n3920;
  assign n4735 = n3920 & pi0590;
  assign n4736 = pi0098 & ~pi0592;
  assign n4737 = n4736 & pi1199;
  assign n4738 = ~n4735 & ~n4737;
  assign n4739 = ~n4734 & ~n4738;
  assign n4740 = ~n4733 & ~n4739;
  assign n4741 = n4731 & n4740;
  assign n4742 = n3625 & n3933;
  assign n4743 = ~n4741 & n4742;
  assign n4744 = ~n3698 & n4743;
  assign n4745 = ~n4729 & n4744;
  assign n4746 = n4731 & ~n4737;
  assign n4747 = ~n4746 & n3956;
  assign n4748 = ~n4745 & ~n4747;
  assign n4749 = ~n4748 & n3869;
  assign n4750 = ~n4749 & ~n3925;
  assign n4751 = n3927 & ~pi0080;
  assign po0238 = ~n4750 & n4751;
  assign n4753 = pi0081 & ~pi0314;
  assign n4754 = ~n4753 & ~pi0068;
  assign po0239 = ~n4426 & ~n4754;
  assign n4756 = ~pi0066 & ~pi0069;
  assign n4757 = ~n4555 & ~n4756;
  assign po0240 = n4281 & n4757;
  assign n4759 = ~pi0068 & pi0084;
  assign n4760 = n2506 & n4759;
  assign n4761 = n4576 & n4760;
  assign n4762 = n4547 & ~pi0314;
  assign n4763 = n4545 & n4762;
  assign po0241 = n4761 | n4763;
  assign n4765 = ~n4400 & pi0299;
  assign n4766 = ~n4380 & ~n4765;
  assign po0242 = n4539 & n4766;
  assign n4768 = n4579 & ~pi0314;
  assign n4769 = ~n4768 & ~pi0067;
  assign po0243 = n4576 & ~n4769;
  assign po0244 = n4560 & ~n4553;
  assign po0245 = n3489 & n4546;
  assign n4773 = n3412 & pi0104;
  assign n4774 = n4281 & n4773;
  assign n4775 = n4774 & n3920;
  assign n4776 = n3449 & pi0088;
  assign n4777 = n4286 & n4776;
  assign po0246 = n4775 | n4777;
  assign n4779 = pi0089 & pi0841;
  assign n4780 = ~pi0024 & pi0070;
  assign n4781 = ~n4779 & ~n4780;
  assign po0247 = n3498 & ~n4781;
  assign n4783 = n4592 & ~pi1050;
  assign n4784 = n4507 & pi0841;
  assign po0248 = n4783 | n4784;
  assign n4786 = ~n2650 & ~pi0024;
  assign n4787 = n3678 & ~n4786;
  assign n4788 = n4275 & n2650;
  assign n4789 = ~n4787 & ~n4788;
  assign n4790 = ~n4789 & n4445;
  assign n4791 = n3631 & n3728;
  assign po0249 = n4790 | n4791;
  assign n4793 = ~pi0039 & pi0092;
  assign n4794 = n4595 & n4793;
  assign n4795 = ~n3470 & ~n4794;
  assign po0250 = n2802 & ~n4795;
  assign n4797 = n3498 & n3375;
  assign n4798 = n2779 & n2825;
  assign n4799 = n4798 & ~pi1050;
  assign po0251 = n4797 | n4799;
  assign n4801 = n4282 & pi0049;
  assign n4802 = n3709 & ~po0840;
  assign n4803 = n4450 & n4802;
  assign po0252 = n4801 | n4803;
  assign n4805 = ~n4562 & ~n4564;
  assign n4806 = ~n4561 & ~n4805;
  assign n4807 = n4806 & ~n4567;
  assign n4808 = pi0089 & ~pi0332;
  assign n4809 = n4282 & n4808;
  assign n4810 = ~n4807 & ~n4809;
  assign n4811 = ~pi0032 & ~pi0040;
  assign n4812 = n2748 & n4811;
  assign n4813 = n4812 & pi0095;
  assign n4814 = n2623 & n4813;
  assign n4815 = n4814 & pi0024;
  assign po0253 = ~n4810 | n4815;
  assign n4817 = n4602 & ~pi0095;
  assign n4818 = ~n2648 & n4817;
  assign n4819 = ~pi0024 & pi0095;
  assign n4820 = n4819 & ~pi0096;
  assign n4821 = ~n4818 & ~n4820;
  assign n4822 = ~n4821 & n4812;
  assign po0254 = ~n2624 & n4822;
  assign n4824 = ~n2650 & ~n4599;
  assign n4825 = n4277 & n4824;
  assign n4826 = n2634 & n4825;
  assign n4827 = n4568 & pi0593;
  assign po0255 = n4826 | n4827;
  assign n4829 = ~n4592 & ~n4798;
  assign n4830 = pi0314 & pi1050;
  assign po0256 = ~n4829 & n4830;
  assign n4832 = n4354 & n3434;
  assign n4833 = n4832 ^ ~pi0099;
  assign n4834 = ~n4833 & n3695;
  assign n4835 = n4375 & pi0152;
  assign n4836 = n4835 & pi0161;
  assign n4837 = n4374 & pi0174;
  assign n4838 = n4837 & pi0144;
  assign n4839 = ~n4836 & ~n4838;
  assign n4840 = n4410 & ~n4839;
  assign po0257 = n4834 | n4840;
  assign n4842 = n2665 & ~n3412;
  assign n4843 = ~n4842 & pi0683;
  assign n4844 = ~n4843 & ~n3453;
  assign n4845 = n4844 & n3708;
  assign n4846 = ~n4845 & n3983;
  assign n4847 = ~n4846 & n3537;
  assign n4848 = po0840 & n3987;
  assign n4849 = ~n3986 & n4848;
  assign n4850 = ~n4847 & ~n4849;
  assign po0258 = n3536 & ~n4850;
  assign n4852 = n4354 ^ ~pi0101;
  assign n4853 = ~n4852 & n3695;
  assign n4854 = n4835 & ~pi0161;
  assign n4855 = n4837 & ~pi0144;
  assign n4856 = ~n4854 & ~n4855;
  assign n4857 = n4410 & ~n4856;
  assign po0259 = n4853 | n4857;
  assign po0260 = n4286 & pi0065;
  assign po0261 = n2891 & ~n3494;
  assign n4861 = n4774 & ~n3920;
  assign n4862 = n4449 & n4337;
  assign n4863 = n4862 & ~n4255;
  assign po0262 = n4861 | n4863;
  assign n4865 = n4433 & pi0106;
  assign n4866 = n4485 & ~pi0024;
  assign po0264 = n4865 | n4866;
  assign po0265 = n4529 & ~pi0999;
  assign n4869 = ~n4729 & ~n3629;
  assign n4870 = ~n4295 & pi0108;
  assign n4871 = ~n4870 & ~pi0098;
  assign n4872 = n4439 & ~n4871;
  assign po0266 = n4869 | n4872;
  assign po0267 = n4439 & n4623;
  assign n4875 = n3489 & n4459;
  assign n4876 = n4875 & pi0314;
  assign n4877 = n4862 & n4255;
  assign po0268 = n4876 | n4877;
  assign n4879 = n2748 & ~pi0024;
  assign n4880 = n4586 & n4879;
  assign n4881 = n4875 & ~pi0314;
  assign po0269 = n4880 | n4881;
  assign po0270 = ~pi0124 | pi0468;
  assign n4884 = n4354 & n3435;
  assign n4885 = n4884 ^ ~pi0113;
  assign po0271 = ~n4885 & n3695;
  assign n4887 = n4370 ^ ~pi0114;
  assign po0272 = ~n4887 & n3695;
  assign n4889 = n4369 & ~pi0116;
  assign n4890 = n4889 ^ ~pi0115;
  assign po0273 = ~n4890 & n3695;
  assign n4892 = n4369 ^ ~pi0116;
  assign po0274 = ~n4892 & n3695;
  assign n4894 = ~n4004 & n2743;
  assign n4895 = ~pi0038 & pi0039;
  assign n4896 = n4041 & n4895;
  assign n4897 = ~n2761 & ~pi0092;
  assign n4898 = ~n4896 & n4897;
  assign n4899 = n2738 & ~pi0054;
  assign n4900 = ~n2765 & ~n2741;
  assign n4901 = n4899 & ~n4900;
  assign n4902 = ~n4898 & n4901;
  assign n4903 = n2750 & n4902;
  assign n4904 = n4010 & ~pi0954;
  assign n4905 = n4904 & ~n4007;
  assign n4906 = n4142 & ~pi0079;
  assign n4907 = ~n4906 & pi0118;
  assign n4908 = ~n4905 & ~n4907;
  assign n4909 = ~n4908 & n2740;
  assign n4910 = ~n4903 & ~n4909;
  assign n4911 = ~n4894 & ~n4910;
  assign n4912 = pi0151 & pi0299;
  assign n4913 = pi0173 & ~pi0299;
  assign n4914 = ~n4912 & ~n4913;
  assign n4915 = n4081 & n4914;
  assign n4916 = ~n4915 & n3704;
  assign n4917 = ~n4916 & ~n3506;
  assign n4918 = ~n4099 & ~pi0150;
  assign n4919 = pi0073 & ~pi0168;
  assign n4920 = ~n4918 & ~n4919;
  assign n4921 = ~n4920 & pi0299;
  assign n4922 = ~pi0073 & pi0232;
  assign n4923 = n2627 & n4922;
  assign n4924 = n4099 & ~n4923;
  assign n4925 = ~pi0185 & ~pi0299;
  assign n4926 = ~n4924 & n4925;
  assign n4927 = n4104 & ~pi0190;
  assign n4928 = ~n4926 & ~n4927;
  assign n4929 = ~n4921 & n4928;
  assign n4930 = ~n4917 & n4929;
  assign n4931 = n4894 & ~n4930;
  assign n4932 = ~n4911 & ~n4931;
  assign n4933 = n3545 & pi0190;
  assign n4934 = n3468 & pi0178;
  assign n4935 = ~n4933 & ~n4934;
  assign n4936 = ~n4935 & n4025;
  assign n4937 = n3545 & pi0168;
  assign n4938 = n3468 & pi0157;
  assign n4939 = ~n4937 & ~n4938;
  assign n4940 = ~n4939 & n4027;
  assign n4941 = ~n4936 & ~n4940;
  assign n4942 = pi0039 & ~pi0092;
  assign n4943 = ~n4941 & n4942;
  assign n4944 = ~pi0178 & ~pi0299;
  assign n4945 = ~pi0157 & pi0299;
  assign n4946 = ~n4944 & ~n4945;
  assign n4947 = n4946 & n4793;
  assign n4948 = ~n4943 & ~n4947;
  assign n4949 = n3704 & ~pi0087;
  assign n4950 = n4039 & n4949;
  assign n4951 = ~n4948 & n4950;
  assign n4952 = ~n4951 & n4015;
  assign n4953 = ~n4932 & n4952;
  assign n4954 = ~n4693 & ~pi0163;
  assign n4955 = ~n4954 ^ ~pi0150;
  assign n4956 = ~n4955 & n4071;
  assign n4957 = n2738 & ~n4121;
  assign n4958 = n3704 & pi0165;
  assign n4959 = n4957 & ~n4958;
  assign n4960 = ~n4956 & ~n4959;
  assign n4961 = ~n4960 & ~n2885;
  assign n4962 = n4957 & ~n3704;
  assign n4963 = ~n4962 & n2745;
  assign n4964 = ~n4961 & n4963;
  assign n4965 = n4698 & ~pi0184;
  assign n4966 = ~n4965 ^ ~pi0185;
  assign n4967 = ~n4966 & n4071;
  assign n4968 = n4703 & ~pi0143;
  assign n4969 = ~n4967 & ~n4968;
  assign n4970 = ~n4969 & ~pi0299;
  assign n4971 = n4964 & ~n4970;
  assign n4972 = ~n4953 & n4971;
  assign n4973 = ~n4116 & n4908;
  assign n4974 = n3704 & pi0150;
  assign n4975 = n4116 & n4974;
  assign n4976 = ~n4973 & ~n4975;
  assign n4977 = n4976 & n4123;
  assign n4978 = n4960 & po1038;
  assign n4979 = ~n4977 & n4978;
  assign po0276 = ~n4972 & ~n4979;
  assign n4981 = n2592 & ~pi0109;
  assign n4982 = ~n4981 & n2569;
  assign n4983 = ~n3533 & n4982;
  assign n4984 = ~n2654 & n2574;
  assign n4985 = ~n4983 & n4984;
  assign n4986 = n2891 & ~n4985;
  assign n4987 = n3536 & ~n2847;
  assign n4988 = n4560 & ~n3723;
  assign n4989 = ~n4798 & ~n4988;
  assign n4990 = ~n4987 & n4989;
  assign po0288 = n4986 | ~n4990;
  assign n4992 = po0288 & ~pi0228;
  assign n4993 = pi0128 & pi0228;
  assign po0277 = n4992 | n4993;
  assign n4995 = ~n3738 & ~po1038;
  assign n4996 = ~n3702 & n4995;
  assign po0280 = n4996 | n3956;
  assign n4998 = ~pi0031 & ~pi0080;
  assign n4999 = n4998 & pi0818;
  assign n5000 = n4999 & pi1093;
  assign n5001 = pi0951 & pi0982;
  assign n5002 = n3923 & n5001;
  assign n5003 = n3927 & n5002;
  assign n5004 = ~n5000 & ~n5003;
  assign n5005 = n5004 & ~pi0120;
  assign po0278 = ~po0280 & ~n5005;
  assign n5007 = n4623 & ~pi0024;
  assign n5008 = ~n4088 & n5007;
  assign n5009 = n3498 & n5008;
  assign n5010 = n3461 & pi0181;
  assign n5011 = n3465 & pi0159;
  assign n5012 = ~n5010 & ~n5011;
  assign n5013 = n4304 & ~n5012;
  assign n5014 = ~n4361 & ~n4363;
  assign n5015 = ~n5014 & n3629;
  assign n5016 = ~n5015 & ~n3630;
  assign n5017 = ~n2885 & pi0163;
  assign n5018 = ~n5017 & pi0087;
  assign n5019 = n2885 & pi0184;
  assign n5020 = n5018 & ~n5019;
  assign n5021 = ~n2885 & ~pi0146;
  assign n5022 = ~po1038 & n2659;
  assign n5023 = pi0051 & ~pi0087;
  assign n5024 = ~n5022 & n5023;
  assign n5025 = ~n5021 & n5024;
  assign n5026 = ~n5020 & ~n5025;
  assign n5027 = n5016 & n5026;
  assign n5028 = ~n5013 & ~n5027;
  assign n5029 = ~n5009 & n5028;
  assign n5030 = ~n5029 & n3704;
  assign n5031 = pi0024 & pi0077;
  assign n5032 = ~n5031 & ~pi0086;
  assign n5033 = n5032 & ~n4623;
  assign n5034 = ~n5033 & ~pi0039;
  assign n5035 = n3625 & n5034;
  assign n5036 = n5035 & n2636;
  assign n5037 = n2562 & n5036;
  assign n5038 = n4683 & ~n5007;
  assign n5039 = n5037 & ~n5038;
  assign n5040 = ~n5039 & n3630;
  assign n5041 = n2562 & n5036;
  assign n5042 = pi0039 ^ ~pi0072;
  assign n5043 = n3626 & ~n5042;
  assign n5044 = n3546 & pi0039;
  assign n5045 = n5043 & ~n5044;
  assign n5046 = ~pi0134 & ~pi0135;
  assign n5047 = n5046 & ~pi0136;
  assign n5048 = n5047 & ~pi0130;
  assign n5049 = ~pi0126 & ~pi0132;
  assign n5050 = n5048 & n5049;
  assign n5051 = ~pi0125 & ~pi0133;
  assign n5052 = n5051 & ~pi0121;
  assign n5053 = ~n5050 & n5052;
  assign n5054 = ~n5051 & pi0121;
  assign n5055 = ~n5053 & ~n5054;
  assign n5056 = ~n5045 & n5055;
  assign n5057 = ~n5041 & ~n5056;
  assign n5058 = n5040 & ~n5057;
  assign po0279 = ~n5030 & ~n5058;
  assign n5060 = ~pi0090 & ~pi0111;
  assign n5061 = n5060 & ~pi0072;
  assign n5062 = n3487 & n5061;
  assign n5063 = n3498 & ~n5062;
  assign n5064 = pi0039 & ~pi0110;
  assign n5065 = n3637 & n5064;
  assign n5066 = ~n4413 & n3704;
  assign n5067 = ~pi0039 & pi0110;
  assign n5068 = n3412 & n5067;
  assign n5069 = po1057 & n5068;
  assign n5070 = ~n5066 & n5069;
  assign n5071 = ~n5065 & ~n5070;
  assign po0281 = ~n5063 & n5071;
  assign n5073 = ~n2621 & ~n5033;
  assign n5074 = ~n4586 & ~pi0039;
  assign n5075 = ~n5073 & n5074;
  assign n5076 = ~n5075 & n3624;
  assign n5077 = n3704 & ~pi0287;
  assign n5078 = n2900 & pi0158;
  assign n5079 = n5077 & n5078;
  assign n5080 = n3726 & ~n5079;
  assign n5081 = n2750 & ~n5080;
  assign n5082 = ~n2514 & ~pi0051;
  assign n5083 = n5082 & ~pi0152;
  assign n5084 = pi0051 & pi0172;
  assign n5085 = ~n5083 & ~n5084;
  assign n5086 = n5085 & pi0299;
  assign n5087 = ~n5086 & n3704;
  assign n5088 = ~n5081 & ~n5087;
  assign n5089 = n3623 & ~pi0072;
  assign n5090 = pi0180 & ~pi0287;
  assign n5091 = n3398 & n5090;
  assign n5092 = ~n5091 & pi0224;
  assign n5093 = ~pi0051 & pi0222;
  assign n5094 = n5093 & ~pi0223;
  assign n5095 = n2514 & n5094;
  assign n5096 = ~n5092 & n5095;
  assign n5097 = n5089 & n5096;
  assign n5098 = n5082 & ~pi0174;
  assign n5099 = pi0051 & pi0193;
  assign n5100 = ~n5099 & ~pi0299;
  assign n5101 = ~n5098 & n5100;
  assign n5102 = ~n5097 & n5101;
  assign n5103 = ~n5088 & ~n5102;
  assign n5104 = ~n5103 & pi0039;
  assign n5105 = n5076 & ~n5104;
  assign n5106 = n5087 & ~n5101;
  assign n5107 = ~pi0121 & ~pi0125;
  assign n5108 = n5050 & n5107;
  assign n5109 = ~pi0125 ^ ~pi0133;
  assign n5110 = ~n5108 & ~n5109;
  assign n5111 = ~n5110 & n3630;
  assign n5112 = ~n5106 & ~n5111;
  assign n5113 = ~n5105 & n5112;
  assign n5114 = n2740 & n4942;
  assign n5115 = ~n3548 & n5114;
  assign n5116 = n5089 & n5115;
  assign n5117 = ~n5103 & n5116;
  assign n5118 = ~n5117 & ~pi0087;
  assign n5119 = ~n5113 & n5118;
  assign n5120 = n3704 & pi0087;
  assign n5121 = pi0140 & ~pi0299;
  assign n5122 = ~n4175 & ~n5121;
  assign n5123 = n5120 & ~n5122;
  assign n5124 = ~n5123 & ~po1038;
  assign n5125 = ~n5119 & n5124;
  assign n5126 = n5037 & n2743;
  assign n5127 = n4152 & ~n5032;
  assign n5128 = pi0197 & pi0299;
  assign n5129 = pi0145 & ~pi0299;
  assign n5130 = ~n5128 & ~n5129;
  assign n5131 = n5032 & n5130;
  assign n5132 = ~n5127 & ~n5131;
  assign n5133 = n5132 & n3704;
  assign n5134 = n5126 & ~n5133;
  assign n5135 = ~n5085 & n4949;
  assign n5136 = n5120 & pi0162;
  assign n5137 = ~n5136 & po1038;
  assign n5138 = ~n5135 & n5137;
  assign n5139 = ~n5111 & n5138;
  assign n5140 = ~n5134 & ~n5139;
  assign po0282 = n5125 | ~n5140;
  assign n5142 = n5052 ^ ~pi0126;
  assign n5143 = n3630 & ~n5142;
  assign n5144 = ~n5050 & n5143;
  assign n5145 = ~n5126 & ~n5144;
  assign n5146 = ~n5145 & ~n5045;
  assign n5147 = n5077 & pi0160;
  assign n5148 = ~n5147 & n3465;
  assign n5149 = n5077 & pi0182;
  assign n5150 = ~n5149 & n3461;
  assign n5151 = ~n5148 & ~n5150;
  assign n5152 = n3628 & ~n5151;
  assign n5153 = pi0051 & pi0153;
  assign n5154 = ~pi0051 & ~pi0166;
  assign n5155 = ~n5153 & ~n5154;
  assign n5156 = n4949 & ~n5155;
  assign n5157 = n5156 & po1038;
  assign n5158 = ~n5157 & ~n3630;
  assign n5159 = ~n5152 & ~n5158;
  assign n5160 = ~n5146 & n5159;
  assign n5161 = n4946 & ~n5032;
  assign n5162 = ~n4183 & n5032;
  assign n5163 = ~n5161 & ~n5162;
  assign n5164 = n5126 & ~n5163;
  assign n5165 = n5082 & n4646;
  assign n5166 = n4641 & pi0051;
  assign n5167 = n5153 & pi0299;
  assign n5168 = ~n5166 & ~n5167;
  assign n5169 = ~n5165 & n5168;
  assign n5170 = ~po1038 & ~pi0087;
  assign n5171 = ~n5169 & n5170;
  assign n5172 = ~n2885 & ~pi0150;
  assign n5173 = ~po1038 & n4925;
  assign n5174 = ~n5173 & pi0087;
  assign n5175 = ~n5172 & n5174;
  assign n5176 = ~n5171 & ~n5175;
  assign n5177 = ~n5164 & n5176;
  assign n5178 = ~n5177 & n3704;
  assign po0283 = ~n5160 & ~n5178;
  assign n5180 = n3709 & pi0250;
  assign n5181 = ~n5180 & pi0127;
  assign n5182 = ~n5181 & pi0094;
  assign n5183 = n5180 & ~po0740;
  assign n5184 = n5182 & ~n5183;
  assign n5185 = ~n5184 & pi0129;
  assign po0284 = ~n4729 & n5185;
  assign n5187 = ~n3709 & ~pi0100;
  assign n5188 = ~n5187 & ~pi0250;
  assign n5189 = ~n5188 & pi0129;
  assign n5190 = ~n5189 & ~n2737;
  assign n5191 = n5188 & ~po0740;
  assign n5192 = n5190 & ~n5191;
  assign n5193 = ~n2804 & ~n5192;
  assign po0286 = n2891 | n5193;
  assign n5195 = n2927 & pi0140;
  assign n5196 = n2900 & n4175;
  assign n5197 = ~n5195 & ~n5196;
  assign n5198 = ~n5197 & n5077;
  assign n5199 = ~n5198 & n3726;
  assign n5200 = n2750 & ~n5199;
  assign n5201 = ~n5200 & pi0039;
  assign n5202 = n5076 & ~n5201;
  assign n5203 = n5052 & n5049;
  assign n5204 = n5203 & ~pi0130;
  assign n5205 = n5204 & ~n5047;
  assign n5206 = ~n5203 & pi0130;
  assign n5207 = ~n5206 & n2514;
  assign n5208 = ~n5205 & n5207;
  assign n5209 = ~n5116 & n5208;
  assign n5210 = n4067 & ~n2514;
  assign n5211 = ~n5209 & ~n5210;
  assign n5212 = n5211 & n5170;
  assign n5213 = ~n5202 & n5212;
  assign n5214 = ~n2514 & n3704;
  assign n5215 = n5214 & pi0169;
  assign n5216 = po1038 & ~n5120;
  assign n5217 = ~n5215 & n5216;
  assign n5218 = ~n5208 & n5217;
  assign n5219 = ~n5213 & ~n5218;
  assign n5220 = ~n5219 & ~pi0051;
  assign n5221 = ~n2885 & ~pi0167;
  assign n5222 = ~po1038 & n4190;
  assign n5223 = ~n5222 & n3704;
  assign n5224 = ~n5221 & n5223;
  assign n5225 = ~n5224 & pi0087;
  assign po0287 = n5220 | n5225;
  assign n5227 = n3628 & ~n3548;
  assign n5228 = ~n5227 & n3630;
  assign n5229 = ~n5041 & n5228;
  assign n5230 = n3704 & ~n4651;
  assign n5231 = ~pi0024 & pi0077;
  assign n5232 = ~n5230 & n5231;
  assign n5233 = n3464 & pi0149;
  assign n5234 = n2927 & pi0183;
  assign n5235 = ~n5233 & ~n5234;
  assign n5236 = ~n5232 & ~n5235;
  assign n5237 = n5236 & n5077;
  assign n5238 = n5237 & n3630;
  assign n5239 = ~n5229 & ~n5238;
  assign n5240 = ~n5048 & n5203;
  assign n5241 = n5052 & ~pi0126;
  assign n5242 = ~n5241 & pi0132;
  assign n5243 = ~n5240 & ~n5242;
  assign n5244 = ~n5045 & ~n5243;
  assign n5245 = ~n5239 & ~n5244;
  assign n5246 = n5126 & ~n5232;
  assign n5247 = n2885 & ~pi0190;
  assign n5248 = ~n5247 & ~n2514;
  assign n5249 = ~n2885 & ~pi0168;
  assign n5250 = n5248 & ~n5249;
  assign n5251 = ~n5250 & n3629;
  assign n5252 = n2885 & pi0173;
  assign n5253 = ~n5252 & n5023;
  assign n5254 = ~n2885 & pi0151;
  assign n5255 = n5253 & ~n5254;
  assign n5256 = ~n2885 & pi0164;
  assign n5257 = ~po1038 & n4018;
  assign n5258 = ~n5257 & pi0087;
  assign n5259 = ~n5256 & n5258;
  assign n5260 = ~n5259 & n3704;
  assign n5261 = ~n5255 & n5260;
  assign n5262 = ~n5251 & n5261;
  assign n5263 = ~n5246 & ~n5262;
  assign po0289 = ~n5245 & n5263;
  assign n5265 = n2927 & pi0145;
  assign n5266 = n2900 & n5128;
  assign n5267 = ~n5265 & ~n5266;
  assign n5268 = ~n5267 & n5077;
  assign n5269 = n3726 & ~pi0072;
  assign n5270 = ~n5268 & n5269;
  assign n5271 = ~n5270 & ~n5042;
  assign n5272 = ~n4729 & n5271;
  assign n5273 = n3973 & ~pi0086;
  assign n5274 = ~n5273 & ~n4050;
  assign n5275 = n5126 & ~n5274;
  assign n5276 = ~n5108 & ~pi0133;
  assign n5277 = n5228 & ~n5276;
  assign n5278 = ~n2885 & ~pi0149;
  assign n5279 = ~n5278 & n5120;
  assign n5280 = n2885 & ~pi0183;
  assign n5281 = n5279 & ~n5280;
  assign n5282 = ~n5277 & ~n5281;
  assign n5283 = ~n5126 & ~n5282;
  assign n5284 = ~n5275 & ~n5283;
  assign po0290 = ~n5272 & n5284;
  assign n5286 = ~n5041 & n3629;
  assign n5287 = n5204 & ~pi0136;
  assign n5288 = n5287 & ~pi0135;
  assign n5289 = ~n5288 & pi0134;
  assign n5290 = ~n5045 & ~n5289;
  assign n5291 = n2927 & pi0186;
  assign n5292 = n2900 & n4017;
  assign n5293 = ~n5291 & ~n5292;
  assign n5294 = ~n5293 & n5077;
  assign n5295 = n5269 & ~n5294;
  assign n5296 = n5043 & ~n5295;
  assign n5297 = ~n5290 & ~n5296;
  assign n5298 = ~n5297 & n2514;
  assign n5299 = ~n2885 & ~pi0171;
  assign n5300 = n2885 & ~pi0192;
  assign n5301 = ~n5299 & ~n5300;
  assign n5302 = n5301 & n5214;
  assign n5303 = ~n5298 & ~n5302;
  assign po0291 = n5286 & n5303;
  assign n5305 = n3464 & pi0150;
  assign n5306 = n2927 & pi0185;
  assign n5307 = ~n5305 & ~n5306;
  assign n5308 = ~n5307 & n5077;
  assign n5309 = n5227 & ~n5308;
  assign n5310 = ~n5309 & n2514;
  assign n5311 = n5288 & pi0134;
  assign n5312 = ~n5287 & pi0135;
  assign n5313 = ~n5311 & ~n5312;
  assign n5314 = ~n5045 & ~n5313;
  assign n5315 = n5310 & ~n5314;
  assign n5316 = ~n2885 & ~pi0170;
  assign n5317 = n2885 & ~pi0194;
  assign n5318 = ~n5316 & ~n5317;
  assign n5319 = n5318 & n5214;
  assign n5320 = ~n5315 & ~n5319;
  assign po0292 = n5286 & n5320;
  assign n5322 = n3464 & pi0163;
  assign n5323 = n2927 & pi0184;
  assign n5324 = ~n5322 & ~n5323;
  assign n5325 = ~n5324 & n5077;
  assign n5326 = ~n5325 & n3726;
  assign n5327 = n5089 & ~n5326;
  assign n5328 = n2514 & pi0039;
  assign n5329 = ~n5327 & n5328;
  assign n5330 = n3704 & ~n4197;
  assign n5331 = ~n5330 & ~n2514;
  assign n5332 = n3625 & ~n5331;
  assign n5333 = ~n5329 & n5332;
  assign n5334 = ~n5075 & n5333;
  assign n5335 = ~n2885 & ~pi0148;
  assign n5336 = ~n5335 & n5214;
  assign n5337 = n2885 & ~pi0141;
  assign n5338 = n5336 & ~n5337;
  assign n5339 = n5287 & ~n5046;
  assign n5340 = ~n5204 & pi0136;
  assign n5341 = ~n5340 & n2514;
  assign n5342 = ~n5339 & n5341;
  assign n5343 = ~n5338 & ~n5342;
  assign n5344 = ~n5227 & ~n5343;
  assign n5345 = ~n5344 & n3629;
  assign po0293 = ~n5334 & n5345;
  assign n5347 = n4411 & ~pi0198;
  assign n5348 = n4412 & ~pi0210;
  assign n5349 = ~n5347 & ~n5348;
  assign n5350 = n3704 & pi0039;
  assign n5351 = ~n5349 & n5350;
  assign n5352 = ~n4378 & n5351;
  assign n5353 = ~pi0039 & pi0137;
  assign po0294 = n5352 | n5353;
  assign n5355 = ~n4000 & ~pi0039;
  assign n5356 = n4039 & n3470;
  assign n5357 = ~n5355 & ~n5356;
  assign n5358 = n2745 & n2741;
  assign n5359 = ~n5357 & n5358;
  assign n5360 = n2788 & n4123;
  assign n5361 = ~n5359 & n5360;
  assign n5362 = n5361 & n4594;
  assign n5363 = n4904 & n4006;
  assign n5364 = n5363 & ~n4005;
  assign n5365 = n4904 & ~pi0139;
  assign n5366 = ~n5365 & pi0138;
  assign n5367 = ~n5364 & ~n5366;
  assign n5368 = n5362 & ~n5367;
  assign n5369 = ~n4594 & ~n5330;
  assign po0295 = n5368 | n5369;
  assign n5371 = n4904 ^ ~pi0139;
  assign n5372 = ~n5371 & ~n4007;
  assign n5373 = n5362 & n5372;
  assign n5374 = ~n4594 & ~n4067;
  assign po0296 = n5373 | n5374;
  assign n5376 = n4302 & ~po0950;
  assign n5377 = n4224 & ~pi0841;
  assign n5378 = n2601 & n5377;
  assign n5379 = ~pi0045 & ~pi0047;
  assign n5380 = n5379 & ~pi0102;
  assign n5381 = n5380 & ~n4294;
  assign n5382 = ~n5378 & n5381;
  assign n5383 = ~n2506 & ~pi0047;
  assign n5384 = ~n5383 & ~pi0252;
  assign n5385 = ~n5382 & ~n5384;
  assign n5386 = ~n5385 & ~pi0040;
  assign n5387 = ~n5376 & n5386;
  assign n5388 = n4585 & n5387;
  assign n5389 = ~n4729 & ~n5388;
  assign n5390 = ~n4561 & ~n3723;
  assign n5391 = ~n4311 & ~pi0287;
  assign n5392 = ~n5391 & ~pi0120;
  assign n5393 = ~n3432 & ~n5392;
  assign n5394 = n3631 & n5393;
  assign n5395 = ~n5390 & ~n5394;
  assign n5396 = ~n5389 & n5395;
  assign n5397 = ~n5396 & n3923;
  assign n5398 = n3923 & pi0832;
  assign n5399 = ~n5397 & ~n5398;
  assign n5400 = n5399 & ~pi0140;
  assign n5401 = ~pi0618 ^ ~pi1154;
  assign n5402 = n5401 & pi0781;
  assign n5403 = ~pi0609 ^ ~pi1155;
  assign n5404 = n5403 & pi0785;
  assign n5405 = ~n5402 & ~n5404;
  assign n5406 = ~pi0630 ^ ~pi1157;
  assign n5407 = n5406 & pi0787;
  assign n5408 = pi0626 ^ ~pi1158;
  assign n5409 = ~n5408 & pi0788;
  assign n5410 = ~n5407 & ~n5409;
  assign n5411 = n5405 & n5410;
  assign n5412 = pi0644 ^ ~pi1160;
  assign n5413 = ~n5412 & pi0790;
  assign n5414 = ~n5413 & pi0603;
  assign n5415 = n5411 & n5414;
  assign n5416 = pi0619 ^ ~pi1159;
  assign n5417 = ~n5416 & pi0789;
  assign n5418 = pi0608 ^ ~pi1153;
  assign n5419 = ~n5418 & pi0778;
  assign n5420 = ~n5417 & ~n5419;
  assign n5421 = ~pi0629 ^ ~pi1156;
  assign n5422 = n5421 & pi0792;
  assign n5423 = n5420 & ~n5422;
  assign n5424 = n5415 & n5423;
  assign n5425 = pi0621 & pi1091;
  assign n5426 = n5424 & ~n5425;
  assign n5427 = pi0715 ^ ~pi1160;
  assign n5428 = ~n5427 & pi0790;
  assign n5429 = ~pi0641 ^ ~pi1158;
  assign n5430 = n5429 & pi0788;
  assign n5431 = ~n5428 & ~n5430;
  assign n5432 = ~pi0625 ^ ~pi1153;
  assign n5433 = n5432 & pi0778;
  assign n5434 = n5431 & ~n5433;
  assign n5435 = pi0660 ^ ~pi1155;
  assign n5436 = ~n5435 & pi0785;
  assign n5437 = ~n5436 & pi0680;
  assign n5438 = ~pi0627 ^ ~pi1154;
  assign n5439 = n5438 & pi0781;
  assign n5440 = ~pi0647 ^ ~pi1157;
  assign n5441 = n5440 & pi0787;
  assign n5442 = ~n5439 & ~n5441;
  assign n5443 = n5437 & n5442;
  assign n5444 = n5434 & n5443;
  assign n5445 = pi0628 ^ ~pi1156;
  assign n5446 = ~n5445 & pi0792;
  assign n5447 = pi0648 ^ ~pi1159;
  assign n5448 = ~n5447 & pi0789;
  assign n5449 = ~n5446 & ~n5448;
  assign n5450 = n5444 & n5449;
  assign n5451 = pi0665 & pi1091;
  assign n5452 = n5450 & ~n5451;
  assign n5453 = ~n5426 & n5452;
  assign n5454 = n5453 & ~pi0738;
  assign n5455 = n5426 & ~pi0761;
  assign n5456 = ~n5454 & ~n5455;
  assign n5457 = ~n5399 & ~n5456;
  assign po0297 = n5400 | n5457;
  assign n5459 = n5399 & ~pi0141;
  assign n5460 = n5453 & pi0706;
  assign n5461 = n5426 & pi0749;
  assign n5462 = ~n5460 & ~n5461;
  assign n5463 = ~n5399 & ~n5462;
  assign po0298 = n5459 | n5463;
  assign n5465 = n5453 & pi0735;
  assign n5466 = n5426 & pi0743;
  assign n5467 = ~n5465 & ~n5466;
  assign n5468 = ~n5399 & n5467;
  assign n5469 = n5399 & ~pi0142;
  assign po0299 = ~n5468 & ~n5469;
  assign n5471 = n5399 & ~pi0143;
  assign n5472 = n5453 & pi0687;
  assign n5473 = n5426 & ~pi0774;
  assign n5474 = ~n5472 & ~n5473;
  assign n5475 = ~n5399 & ~n5474;
  assign po0300 = n5471 | n5475;
  assign n5477 = n5453 & pi0736;
  assign n5478 = n5426 & pi0758;
  assign n5479 = ~n5477 & ~n5478;
  assign n5480 = ~n5399 & n5479;
  assign n5481 = n5399 & ~pi0144;
  assign po0301 = ~n5480 & ~n5481;
  assign n5483 = n5399 & ~pi0145;
  assign n5484 = n5453 & ~pi0698;
  assign n5485 = n5426 & ~pi0767;
  assign n5486 = ~n5484 & ~n5485;
  assign n5487 = ~n5399 & ~n5486;
  assign po0302 = n5483 | n5487;
  assign n5489 = pi0907 & ~pi0947;
  assign n5490 = n5489 & pi0735;
  assign n5491 = pi0743 & pi0947;
  assign n5492 = ~n5490 & ~n5491;
  assign n5493 = ~n5399 & n5492;
  assign n5494 = n5399 & ~pi0146;
  assign po0303 = ~n5493 & ~n5494;
  assign n5496 = n5399 & ~pi0147;
  assign n5497 = n5489 & pi0726;
  assign n5498 = ~pi0770 & pi0947;
  assign n5499 = ~n5497 & ~n5498;
  assign n5500 = ~n5399 & ~n5499;
  assign po0304 = n5496 | n5500;
  assign n5502 = n5399 & ~pi0148;
  assign n5503 = n5489 & pi0706;
  assign n5504 = pi0749 & pi0947;
  assign n5505 = ~n5503 & ~n5504;
  assign n5506 = ~n5399 & ~n5505;
  assign po0305 = n5502 | n5506;
  assign n5508 = ~n3422 & ~n5392;
  assign n5509 = n3420 & n3721;
  assign n5510 = n3720 & ~n4040;
  assign n5511 = ~n5509 & ~n5510;
  assign n5512 = ~n5508 & n5511;
  assign n5513 = n3631 & ~n5512;
  assign n5514 = ~n5389 & ~n5513;
  assign n5515 = ~n5514 & n3923;
  assign n5516 = ~n5515 & ~n5398;
  assign n5517 = n5489 & ~pi0725;
  assign n5518 = ~pi0755 & pi0947;
  assign n5519 = ~n5517 & ~n5518;
  assign n5520 = ~n5516 & ~n5519;
  assign n5521 = n5399 & ~pi0149;
  assign po0306 = n5520 | n5521;
  assign n5523 = n5489 & ~pi0701;
  assign n5524 = ~pi0751 & pi0947;
  assign n5525 = ~n5523 & ~n5524;
  assign n5526 = ~n5516 & ~n5525;
  assign n5527 = n5399 & ~pi0150;
  assign po0307 = n5526 | n5527;
  assign n5529 = n5399 & ~pi0151;
  assign n5530 = n5489 & ~pi0723;
  assign n5531 = ~pi0745 & pi0947;
  assign n5532 = ~n5530 & ~n5531;
  assign n5533 = ~n5399 & ~n5532;
  assign po0308 = n5529 | n5533;
  assign n5535 = n5489 & pi0696;
  assign n5536 = pi0759 & pi0947;
  assign n5537 = ~n5535 & ~n5536;
  assign n5538 = ~n5399 & n5537;
  assign n5539 = n5399 & ~pi0152;
  assign po0309 = ~n5538 & ~n5539;
  assign n5541 = n5399 & ~pi0153;
  assign n5542 = n5489 & pi0700;
  assign n5543 = pi0766 & pi0947;
  assign n5544 = ~n5542 & ~n5543;
  assign n5545 = ~n5399 & ~n5544;
  assign po0310 = n5541 | n5545;
  assign n5547 = n5489 & ~pi0704;
  assign n5548 = ~pi0742 & pi0947;
  assign n5549 = ~n5547 & ~n5548;
  assign n5550 = ~n5516 & ~n5549;
  assign n5551 = n5399 & ~pi0154;
  assign po0311 = n5550 | n5551;
  assign n5553 = n5489 & ~pi0686;
  assign n5554 = ~pi0757 & pi0947;
  assign n5555 = ~n5553 & ~n5554;
  assign n5556 = ~n5516 & ~n5555;
  assign n5557 = n5399 & ~pi0155;
  assign po0312 = n5556 | n5557;
  assign n5559 = n5489 & ~pi0724;
  assign n5560 = ~pi0741 & pi0947;
  assign n5561 = ~n5559 & ~n5560;
  assign n5562 = ~n5516 & ~n5561;
  assign n5563 = n5399 & ~pi0156;
  assign po0313 = n5562 | n5563;
  assign n5565 = n5399 & ~pi0157;
  assign n5566 = n5489 & ~pi0688;
  assign n5567 = ~pi0760 & pi0947;
  assign n5568 = ~n5566 & ~n5567;
  assign n5569 = ~n5399 & ~n5568;
  assign po0314 = n5565 | n5569;
  assign n5571 = n5489 & ~pi0702;
  assign n5572 = ~pi0753 & pi0947;
  assign n5573 = ~n5571 & ~n5572;
  assign n5574 = ~n5516 & ~n5573;
  assign n5575 = n5399 & ~pi0158;
  assign po0315 = n5574 | n5575;
  assign n5577 = n5399 & ~pi0159;
  assign n5578 = n5489 & ~pi0709;
  assign n5579 = ~pi0754 & pi0947;
  assign n5580 = ~n5578 & ~n5579;
  assign n5581 = ~n5399 & ~n5580;
  assign po0316 = n5577 | n5581;
  assign n5583 = n5399 & ~pi0160;
  assign n5584 = n5489 & ~pi0734;
  assign n5585 = ~pi0756 & pi0947;
  assign n5586 = ~n5584 & ~n5585;
  assign n5587 = ~n5399 & ~n5586;
  assign po0317 = n5583 | n5587;
  assign n5589 = n5489 & pi0736;
  assign n5590 = pi0758 & pi0947;
  assign n5591 = ~n5589 & ~n5590;
  assign n5592 = ~n5399 & n5591;
  assign n5593 = n5399 & ~pi0161;
  assign po0318 = ~n5592 & ~n5593;
  assign n5595 = n5399 & ~pi0162;
  assign n5596 = n5489 & ~pi0738;
  assign n5597 = ~pi0761 & pi0947;
  assign n5598 = ~n5596 & ~n5597;
  assign n5599 = ~n5399 & ~n5598;
  assign po0319 = n5595 | n5599;
  assign n5601 = n5399 & ~pi0163;
  assign n5602 = n5489 & ~pi0737;
  assign n5603 = ~pi0777 & pi0947;
  assign n5604 = ~n5602 & ~n5603;
  assign n5605 = ~n5399 & ~n5604;
  assign po0320 = n5601 | n5605;
  assign n5607 = n5399 & ~pi0164;
  assign n5608 = n5489 & pi0703;
  assign n5609 = ~pi0752 & pi0947;
  assign n5610 = ~n5608 & ~n5609;
  assign n5611 = ~n5399 & ~n5610;
  assign po0321 = n5607 | n5611;
  assign n5613 = n5489 & pi0687;
  assign n5614 = ~pi0774 & pi0947;
  assign n5615 = ~n5613 & ~n5614;
  assign n5616 = ~n5516 & ~n5615;
  assign n5617 = n5399 & ~pi0165;
  assign po0322 = n5616 | n5617;
  assign n5619 = n5489 & pi0727;
  assign n5620 = pi0772 & pi0947;
  assign n5621 = ~n5619 & ~n5620;
  assign n5622 = ~n5399 & n5621;
  assign n5623 = n5399 & ~pi0166;
  assign po0323 = ~n5622 & ~n5623;
  assign n5625 = n5399 & ~pi0167;
  assign n5626 = n5489 & pi0705;
  assign n5627 = ~pi0768 & pi0947;
  assign n5628 = ~n5626 & ~n5627;
  assign n5629 = ~n5399 & ~n5628;
  assign po0324 = n5625 | n5629;
  assign n5631 = n5399 & ~pi0168;
  assign n5632 = n5489 & pi0699;
  assign n5633 = pi0763 & pi0947;
  assign n5634 = ~n5632 & ~n5633;
  assign n5635 = ~n5399 & ~n5634;
  assign po0325 = n5631 | n5635;
  assign n5637 = n5399 & ~pi0169;
  assign n5638 = n5489 & pi0729;
  assign n5639 = pi0746 & pi0947;
  assign n5640 = ~n5638 & ~n5639;
  assign n5641 = ~n5399 & ~n5640;
  assign po0326 = n5637 | n5641;
  assign n5643 = n5399 & ~pi0170;
  assign n5644 = n5489 & pi0730;
  assign n5645 = pi0748 & pi0947;
  assign n5646 = ~n5644 & ~n5645;
  assign n5647 = ~n5399 & ~n5646;
  assign po0327 = n5643 | n5647;
  assign n5649 = n5399 & ~pi0171;
  assign n5650 = n5489 & pi0691;
  assign n5651 = pi0764 & pi0947;
  assign n5652 = ~n5650 & ~n5651;
  assign n5653 = ~n5399 & ~n5652;
  assign po0328 = n5649 | n5653;
  assign n5655 = n5399 & ~pi0172;
  assign n5656 = n5489 & pi0690;
  assign n5657 = pi0739 & pi0947;
  assign n5658 = ~n5656 & ~n5657;
  assign n5659 = ~n5399 & ~n5658;
  assign po0329 = n5655 | n5659;
  assign n5661 = n5399 & ~pi0173;
  assign n5662 = n5453 & ~pi0723;
  assign n5663 = n5426 & ~pi0745;
  assign n5664 = ~n5662 & ~n5663;
  assign n5665 = ~n5399 & ~n5664;
  assign po0330 = n5661 | n5665;
  assign n5667 = n5453 & pi0696;
  assign n5668 = n5426 & pi0759;
  assign n5669 = ~n5667 & ~n5668;
  assign n5670 = ~n5399 & n5669;
  assign n5671 = n5399 & ~pi0174;
  assign po0331 = ~n5670 & ~n5671;
  assign n5673 = n5399 & ~pi0175;
  assign n5674 = n5453 & pi0700;
  assign n5675 = n5426 & pi0766;
  assign n5676 = ~n5674 & ~n5675;
  assign n5677 = ~n5399 & ~n5676;
  assign po0332 = n5673 | n5677;
  assign n5679 = n5399 & ~pi0176;
  assign n5680 = n5453 & ~pi0704;
  assign n5681 = n5426 & ~pi0742;
  assign n5682 = ~n5680 & ~n5681;
  assign n5683 = ~n5399 & ~n5682;
  assign po0333 = n5679 | n5683;
  assign n5685 = n5399 & ~pi0177;
  assign n5686 = n5453 & ~pi0686;
  assign n5687 = n5426 & ~pi0757;
  assign n5688 = ~n5686 & ~n5687;
  assign n5689 = ~n5399 & ~n5688;
  assign po0334 = n5685 | n5689;
  assign n5691 = n5399 & ~pi0178;
  assign n5692 = n5453 & ~pi0688;
  assign n5693 = n5426 & ~pi0760;
  assign n5694 = ~n5692 & ~n5693;
  assign n5695 = ~n5399 & ~n5694;
  assign po0335 = n5691 | n5695;
  assign n5697 = n5399 & ~pi0179;
  assign n5698 = n5453 & ~pi0724;
  assign n5699 = n5426 & ~pi0741;
  assign n5700 = ~n5698 & ~n5699;
  assign n5701 = ~n5399 & ~n5700;
  assign po0336 = n5697 | n5701;
  assign n5703 = n5399 & ~pi0180;
  assign n5704 = n5453 & ~pi0702;
  assign n5705 = n5426 & ~pi0753;
  assign n5706 = ~n5704 & ~n5705;
  assign n5707 = ~n5399 & ~n5706;
  assign po0337 = n5703 | n5707;
  assign n5709 = n5399 & ~pi0181;
  assign n5710 = n5453 & ~pi0709;
  assign n5711 = n5426 & ~pi0754;
  assign n5712 = ~n5710 & ~n5711;
  assign n5713 = ~n5399 & ~n5712;
  assign po0338 = n5709 | n5713;
  assign n5715 = n5399 & ~pi0182;
  assign n5716 = n5453 & ~pi0734;
  assign n5717 = n5426 & ~pi0756;
  assign n5718 = ~n5716 & ~n5717;
  assign n5719 = ~n5399 & ~n5718;
  assign po0339 = n5715 | n5719;
  assign n5721 = n5399 & ~pi0183;
  assign n5722 = n5453 & ~pi0725;
  assign n5723 = n5426 & ~pi0755;
  assign n5724 = ~n5722 & ~n5723;
  assign n5725 = ~n5399 & ~n5724;
  assign po0340 = n5721 | n5725;
  assign n5727 = n5399 & ~pi0184;
  assign n5728 = n5453 & ~pi0737;
  assign n5729 = n5426 & ~pi0777;
  assign n5730 = ~n5728 & ~n5729;
  assign n5731 = ~n5399 & ~n5730;
  assign po0341 = n5727 | n5731;
  assign n5733 = n5399 & ~pi0185;
  assign n5734 = n5453 & ~pi0701;
  assign n5735 = n5426 & ~pi0751;
  assign n5736 = ~n5734 & ~n5735;
  assign n5737 = ~n5399 & ~n5736;
  assign po0342 = n5733 | n5737;
  assign n5739 = n5399 & ~pi0186;
  assign n5740 = n5453 & pi0703;
  assign n5741 = n5426 & ~pi0752;
  assign n5742 = ~n5740 & ~n5741;
  assign n5743 = ~n5399 & ~n5742;
  assign po0343 = n5739 | n5743;
  assign n5745 = n5399 & ~pi0187;
  assign n5746 = n5453 & pi0726;
  assign n5747 = n5426 & ~pi0770;
  assign n5748 = ~n5746 & ~n5747;
  assign n5749 = ~n5399 & ~n5748;
  assign po0344 = n5745 | n5749;
  assign n5751 = n5399 & ~pi0188;
  assign n5752 = n5453 & pi0705;
  assign n5753 = n5426 & ~pi0768;
  assign n5754 = ~n5752 & ~n5753;
  assign n5755 = ~n5399 & ~n5754;
  assign po0345 = n5751 | n5755;
  assign n5757 = n5453 & pi0727;
  assign n5758 = n5426 & pi0772;
  assign n5759 = ~n5757 & ~n5758;
  assign n5760 = ~n5399 & n5759;
  assign n5761 = n5399 & ~pi0189;
  assign po0346 = ~n5760 & ~n5761;
  assign n5763 = n5399 & ~pi0190;
  assign n5764 = n5453 & pi0699;
  assign n5765 = n5426 & pi0763;
  assign n5766 = ~n5764 & ~n5765;
  assign n5767 = ~n5399 & ~n5766;
  assign po0347 = n5763 | n5767;
  assign n5769 = n5399 & ~pi0191;
  assign n5770 = n5453 & pi0729;
  assign n5771 = n5426 & pi0746;
  assign n5772 = ~n5770 & ~n5771;
  assign n5773 = ~n5399 & ~n5772;
  assign po0348 = n5769 | n5773;
  assign n5775 = n5399 & ~pi0192;
  assign n5776 = n5453 & pi0691;
  assign n5777 = n5426 & pi0764;
  assign n5778 = ~n5776 & ~n5777;
  assign n5779 = ~n5399 & ~n5778;
  assign po0349 = n5775 | n5779;
  assign n5781 = n5399 & ~pi0193;
  assign n5782 = n5453 & pi0690;
  assign n5783 = n5426 & pi0739;
  assign n5784 = ~n5782 & ~n5783;
  assign n5785 = ~n5399 & ~n5784;
  assign po0350 = n5781 | n5785;
  assign n5787 = n5399 & ~pi0194;
  assign n5788 = n5453 & pi0730;
  assign n5789 = n5426 & pi0748;
  assign n5790 = ~n5788 & ~n5789;
  assign n5791 = ~n5399 & ~n5790;
  assign po0351 = n5787 | n5791;
  assign n5793 = n5363 & ~pi0196;
  assign n5794 = ~n5793 & pi0195;
  assign n5795 = n5362 & n5794;
  assign n5796 = pi0192 & ~pi0299;
  assign n5797 = pi0171 & pi0299;
  assign n5798 = ~n5796 & ~n5797;
  assign n5799 = n3704 & ~n5798;
  assign n5800 = ~n4594 & ~n5799;
  assign po0352 = n5795 | n5800;
  assign n5802 = n5793 & pi0195;
  assign n5803 = ~n5363 & pi0196;
  assign n5804 = ~n5802 & ~n5803;
  assign n5805 = n5362 & ~n5804;
  assign n5806 = pi0194 & ~pi0299;
  assign n5807 = pi0170 & pi0299;
  assign n5808 = ~n5806 & ~n5807;
  assign n5809 = n3704 & ~n5808;
  assign n5810 = ~n4594 & ~n5809;
  assign po0353 = n5805 | n5810;
  assign n5812 = n5399 & ~pi0197;
  assign n5813 = n5489 & ~pi0698;
  assign n5814 = ~pi0767 & pi0947;
  assign n5815 = ~n5813 & ~n5814;
  assign n5816 = ~n5399 & ~n5815;
  assign po0354 = n5812 | n5816;
  assign n5818 = ~n5397 & ~pi0198;
  assign n5819 = n5453 & pi0634;
  assign n5820 = n5426 & pi0633;
  assign n5821 = ~n5819 & ~n5820;
  assign n5822 = n5397 & n5821;
  assign po0355 = ~n5818 & ~n5822;
  assign n5824 = ~n5397 & pi0199;
  assign n5825 = n5453 & pi0637;
  assign n5826 = n5426 & pi0617;
  assign n5827 = ~n5825 & ~n5826;
  assign n5828 = n5397 & ~n5827;
  assign po0356 = n5824 | n5828;
  assign n5830 = ~n5397 & ~pi0200;
  assign n5831 = n5453 & pi0643;
  assign n5832 = n5426 & pi0606;
  assign n5833 = ~n5831 & ~n5832;
  assign n5834 = n5397 & n5833;
  assign po0357 = ~n5830 & ~n5834;
  assign n5836 = n4439 & ~n2537;
  assign n5837 = ~n2776 & ~pi0332;
  assign n5838 = ~n5836 & n5837;
  assign n5839 = n2885 & pi0198;
  assign n5840 = ~n2885 & pi0210;
  assign n5841 = ~n5839 & ~n5840;
  assign n5842 = ~n5841 & pi0096;
  assign n5843 = ~pi0032 & pi0070;
  assign n5844 = ~n5842 & n5843;
  assign n5845 = n4097 & ~pi0070;
  assign n5846 = n5841 & n5845;
  assign n5847 = ~n5844 & ~n5846;
  assign n5848 = ~n5847 & pi0233;
  assign n5849 = n5848 & pi0237;
  assign n5850 = n5838 & ~n5849;
  assign n5851 = n2885 & n3398;
  assign n5852 = n3583 & ~n5851;
  assign n5853 = ~n3581 & ~pi0587;
  assign n5854 = n5853 & n2885;
  assign n5855 = ~n5852 & ~n5854;
  assign n5856 = ~n5855 & ~pi0332;
  assign n5857 = ~n5850 & ~n5856;
  assign n5858 = ~n5857 & ~pi0201;
  assign n5859 = n5842 & pi0237;
  assign n5860 = n5855 & pi0233;
  assign n5861 = n5859 & n5860;
  assign po0358 = n5858 | n5861;
  assign n5863 = ~n5847 & ~pi0233;
  assign n5864 = n5863 & pi0237;
  assign n5865 = n5838 & ~n5864;
  assign n5866 = ~n5865 & ~n5856;
  assign n5867 = ~n5866 & ~pi0202;
  assign n5868 = n5855 & ~pi0233;
  assign n5869 = n5859 & n5868;
  assign po0359 = n5867 | n5869;
  assign n5871 = n5863 & ~pi0237;
  assign n5872 = n5838 & ~n5871;
  assign n5873 = ~n5872 & ~n5856;
  assign n5874 = ~n5873 & ~pi0203;
  assign n5875 = n5842 & ~pi0237;
  assign n5876 = n5868 & n5875;
  assign po0360 = n5874 | n5876;
  assign n5878 = n2885 & ~pi0602;
  assign n5879 = ~n5878 & n3398;
  assign n5880 = ~n2885 & ~pi0907;
  assign n5881 = n5879 & ~n5880;
  assign n5882 = ~n5881 & ~n3575;
  assign n5883 = n5882 & ~pi0332;
  assign n5884 = ~n5850 & ~n5883;
  assign n5885 = ~n5884 & ~pi0204;
  assign n5886 = n5859 & ~n5882;
  assign n5887 = n5886 & pi0233;
  assign po0361 = n5885 | n5887;
  assign n5889 = ~n5865 & ~n5883;
  assign n5890 = ~n5889 & ~pi0205;
  assign n5891 = n5886 & ~pi0233;
  assign po0362 = n5890 | n5891;
  assign n5893 = n5848 & ~pi0237;
  assign n5894 = n5838 & ~n5893;
  assign n5895 = ~n5894 & ~n5883;
  assign n5896 = ~n5895 & ~pi0206;
  assign n5897 = n5875 & ~n5882;
  assign n5898 = n5897 & pi0233;
  assign po0363 = n5896 | n5898;
  assign n5900 = ~n5397 & pi0207;
  assign n5901 = n5453 & pi0710;
  assign n5902 = n5426 & pi0623;
  assign n5903 = ~n5901 & ~n5902;
  assign n5904 = n5397 & n5903;
  assign po0364 = ~n5900 & ~n5904;
  assign n5906 = ~n5397 & pi0208;
  assign n5907 = n5453 & pi0638;
  assign n5908 = n5426 & pi0607;
  assign n5909 = ~n5907 & ~n5908;
  assign n5910 = n5397 & n5909;
  assign po0365 = ~n5906 & ~n5910;
  assign n5912 = ~n5397 & pi0209;
  assign n5913 = n5453 & pi0639;
  assign n5914 = n5426 & pi0622;
  assign n5915 = ~n5913 & ~n5914;
  assign n5916 = n5397 & n5915;
  assign po0366 = ~n5912 & ~n5916;
  assign n5918 = ~n5397 & ~pi0210;
  assign n5919 = n5489 & pi0634;
  assign n5920 = pi0633 & pi0947;
  assign n5921 = ~n5919 & ~n5920;
  assign n5922 = n5397 & n5921;
  assign po0367 = ~n5918 & ~n5922;
  assign n5924 = ~n5397 & ~pi0211;
  assign n5925 = n5489 & pi0643;
  assign n5926 = pi0606 & pi0947;
  assign n5927 = ~n5925 & ~n5926;
  assign n5928 = n5397 & n5927;
  assign po0368 = ~n5924 & ~n5928;
  assign n5930 = ~n5397 & ~pi0212;
  assign n5931 = n5489 & pi0638;
  assign n5932 = pi0607 & pi0947;
  assign n5933 = ~n5931 & ~n5932;
  assign n5934 = n5515 & ~n5933;
  assign po0369 = n5930 | n5934;
  assign n5936 = ~n5397 & ~pi0213;
  assign n5937 = n5489 & pi0639;
  assign n5938 = pi0622 & pi0947;
  assign n5939 = ~n5937 & ~n5938;
  assign n5940 = n5515 & ~n5939;
  assign po0370 = n5936 | n5940;
  assign n5942 = ~n5397 & pi0214;
  assign n5943 = n5489 & pi0710;
  assign n5944 = pi0623 & pi0947;
  assign n5945 = ~n5943 & ~n5944;
  assign n5946 = n5397 & n5945;
  assign po0371 = ~n5942 & ~n5946;
  assign n5948 = ~n5397 & ~pi0215;
  assign n5949 = n5489 & pi0681;
  assign n5950 = pi0642 & pi0947;
  assign n5951 = ~n5949 & ~n5950;
  assign n5952 = n5397 & n5951;
  assign po0372 = ~n5948 & ~n5952;
  assign n5954 = ~n5397 & ~pi0216;
  assign n5955 = n5489 & pi0662;
  assign n5956 = pi0614 & pi0947;
  assign n5957 = ~n5955 & ~n5956;
  assign n5958 = n5397 & n5957;
  assign po0373 = ~n5954 & ~n5958;
  assign n5960 = ~n5397 & pi0217;
  assign n5961 = n5453 & ~pi0695;
  assign n5962 = n5426 & pi0612;
  assign n5963 = ~n5961 & ~n5962;
  assign n5964 = n5397 & n5963;
  assign po0374 = ~n5960 & ~n5964;
  assign n5966 = ~n5872 & ~n5883;
  assign n5967 = ~n5966 & ~pi0218;
  assign n5968 = n5897 & ~pi0233;
  assign po0375 = n5967 | n5968;
  assign n5970 = ~n5397 & pi0219;
  assign n5971 = n5489 & pi0637;
  assign n5972 = pi0617 & pi0947;
  assign n5973 = ~n5971 & ~n5972;
  assign n5974 = n5515 & ~n5973;
  assign po0376 = n5970 | n5974;
  assign n5976 = ~n5894 & ~n5856;
  assign n5977 = ~n5976 & ~pi0220;
  assign n5978 = n5860 & n5875;
  assign po0377 = n5977 | n5978;
  assign n5980 = ~n5397 & ~pi0221;
  assign n5981 = n5489 & pi0661;
  assign n5982 = pi0616 & pi0947;
  assign n5983 = ~n5981 & ~n5982;
  assign n5984 = n5397 & n5983;
  assign po0378 = ~n5980 & ~n5984;
  assign n5986 = ~n5397 & ~pi0222;
  assign n5987 = n5453 & pi0661;
  assign n5988 = n5426 & pi0616;
  assign n5989 = ~n5987 & ~n5988;
  assign n5990 = n5397 & n5989;
  assign po0379 = ~n5986 & ~n5990;
  assign n5992 = ~n5397 & ~pi0223;
  assign n5993 = n5453 & pi0681;
  assign n5994 = n5426 & pi0642;
  assign n5995 = ~n5993 & ~n5994;
  assign n5996 = n5397 & n5995;
  assign po0380 = ~n5992 & ~n5996;
  assign n5998 = ~n5397 & ~pi0224;
  assign n5999 = n5453 & pi0662;
  assign n6000 = n5426 & pi0614;
  assign n6001 = ~n5999 & ~n6000;
  assign n6002 = n5397 & n6001;
  assign po0381 = ~n5998 & ~n6002;
  assign n6004 = n2693 & n2748;
  assign n6005 = pi0070 & pi0332;
  assign n6006 = ~n2703 & ~n6005;
  assign n6007 = n2891 & ~n6006;
  assign n6008 = n4987 & n2669;
  assign n6009 = ~pi0055 & ~pi0137;
  assign n6010 = ~n6008 & n6009;
  assign n6011 = ~n2804 & ~n6010;
  assign n6012 = ~n6007 & ~n6011;
  assign po0382 = n6004 | ~n6012;
  assign n6014 = n2891 & n3386;
  assign n6015 = n2787 & ~n2799;
  assign n6016 = n4814 & pi0479;
  assign n6017 = n2803 & ~n6016;
  assign n6018 = ~n6015 & n6017;
  assign po0393 = n6014 | ~n6018;
  assign n6020 = po0393 & ~pi0228;
  assign n6021 = pi0228 & pi0231;
  assign po0383 = n6020 | n6021;
  assign n6023 = n4275 & pi1093;
  assign n6024 = n2676 & ~pi0058;
  assign n6025 = n6024 & n2577;
  assign n6026 = ~n6025 & ~pi0072;
  assign n6027 = ~n4429 & n6026;
  assign n6028 = ~n6023 & n6027;
  assign n6029 = n2891 & ~n6028;
  assign n6030 = ~n6029 & ~n4590;
  assign n6031 = po0840 & pi0036;
  assign po0384 = n6030 | n6031;
  assign n6033 = ~n3450 & ~n2640;
  assign n6034 = ~po1038 & n2863;
  assign n6035 = ~n6033 & n6034;
  assign n6036 = ~n2639 & n6035;
  assign n6037 = ~n6036 & ~pi0228;
  assign n6038 = ~n6037 & ~pi0039;
  assign n6039 = n4806 & pi1091;
  assign po0385 = n6038 | n6039;
  assign n6041 = po0740 & ~pi0047;
  assign n6042 = n2545 & n6041;
  assign n6043 = n6042 & ~n4039;
  assign po0387 = ~n5396 & ~n6043;
  assign po1049 = ~n4014 | pi0064;
  assign n6046 = ~pi0065 ^ ~pi0102;
  assign n6047 = ~po1049 & n6046;
  assign n6048 = n6047 & n2525;
  assign n6049 = ~n6048 & ~n4236;
  assign n6050 = ~n3479 & n6049;
  assign n6051 = ~n2804 & ~po0223;
  assign po0389 = n6050 | n6051;
  assign n6053 = n4471 & pi1155;
  assign n6054 = n4379 & pi1156;
  assign n6055 = ~n6053 & ~n6054;
  assign n6056 = pi0199 & ~pi0200;
  assign n6057 = n6056 & pi1154;
  assign n6058 = n6055 & ~n6057;
  assign n6059 = ~pi0207 & pi0208;
  assign n6060 = ~n6058 & n6059;
  assign n6061 = n6056 & pi1155;
  assign n6062 = n4471 & pi1156;
  assign n6063 = ~n6061 & ~n6062;
  assign n6064 = n4379 & pi1157;
  assign n6065 = n6063 & ~n6064;
  assign n6066 = pi0207 & ~pi0208;
  assign n6067 = ~n6065 & n6066;
  assign n6068 = ~n6060 & ~n6067;
  assign n6069 = n2885 & ~pi0209;
  assign n6070 = n6068 & n6069;
  assign n6071 = n4471 & pi1154;
  assign n6072 = n6056 & pi1153;
  assign n6073 = ~n6071 & ~n6072;
  assign n6074 = n4379 & pi1155;
  assign n6075 = n6073 & ~n6074;
  assign n6076 = ~n6075 & n4382;
  assign n6077 = n6070 & ~n6076;
  assign n6078 = pi0200 & pi1143;
  assign n6079 = ~pi0200 & pi1144;
  assign n6080 = ~n6078 & ~n6079;
  assign n6081 = pi0207 ^ ~pi0208;
  assign n6082 = ~n6080 & ~n6081;
  assign n6083 = n4382 & ~pi0200;
  assign n6084 = n6083 & pi1143;
  assign n6085 = ~n6082 & ~n6084;
  assign n6086 = ~n4379 & pi1142;
  assign n6087 = ~n4383 & n6086;
  assign n6088 = n6085 & ~n6087;
  assign n6089 = ~pi0207 & ~pi0208;
  assign n6090 = ~n6089 & ~pi0200;
  assign n6091 = n6090 & pi1142;
  assign n6092 = ~n6091 & pi0199;
  assign n6093 = ~n6088 & ~n6092;
  assign n6094 = n2885 & pi0209;
  assign n6095 = ~n6093 & n6094;
  assign n6096 = ~n6095 & pi0230;
  assign n6097 = ~n6077 & n6096;
  assign n6098 = ~pi0219 & pi1156;
  assign n6099 = pi0219 & pi1154;
  assign n6100 = ~n6098 & ~n6099;
  assign n6101 = n6100 & ~pi0214;
  assign n6102 = ~n6101 & ~pi0211;
  assign n6103 = pi0219 & pi1153;
  assign n6104 = ~pi0219 & pi1155;
  assign n6105 = ~n6103 & ~n6104;
  assign n6106 = n6105 & pi0214;
  assign n6107 = n6102 & ~n6106;
  assign n6108 = ~pi0214 & ~pi1155;
  assign n6109 = n4468 & ~n6108;
  assign n6110 = pi0214 & ~pi1154;
  assign n6111 = n6109 & ~n6110;
  assign n6112 = ~n6107 & ~n6111;
  assign n6113 = ~n6112 & pi0212;
  assign n6114 = ~n2885 & ~pi0213;
  assign n6115 = pi0219 & pi1155;
  assign n6116 = ~pi0219 & pi1157;
  assign n6117 = ~n6115 & ~n6116;
  assign n6118 = n6117 & ~pi0211;
  assign n6119 = ~n6098 & pi0211;
  assign n6120 = ~pi0212 & pi0214;
  assign n6121 = ~n6119 & n6120;
  assign n6122 = ~n6118 & n6121;
  assign n6123 = n6114 & ~n6122;
  assign n6124 = ~n6113 & n6123;
  assign n6125 = ~pi0212 & ~pi0214;
  assign n6126 = n4467 & ~n6125;
  assign n6127 = n6126 & pi1143;
  assign n6128 = n4385 & n4468;
  assign n6129 = n4465 & ~n6125;
  assign n6130 = ~n6128 & ~n6129;
  assign n6131 = ~n6130 & pi1142;
  assign n6132 = pi0212 ^ ~pi0214;
  assign n6133 = n4400 & ~n6132;
  assign n6134 = n6133 & pi1144;
  assign n6135 = ~n6131 & ~n6134;
  assign n6136 = ~n6127 & n6135;
  assign n6137 = ~n2885 & pi0213;
  assign n6138 = n6136 & n6137;
  assign n6139 = ~n6124 & ~n6138;
  assign n6140 = n6097 & n6139;
  assign n6141 = ~pi0230 & ~pi0233;
  assign po0390 = n6140 | n6141;
  assign n6143 = n2885 & n6089;
  assign n6144 = ~n2885 & n6125;
  assign n6145 = ~n6143 & ~n6144;
  assign n6146 = n4476 & n6145;
  assign n6147 = n6146 & ~n4390;
  assign n6148 = n6147 & pi1152;
  assign n6149 = n4476 & ~pi1153;
  assign n6150 = n4390 & n6145;
  assign n6151 = ~n6149 & n6150;
  assign n6152 = ~n4476 & ~pi1154;
  assign n6153 = n6151 & ~n6152;
  assign n6154 = ~n6148 & ~n6153;
  assign n6155 = ~n6094 & ~n6137;
  assign n6156 = n6154 & n6155;
  assign n6157 = n6147 & pi1154;
  assign n6158 = n6126 & pi1155;
  assign n6159 = n6133 & pi1156;
  assign n6160 = n6137 & ~n6159;
  assign n6161 = ~n6158 & n6160;
  assign n6162 = ~n6055 & ~n6081;
  assign n6163 = n6074 & n4382;
  assign n6164 = ~n6162 & ~n6163;
  assign n6165 = n6094 & n6164;
  assign n6166 = ~n6161 & ~n6165;
  assign n6167 = ~n6157 & ~n6166;
  assign n6168 = ~n6167 & pi0230;
  assign n6169 = ~n6156 & n6168;
  assign n6170 = ~pi0230 & pi0234;
  assign po0391 = n6169 | n6170;
  assign n6172 = ~n6075 & ~pi0209;
  assign n6173 = ~n6065 & pi0209;
  assign n6174 = ~n6172 & ~n6173;
  assign n6175 = ~n6174 & ~n6081;
  assign n6176 = n4471 & pi1153;
  assign n6177 = n4379 & pi1154;
  assign n6178 = ~n6176 & ~n6177;
  assign n6179 = n6069 & n6178;
  assign n6180 = n6055 & pi0209;
  assign n6181 = ~n6180 & n4382;
  assign n6182 = ~n6181 & n2885;
  assign n6183 = ~n6179 & ~n6182;
  assign n6184 = ~n6175 & ~n6183;
  assign n6185 = ~pi0213 & pi1154;
  assign n6186 = pi0213 & pi1156;
  assign n6187 = ~n6185 & ~n6186;
  assign n6188 = n6126 & ~n6187;
  assign n6189 = n6105 & ~pi0213;
  assign n6190 = ~n6132 & ~pi0211;
  assign n6191 = ~n6189 & n6190;
  assign n6192 = n6117 & pi0213;
  assign n6193 = n6191 & ~n6192;
  assign n6194 = ~pi0213 & pi1153;
  assign n6195 = pi0213 & pi1155;
  assign n6196 = ~n6194 & ~n6195;
  assign n6197 = n6128 & ~n6196;
  assign n6198 = ~n2885 & ~n6197;
  assign n6199 = ~n6193 & n6198;
  assign n6200 = ~n6188 & n6199;
  assign n6201 = ~n6200 & pi0230;
  assign n6202 = ~n6184 & n6201;
  assign n6203 = ~pi0230 & pi0235;
  assign po0392 = n6202 | n6203;
  assign n6205 = n6117 & ~pi0214;
  assign n6206 = n6100 & pi0214;
  assign n6207 = ~n6205 & ~n6206;
  assign n6208 = n6207 & ~pi0211;
  assign n6209 = pi0214 & ~pi1155;
  assign n6210 = n4468 & ~n6209;
  assign n6211 = ~pi0214 & ~pi1156;
  assign n6212 = n6210 & ~n6211;
  assign n6213 = ~n6208 & ~n6212;
  assign n6214 = ~n6213 & pi0212;
  assign n6215 = n4465 & pi1156;
  assign n6216 = n4468 & pi1157;
  assign n6217 = ~n6215 & ~n6216;
  assign n6218 = n4400 & pi1158;
  assign n6219 = n6217 & ~n6218;
  assign n6220 = ~n6219 & n6120;
  assign n6221 = ~n6214 & ~n6220;
  assign n6222 = ~n6221 & n6114;
  assign n6223 = ~n6065 & n6059;
  assign n6224 = n4471 & pi1157;
  assign n6225 = n6056 & pi1156;
  assign n6226 = ~n6224 & ~n6225;
  assign n6227 = n4379 & pi1158;
  assign n6228 = n6226 & ~n6227;
  assign n6229 = ~n6228 & n6066;
  assign n6230 = ~n6223 & ~n6229;
  assign n6231 = ~n6058 & n4382;
  assign n6232 = n6230 & ~n6231;
  assign n6233 = ~n6232 & n6069;
  assign n6234 = ~n6130 & pi1143;
  assign n6235 = ~n6132 & ~pi0219;
  assign n6236 = ~pi0211 & pi1145;
  assign n6237 = pi0211 & pi1144;
  assign n6238 = ~n6236 & ~n6237;
  assign n6239 = n6235 & ~n6238;
  assign n6240 = n4401 & pi1144;
  assign n6241 = ~n6239 & ~n6240;
  assign n6242 = ~n6234 & n6241;
  assign n6243 = n6137 & ~n6242;
  assign n6244 = ~n6243 & pi0230;
  assign n6245 = ~n6233 & n6244;
  assign n6246 = ~n6222 & n6245;
  assign n6247 = ~n6081 & pi0200;
  assign n6248 = ~n6083 & ~n6247;
  assign n6249 = ~n6248 & pi1144;
  assign n6250 = n4382 & n6078;
  assign n6251 = ~n6249 & ~n6250;
  assign n6252 = ~n6251 & ~pi0199;
  assign n6253 = n4383 & pi1145;
  assign n6254 = pi0199 & pi1143;
  assign n6255 = ~n6253 & ~n6254;
  assign n6256 = ~n6255 & n6090;
  assign n6257 = ~n6252 & ~n6256;
  assign n6258 = ~n6257 & n6094;
  assign n6259 = n6246 & ~n6258;
  assign n6260 = ~pi0230 & pi0237;
  assign po0394 = ~n6259 & ~n6260;
  assign n6262 = n6147 & pi1151;
  assign n6263 = n4476 & ~pi1152;
  assign n6264 = n6150 & ~n6263;
  assign n6265 = ~n4476 & ~pi1153;
  assign n6266 = n6264 & ~n6265;
  assign n6267 = ~n6262 & ~n6266;
  assign n6268 = n6267 & n6155;
  assign n6269 = ~n6072 & n4382;
  assign n6270 = ~n6269 & ~n6089;
  assign n6271 = ~n6075 & n6270;
  assign n6272 = n6094 & ~n6271;
  assign n6273 = ~n6178 & n4382;
  assign n6274 = n6272 & ~n6273;
  assign n6275 = ~n6130 & pi1153;
  assign n6276 = n4401 & pi1154;
  assign n6277 = ~pi0211 & pi1155;
  assign n6278 = pi0211 & pi1154;
  assign n6279 = ~n6277 & ~n6278;
  assign n6280 = n6235 & ~n6279;
  assign n6281 = ~n6276 & ~n6280;
  assign n6282 = ~n6275 & n6281;
  assign n6283 = n6137 & n6282;
  assign n6284 = ~n6283 & pi0230;
  assign n6285 = ~n6274 & n6284;
  assign n6286 = ~n6268 & n6285;
  assign n6287 = ~pi0230 & pi0238;
  assign po0395 = n6286 | n6287;
  assign n6289 = n6213 & ~pi0213;
  assign n6290 = n6219 & pi0213;
  assign n6291 = ~n2885 & n6120;
  assign n6292 = ~n6290 & n6291;
  assign n6293 = ~n6289 & n6292;
  assign n6294 = n6228 & pi0209;
  assign n6295 = n6058 & ~pi0209;
  assign n6296 = ~n6294 & ~n6295;
  assign n6297 = n2885 & n6066;
  assign n6298 = n6296 & n6297;
  assign n6299 = ~n6298 & pi0230;
  assign n6300 = ~n6293 & n6299;
  assign n6301 = ~pi0230 & ~pi0239;
  assign po0396 = ~n6300 & ~n6301;
  assign n6303 = n6147 & pi1145;
  assign n6304 = ~n4476 & ~pi1147;
  assign n6305 = n6150 & ~n6304;
  assign n6306 = n4476 & ~pi1146;
  assign n6307 = n6305 & ~n6306;
  assign n6308 = ~n6303 & ~n6307;
  assign n6309 = ~n6308 & n6155;
  assign n6310 = n6147 & pi1147;
  assign n6311 = ~n4476 & ~pi1149;
  assign n6312 = n6150 & ~n6311;
  assign n6313 = n4476 & ~pi1148;
  assign n6314 = n6312 & ~n6313;
  assign n6315 = ~n6310 & ~n6314;
  assign n6316 = ~n6315 & ~n6155;
  assign n6317 = ~n6309 & ~n6316;
  assign n6318 = n6317 & pi0230;
  assign n6319 = ~pi0230 & ~pi0240;
  assign po0397 = ~n6318 & ~n6319;
  assign n6321 = n6147 & pi1149;
  assign n6322 = ~n4476 & ~pi1151;
  assign n6323 = n6150 & ~n6322;
  assign n6324 = n4476 & ~pi1150;
  assign n6325 = n6323 & ~n6324;
  assign n6326 = ~n6321 & ~n6325;
  assign n6327 = ~n6326 & n6155;
  assign n6328 = ~n6267 & ~n6155;
  assign n6329 = ~n6327 & ~n6328;
  assign n6330 = n6329 & pi0230;
  assign n6331 = ~pi0230 & ~pi0241;
  assign po0398 = ~n6330 & ~n6331;
  assign n6333 = n6147 & pi1144;
  assign n6334 = n4476 & ~pi1145;
  assign n6335 = n6150 & ~n6334;
  assign n6336 = ~n4476 & ~pi1146;
  assign n6337 = n6335 & ~n6336;
  assign n6338 = ~n6333 & ~n6337;
  assign n6339 = n6338 & ~n6155;
  assign n6340 = n6136 & n6114;
  assign n6341 = ~n6093 & n6069;
  assign n6342 = ~n6341 & pi0230;
  assign n6343 = ~n6340 & n6342;
  assign n6344 = ~n6339 & n6343;
  assign n6345 = ~pi0230 & pi0242;
  assign po0399 = n6344 | n6345;
  assign n6347 = ~po1038 & n4541;
  assign n6348 = ~n6347 & pi0081;
  assign n6349 = ~n4389 & n6348;
  assign n6350 = ~pi0083 & ~pi0085;
  assign n6351 = ~n6349 & n6350;
  assign n6352 = ~n6351 & pi0314;
  assign n6353 = n6352 & pi0802;
  assign n6354 = n6353 & pi0276;
  assign n6355 = n6354 & pi0271;
  assign n6356 = n6355 & pi0273;
  assign n6357 = n6356 & pi0283;
  assign n6358 = n6357 & pi0272;
  assign n6359 = n6358 & pi0275;
  assign n6360 = n6359 & pi0268;
  assign n6361 = n6360 & pi0253;
  assign n6362 = n6361 & pi0254;
  assign n6363 = n6362 & pi0267;
  assign n6364 = n6363 & ~pi0263;
  assign n6365 = ~n6364 ^ ~pi0243;
  assign n6366 = ~pi0230 & ~pi1091;
  assign n6367 = ~n6365 & n6366;
  assign n6368 = n2885 & ~n6056;
  assign n6369 = ~n4466 & ~n6368;
  assign n6370 = n6369 & pi1157;
  assign n6371 = ~n2885 & ~n4400;
  assign n6372 = ~n6371 & ~n4381;
  assign n6373 = n6372 & pi1155;
  assign n6374 = ~n6370 & ~n6373;
  assign n6375 = ~n2885 & ~n4468;
  assign n6376 = ~n6375 & ~n4473;
  assign n6377 = n6376 & pi1156;
  assign n6378 = n6374 & ~n6377;
  assign n6379 = ~n6378 & ~n6366;
  assign po0400 = n6367 | n6379;
  assign n6381 = n6308 & ~n6155;
  assign n6382 = n6257 & n6069;
  assign n6383 = n6114 & n6242;
  assign n6384 = ~n6383 & pi0230;
  assign n6385 = ~n6382 & n6384;
  assign n6386 = ~n6381 & n6385;
  assign n6387 = ~pi0230 & pi0244;
  assign po0401 = n6386 | n6387;
  assign n6389 = ~n6338 & n6155;
  assign n6390 = n6147 & pi1146;
  assign n6391 = ~n4476 & ~pi1148;
  assign n6392 = n6150 & ~n6391;
  assign n6393 = n4476 & ~pi1147;
  assign n6394 = n6392 & ~n6393;
  assign n6395 = ~n6390 & ~n6394;
  assign n6396 = ~n6395 & ~n6155;
  assign n6397 = ~n6389 & ~n6396;
  assign n6398 = n6397 & pi0230;
  assign n6399 = ~pi0230 & ~pi0245;
  assign po0402 = ~n6398 & ~n6399;
  assign n6401 = ~n6395 & n6155;
  assign n6402 = n6147 & pi1148;
  assign n6403 = ~n4476 & ~pi1150;
  assign n6404 = n6150 & ~n6403;
  assign n6405 = n4476 & ~pi1149;
  assign n6406 = n6404 & ~n6405;
  assign n6407 = ~n6402 & ~n6406;
  assign n6408 = ~n6407 & ~n6155;
  assign n6409 = ~n6401 & ~n6408;
  assign n6410 = n6409 & pi0230;
  assign n6411 = ~pi0230 & ~pi0246;
  assign po0403 = ~n6410 & ~n6411;
  assign n6413 = ~n6315 & n6155;
  assign n6414 = ~n6326 & ~n6155;
  assign n6415 = ~n6413 & ~n6414;
  assign n6416 = n6415 & pi0230;
  assign n6417 = ~pi0230 & ~pi0247;
  assign po0404 = ~n6416 & ~n6417;
  assign n6419 = ~n6407 & n6155;
  assign n6420 = n6147 & pi1150;
  assign n6421 = ~n4476 & ~pi1152;
  assign n6422 = n6150 & ~n6421;
  assign n6423 = n4476 & ~pi1151;
  assign n6424 = n6422 & ~n6423;
  assign n6425 = ~n6420 & ~n6424;
  assign n6426 = ~n6425 & ~n6155;
  assign n6427 = ~n6419 & ~n6426;
  assign n6428 = n6427 & pi0230;
  assign n6429 = ~pi0230 & ~pi0248;
  assign po0405 = ~n6428 & ~n6429;
  assign n6431 = ~n6425 & n6155;
  assign n6432 = ~n6154 & ~n6155;
  assign n6433 = ~n6431 & ~n6432;
  assign n6434 = n6433 & pi0230;
  assign n6435 = ~pi0230 & ~pi0249;
  assign po0406 = ~n6434 & ~n6435;
  assign n6437 = ~n4987 & ~n4450;
  assign po0407 = ~n6437 & ~pi0250;
  assign n6439 = n4379 & pi0897;
  assign n6440 = n4471 & ~pi0476;
  assign n6441 = ~n6439 & ~n6440;
  assign n6442 = n6441 & pi0251;
  assign n6443 = pi0200 & pi1039;
  assign n6444 = ~pi0200 & pi1053;
  assign n6445 = ~n6443 & ~n6444;
  assign n6446 = ~n6441 & ~n6445;
  assign po0408 = n6442 | n6446;
  assign n6448 = n3420 & ~n3431;
  assign n6449 = n3631 & n6448;
  assign n6450 = ~n3927 & pi1093;
  assign n6451 = pi0252 & pi1092;
  assign n6452 = ~n6450 & n6451;
  assign po0409 = n6449 | n6452;
  assign n6454 = ~n6360 ^ ~pi0253;
  assign n6455 = n6454 & n6366;
  assign n6456 = n6369 & pi1153;
  assign n6457 = n6372 & pi1151;
  assign n6458 = ~n6456 & ~n6457;
  assign n6459 = n6376 & pi1152;
  assign n6460 = n6458 & ~n6459;
  assign n6461 = ~n6460 & ~n6366;
  assign po0410 = n6455 | n6461;
  assign n6463 = ~n6361 ^ ~pi0254;
  assign n6464 = n6463 & n6366;
  assign n6465 = n6376 & pi1153;
  assign n6466 = n6372 & pi1152;
  assign n6467 = ~n6465 & ~n6466;
  assign n6468 = n6369 & pi1154;
  assign n6469 = n6467 & ~n6468;
  assign n6470 = ~n6469 & ~n6366;
  assign po0411 = n6464 | n6470;
  assign n6472 = n6441 & pi0255;
  assign n6473 = pi0200 & pi1036;
  assign n6474 = ~pi0200 & pi1049;
  assign n6475 = ~n6473 & ~n6474;
  assign n6476 = ~n6441 & ~n6475;
  assign po0412 = n6472 | n6476;
  assign n6478 = n6441 & pi0256;
  assign n6479 = pi0200 & pi1070;
  assign n6480 = ~pi0200 & pi1048;
  assign n6481 = ~n6479 & ~n6480;
  assign n6482 = ~n6441 & ~n6481;
  assign po0413 = n6478 | n6482;
  assign n6484 = n6441 & pi0257;
  assign n6485 = pi0200 & pi1065;
  assign n6486 = ~pi0200 & pi1084;
  assign n6487 = ~n6485 & ~n6486;
  assign n6488 = ~n6441 & ~n6487;
  assign po0414 = n6484 | n6488;
  assign n6490 = n6441 & pi0258;
  assign n6491 = pi0200 & pi1062;
  assign n6492 = ~pi0200 & pi1072;
  assign n6493 = ~n6491 & ~n6492;
  assign n6494 = ~n6441 & ~n6493;
  assign po0415 = n6490 | n6494;
  assign n6496 = n6441 & pi0259;
  assign n6497 = pi0200 & pi1069;
  assign n6498 = ~pi0200 & pi1059;
  assign n6499 = ~n6497 & ~n6498;
  assign n6500 = ~n6441 & ~n6499;
  assign po0416 = n6496 | n6500;
  assign n6502 = n6441 & pi0260;
  assign n6503 = pi0200 & pi1067;
  assign n6504 = ~pi0200 & pi1044;
  assign n6505 = ~n6503 & ~n6504;
  assign n6506 = ~n6441 & ~n6505;
  assign po0417 = n6502 | n6506;
  assign n6508 = n6441 & pi0261;
  assign n6509 = pi0200 & pi1040;
  assign n6510 = ~pi0200 & pi1037;
  assign n6511 = ~n6509 & ~n6510;
  assign n6512 = ~n6441 & ~n6511;
  assign po0418 = n6508 | n6512;
  assign n6514 = ~pi0228 & pi1093;
  assign n6515 = ~pi0123 & pi0228;
  assign n6516 = ~n6514 & ~n6515;
  assign n6517 = n6150 & ~n6516;
  assign n6518 = n6517 & pi1142;
  assign n6519 = n6516 & ~pi0262;
  assign po0419 = n6518 | n6519;
  assign n6521 = n6363 ^ ~pi0263;
  assign n6522 = n6521 & n6366;
  assign n6523 = n6369 & pi1156;
  assign n6524 = n6372 & pi1154;
  assign n6525 = ~n6523 & ~n6524;
  assign n6526 = n6376 & pi1155;
  assign n6527 = n6525 & ~n6526;
  assign n6528 = ~n6527 & ~n6366;
  assign po0420 = n6522 | n6528;
  assign n6530 = ~n6352 & pi0264;
  assign n6531 = n6352 & ~pi0796;
  assign n6532 = ~n6530 & ~n6531;
  assign n6533 = n6532 & n6366;
  assign n6534 = n6372 & pi1141;
  assign n6535 = n6369 & pi1143;
  assign n6536 = ~n6534 & ~n6535;
  assign n6537 = n6376 & pi1142;
  assign n6538 = n6536 & ~n6537;
  assign n6539 = ~n6538 & ~n6366;
  assign po0421 = n6533 | n6539;
  assign n6541 = ~n6352 & pi0265;
  assign n6542 = n6352 & ~pi0819;
  assign n6543 = ~n6541 & ~n6542;
  assign n6544 = n6543 & n6366;
  assign n6545 = n6372 & pi1142;
  assign n6546 = n6369 & pi1144;
  assign n6547 = ~n6545 & ~n6546;
  assign n6548 = n6376 & pi1143;
  assign n6549 = n6547 & ~n6548;
  assign n6550 = ~n6549 & ~n6366;
  assign po0422 = n6544 | n6550;
  assign n6552 = ~n6352 & ~pi0266;
  assign n6553 = n6352 & ~pi0948;
  assign n6554 = ~n6552 & ~n6553;
  assign n6555 = n6554 & n6366;
  assign n6556 = n6372 & pi1134;
  assign n6557 = n6369 & pi1136;
  assign n6558 = ~n6556 & ~n6557;
  assign n6559 = n6376 & pi1135;
  assign n6560 = n6558 & ~n6559;
  assign n6561 = ~n6560 & ~n6366;
  assign po0423 = n6555 | n6561;
  assign n6563 = ~n6362 ^ ~pi0267;
  assign n6564 = n6563 & n6366;
  assign n6565 = n6376 & pi1154;
  assign n6566 = n6372 & pi1153;
  assign n6567 = ~n6565 & ~n6566;
  assign n6568 = n6369 & pi1155;
  assign n6569 = n6567 & ~n6568;
  assign n6570 = ~n6569 & ~n6366;
  assign po0424 = n6564 | n6570;
  assign n6572 = ~n6359 ^ ~pi0268;
  assign n6573 = n6572 & n6366;
  assign n6574 = n6369 & pi1152;
  assign n6575 = n6372 & pi1150;
  assign n6576 = ~n6574 & ~n6575;
  assign n6577 = n6376 & pi1151;
  assign n6578 = n6576 & ~n6577;
  assign n6579 = ~n6578 & ~n6366;
  assign po0425 = n6573 | n6579;
  assign n6581 = ~n6352 & pi0269;
  assign n6582 = n6352 & ~pi0817;
  assign n6583 = ~n6581 & ~n6582;
  assign n6584 = n6583 & n6366;
  assign n6585 = n6372 & pi1136;
  assign n6586 = n6369 & pi1138;
  assign n6587 = ~n6585 & ~n6586;
  assign n6588 = n6376 & pi1137;
  assign n6589 = n6587 & ~n6588;
  assign n6590 = ~n6589 & ~n6366;
  assign po0426 = n6584 | n6590;
  assign n6592 = ~n6352 & pi0270;
  assign n6593 = n6352 & ~pi0805;
  assign n6594 = ~n6592 & ~n6593;
  assign n6595 = n6594 & n6366;
  assign n6596 = n6372 & pi1139;
  assign n6597 = n6369 & pi1141;
  assign n6598 = ~n6596 & ~n6597;
  assign n6599 = n6376 & pi1140;
  assign n6600 = n6598 & ~n6599;
  assign n6601 = ~n6600 & ~n6366;
  assign po0427 = n6595 | n6601;
  assign n6603 = ~n6354 ^ ~pi0271;
  assign n6604 = n6603 & n6366;
  assign n6605 = n6376 & pi1146;
  assign n6606 = n6372 & pi1145;
  assign n6607 = ~n6605 & ~n6606;
  assign n6608 = n6369 & pi1147;
  assign n6609 = n6607 & ~n6608;
  assign n6610 = ~n6609 & ~n6366;
  assign po0428 = n6604 | n6610;
  assign n6612 = ~n6357 ^ ~pi0272;
  assign n6613 = n6612 & n6366;
  assign n6614 = n6369 & pi1150;
  assign n6615 = n6372 & pi1148;
  assign n6616 = ~n6614 & ~n6615;
  assign n6617 = n6376 & pi1149;
  assign n6618 = n6616 & ~n6617;
  assign n6619 = ~n6618 & ~n6366;
  assign po0429 = n6613 | n6619;
  assign n6621 = ~n6355 ^ ~pi0273;
  assign n6622 = n6621 & n6366;
  assign n6623 = n6372 & pi1146;
  assign n6624 = n6369 & pi1148;
  assign n6625 = ~n6623 & ~n6624;
  assign n6626 = n6376 & pi1147;
  assign n6627 = n6625 & ~n6626;
  assign n6628 = ~n6627 & ~n6366;
  assign po0430 = n6622 | n6628;
  assign n6630 = ~n6352 & pi0274;
  assign n6631 = n6352 & ~pi0659;
  assign n6632 = ~n6630 & ~n6631;
  assign n6633 = n6632 & n6366;
  assign n6634 = n6369 & pi1145;
  assign n6635 = n6372 & pi1143;
  assign n6636 = ~n6634 & ~n6635;
  assign n6637 = n6376 & pi1144;
  assign n6638 = n6636 & ~n6637;
  assign n6639 = ~n6638 & ~n6366;
  assign po0431 = n6633 | n6639;
  assign n6641 = ~n6358 ^ ~pi0275;
  assign n6642 = n6641 & n6366;
  assign n6643 = n6369 & pi1151;
  assign n6644 = n6372 & pi1149;
  assign n6645 = ~n6643 & ~n6644;
  assign n6646 = n6376 & pi1150;
  assign n6647 = n6645 & ~n6646;
  assign n6648 = ~n6647 & ~n6366;
  assign po0432 = n6642 | n6648;
  assign n6650 = ~n6353 ^ ~pi0276;
  assign n6651 = n6650 & n6366;
  assign n6652 = n6369 & pi1146;
  assign n6653 = n6372 & pi1144;
  assign n6654 = ~n6652 & ~n6653;
  assign n6655 = n6376 & pi1145;
  assign n6656 = n6654 & ~n6655;
  assign n6657 = ~n6656 & ~n6366;
  assign po0433 = n6651 | n6657;
  assign n6659 = ~n6352 & pi0277;
  assign n6660 = n6352 & ~pi0820;
  assign n6661 = ~n6659 & ~n6660;
  assign n6662 = n6661 & n6366;
  assign n6663 = n6372 & pi1140;
  assign n6664 = n6369 & pi1142;
  assign n6665 = ~n6663 & ~n6664;
  assign n6666 = n6376 & pi1141;
  assign n6667 = n6665 & ~n6666;
  assign n6668 = ~n6667 & ~n6366;
  assign po0434 = n6662 | n6668;
  assign n6670 = ~n6352 & ~pi0278;
  assign n6671 = n6352 & ~pi0976;
  assign n6672 = ~n6670 & ~n6671;
  assign n6673 = n6672 & n6366;
  assign n6674 = n6372 & pi1132;
  assign n6675 = n6369 & pi1134;
  assign n6676 = ~n6674 & ~n6675;
  assign n6677 = n6376 & pi1133;
  assign n6678 = n6676 & ~n6677;
  assign n6679 = ~n6678 & ~n6366;
  assign po0435 = n6673 | n6679;
  assign n6681 = ~n6352 & ~pi0279;
  assign n6682 = n6352 & ~pi0958;
  assign n6683 = ~n6681 & ~n6682;
  assign n6684 = n6683 & n6366;
  assign n6685 = n6372 & pi1133;
  assign n6686 = n6369 & pi1135;
  assign n6687 = ~n6685 & ~n6686;
  assign n6688 = n6376 & pi1134;
  assign n6689 = n6687 & ~n6688;
  assign n6690 = ~n6689 & ~n6366;
  assign po0436 = n6684 | n6690;
  assign n6692 = ~n6352 & pi0280;
  assign n6693 = n6352 & ~pi0914;
  assign n6694 = ~n6692 & ~n6693;
  assign n6695 = n6694 & n6366;
  assign n6696 = n6372 & pi1135;
  assign n6697 = n6369 & pi1137;
  assign n6698 = ~n6696 & ~n6697;
  assign n6699 = n6376 & pi1136;
  assign n6700 = n6698 & ~n6699;
  assign n6701 = ~n6700 & ~n6366;
  assign po0437 = n6695 | n6701;
  assign n6703 = ~n6352 & pi0281;
  assign n6704 = n6352 & ~pi0830;
  assign n6705 = ~n6703 & ~n6704;
  assign n6706 = n6705 & n6366;
  assign n6707 = n6372 & pi1137;
  assign n6708 = n6369 & pi1139;
  assign n6709 = ~n6707 & ~n6708;
  assign n6710 = n6376 & pi1138;
  assign n6711 = n6709 & ~n6710;
  assign n6712 = ~n6711 & ~n6366;
  assign po0438 = n6706 | n6712;
  assign n6714 = ~n6352 & pi0282;
  assign n6715 = n6352 & ~pi0836;
  assign n6716 = ~n6714 & ~n6715;
  assign n6717 = n6716 & n6366;
  assign n6718 = n6372 & pi1138;
  assign n6719 = n6369 & pi1140;
  assign n6720 = ~n6718 & ~n6719;
  assign n6721 = n6376 & pi1139;
  assign n6722 = n6720 & ~n6721;
  assign n6723 = ~n6722 & ~n6366;
  assign po0439 = n6717 | n6723;
  assign n6725 = ~n6356 ^ ~pi0283;
  assign n6726 = n6725 & n6366;
  assign n6727 = n6369 & pi1149;
  assign n6728 = n6372 & pi1147;
  assign n6729 = ~n6727 & ~n6728;
  assign n6730 = n6376 & pi1148;
  assign n6731 = n6729 & ~n6730;
  assign n6732 = ~n6731 & ~n6366;
  assign po0440 = n6726 | n6732;
  assign n6734 = ~n4476 & pi1143;
  assign n6735 = n6517 & n6734;
  assign n6736 = n6516 & ~pi0284;
  assign po0441 = n6735 | n6736;
  assign po0637 = n4449 & ~n4340;
  assign n6739 = po0637 & ~n3949;
  assign n6740 = n6739 & pi0289;
  assign n6741 = pi0286 & pi0288;
  assign n6742 = n6740 & n6741;
  assign n6743 = ~n6742 ^ ~pi0285;
  assign n6744 = n3949 & ~pi0288;
  assign n6745 = ~po0637 & n6744;
  assign n6746 = n3918 & pi0285;
  assign n6747 = n6745 & n6746;
  assign n6748 = ~n6747 & ~pi0793;
  assign po0442 = n6743 & n6748;
  assign n6750 = n6739 & pi0288;
  assign n6751 = ~n6750 & ~n6745;
  assign n6752 = ~n6751 & pi0286;
  assign n6753 = ~n6752 & ~pi0793;
  assign n6754 = n6745 & ~n3920;
  assign n6755 = ~n6754 & ~n6750;
  assign n6756 = n6755 & ~pi0286;
  assign po0443 = n6753 & ~n6756;
  assign n6758 = ~pi0287 & pi0457;
  assign po0444 = ~n6758 & ~pi0332;
  assign n6760 = n3956 ^ ~pi0288;
  assign n6761 = po0637 ^ ~n6760;
  assign po0445 = n6761 & ~pi0793;
  assign n6763 = ~n6750 & ~pi0289;
  assign n6764 = ~n6740 & pi0286;
  assign n6765 = ~n6763 & n6764;
  assign n6766 = ~n6741 & pi0289;
  assign n6767 = ~n6745 & n6766;
  assign n6768 = ~n6747 & ~n6767;
  assign n6769 = ~n6765 & n6768;
  assign po0446 = ~n6769 & ~pi0793;
  assign n6771 = pi0290 & pi0476;
  assign n6772 = ~pi0476 & pi1048;
  assign po0447 = n6771 | n6772;
  assign n6774 = pi0291 & pi0476;
  assign n6775 = ~pi0476 & pi1049;
  assign po0448 = n6774 | n6775;
  assign n6777 = pi0292 & pi0476;
  assign n6778 = ~pi0476 & pi1084;
  assign po0449 = n6777 | n6778;
  assign n6780 = pi0293 & pi0476;
  assign n6781 = ~pi0476 & pi1059;
  assign po0450 = n6780 | n6781;
  assign n6783 = pi0294 & pi0476;
  assign n6784 = ~pi0476 & pi1072;
  assign po0451 = n6783 | n6784;
  assign n6786 = pi0295 & pi0476;
  assign n6787 = ~pi0476 & pi1053;
  assign po0452 = n6786 | n6787;
  assign n6789 = pi0296 & pi0476;
  assign n6790 = ~pi0476 & pi1037;
  assign po0453 = n6789 | n6790;
  assign n6792 = pi0297 & pi0476;
  assign n6793 = ~pi0476 & pi1044;
  assign po0454 = n6792 | n6793;
  assign n6795 = pi0298 & pi0478;
  assign n6796 = ~pi0478 & pi1044;
  assign po0455 = n6795 | n6796;
  assign n6798 = n4281 & pi0106;
  assign n6799 = pi0039 & ~pi0287;
  assign n6800 = n4480 & n6799;
  assign n6801 = ~n4485 & ~n6800;
  assign n6802 = ~n6798 & n6801;
  assign n6803 = n2776 & ~po1038;
  assign po0456 = ~n6802 | n6803;
  assign n6805 = n2754 & ~pi0024;
  assign n6806 = n6805 & ~pi0312;
  assign n6807 = n6806 ^ ~pi0300;
  assign po0457 = ~n6807 | pi0055;
  assign n6809 = ~pi0300 & ~pi0312;
  assign n6810 = n6805 & n6809;
  assign n6811 = n6810 ^ ~pi0301;
  assign po0458 = n6811 & ~pi0055;
  assign n6813 = n2885 & n2928;
  assign n6814 = ~n2885 & n2901;
  assign n6815 = ~n6813 & ~n6814;
  assign n6816 = ~n6815 & pi0937;
  assign n6817 = ~n2885 & n2717;
  assign n6818 = ~n6817 & ~n3291;
  assign n6819 = ~n6818 & ~pi0237;
  assign n6820 = ~n6816 & ~n6819;
  assign n6821 = n2885 & n2931;
  assign n6822 = ~n2885 & n2904;
  assign n6823 = ~n6821 & ~n6822;
  assign n6824 = ~n6823 & pi0273;
  assign n6825 = n3369 & pi1148;
  assign n6826 = ~n6824 & ~n6825;
  assign po0459 = ~n6820 | ~n6826;
  assign n6828 = pi0303 & pi0478;
  assign n6829 = ~pi0478 & pi1049;
  assign po0460 = n6828 | n6829;
  assign n6831 = pi0304 & pi0478;
  assign n6832 = ~pi0478 & pi1048;
  assign po0461 = n6831 | n6832;
  assign n6834 = pi0305 & pi0478;
  assign n6835 = ~pi0478 & pi1084;
  assign po0462 = n6834 | n6835;
  assign n6837 = pi0306 & pi0478;
  assign n6838 = ~pi0478 & pi1059;
  assign po0463 = n6837 | n6838;
  assign n6840 = pi0307 & pi0478;
  assign n6841 = ~pi0478 & pi1053;
  assign po0464 = n6840 | n6841;
  assign n6843 = pi0308 & pi0478;
  assign n6844 = ~pi0478 & pi1037;
  assign po0465 = n6843 | n6844;
  assign n6846 = pi0309 & pi0478;
  assign n6847 = ~pi0478 & pi1072;
  assign po0466 = n6846 | n6847;
  assign n6849 = ~n6823 & pi0271;
  assign n6850 = ~n6818 & ~pi0233;
  assign n6851 = ~n6849 & ~n6850;
  assign n6852 = n3369 & pi1147;
  assign n6853 = ~n6815 & pi0934;
  assign n6854 = ~n6852 & ~n6853;
  assign po0467 = ~n6851 | ~n6854;
  assign n6856 = n6809 & pi0301;
  assign n6857 = n6805 & n6856;
  assign n6858 = n6857 ^ ~pi0311;
  assign po0468 = n6858 & ~pi0055;
  assign n6860 = n6805 ^ ~pi0312;
  assign po0469 = ~n6860 & ~pi0055;
  assign n6862 = ~n4875 & ~n4862;
  assign n6863 = ~n6862 & ~po0740;
  assign po0634 = ~n6863 & ~n4881;
  assign n6865 = po0634 & ~pi0954;
  assign n6866 = pi0313 & pi0954;
  assign po0470 = ~n6865 & ~n6866;
  assign n6868 = n5204 & n5047;
  assign po0471 = n5229 & n6868;
  assign n6870 = po0637 & ~pi0340;
  assign n6871 = n6870 & pi1080;
  assign n6872 = ~n6870 & pi0315;
  assign po0472 = n6871 | n6872;
  assign n6874 = n6870 & pi1047;
  assign n6875 = ~n6870 & pi0316;
  assign po0473 = n6874 | n6875;
  assign n6877 = po0637 & ~pi0330;
  assign n6878 = n6877 & pi1078;
  assign n6879 = ~n6877 & pi0317;
  assign po0474 = n6878 | n6879;
  assign n6881 = po0637 & ~pi0341;
  assign n6882 = n6881 & pi1074;
  assign n6883 = ~n6881 & pi0318;
  assign po0475 = n6882 | n6883;
  assign n6885 = n6881 & pi1072;
  assign n6886 = ~n6881 & pi0319;
  assign po0476 = n6885 | n6886;
  assign n6888 = n6870 & pi1048;
  assign n6889 = ~n6870 & pi0320;
  assign po0477 = n6888 | n6889;
  assign n6891 = n6870 & pi1058;
  assign n6892 = ~n6870 & pi0321;
  assign po0478 = n6891 | n6892;
  assign n6894 = n6870 & pi1051;
  assign n6895 = ~n6870 & pi0322;
  assign po0479 = n6894 | n6895;
  assign n6897 = n6870 & pi1065;
  assign n6898 = ~n6870 & pi0323;
  assign po0480 = n6897 | n6898;
  assign n6900 = n6881 & pi1086;
  assign n6901 = ~n6881 & pi0324;
  assign po0481 = n6900 | n6901;
  assign n6903 = n6881 & pi1063;
  assign n6904 = ~n6881 & pi0325;
  assign po0482 = n6903 | n6904;
  assign n6906 = n6881 & pi1057;
  assign n6907 = ~n6881 & pi0326;
  assign po0483 = n6906 | n6907;
  assign n6909 = n6870 & pi1040;
  assign n6910 = ~n6870 & pi0327;
  assign po0484 = n6909 | n6910;
  assign n6912 = n6881 & pi1058;
  assign n6913 = ~n6881 & pi0328;
  assign po0485 = n6912 | n6913;
  assign n6915 = n6881 & pi1043;
  assign n6916 = ~n6881 & pi0329;
  assign po0486 = n6915 | n6916;
  assign n6918 = ~po0637 & ~pi0330;
  assign n6919 = ~n6870 & ~n6918;
  assign n6920 = ~n2640 & pi1092;
  assign po0487 = ~n6919 & n6920;
  assign n6922 = ~po0637 & ~pi0331;
  assign n6923 = ~n6881 & ~n6922;
  assign po0488 = ~n6923 & n6920;
  assign n6925 = n2891 & n4284;
  assign n6926 = ~n4420 & ~n4570;
  assign n6927 = n6926 & ~n2763;
  assign po0489 = n6925 | ~n6927;
  assign n6929 = n6881 & pi1040;
  assign n6930 = ~n6881 & pi0333;
  assign po0490 = n6929 | n6930;
  assign n6932 = n6881 & pi1065;
  assign n6933 = ~n6881 & pi0334;
  assign po0491 = n6932 | n6933;
  assign n6935 = n6881 & pi1069;
  assign n6936 = ~n6881 & pi0335;
  assign po0492 = n6935 | n6936;
  assign n6938 = n6877 & pi1070;
  assign n6939 = ~n6877 & pi0336;
  assign po0493 = n6938 | n6939;
  assign n6941 = n6877 & pi1044;
  assign n6942 = ~n6877 & pi0337;
  assign po0494 = n6941 | n6942;
  assign n6944 = n6877 & pi1072;
  assign n6945 = ~n6877 & pi0338;
  assign po0495 = n6944 | n6945;
  assign n6947 = n6877 & pi1086;
  assign n6948 = ~n6877 & pi0339;
  assign po0496 = n6947 | n6948;
  assign n6950 = ~po0637 & ~pi0340;
  assign n6951 = ~n6950 & n6920;
  assign n6952 = po0637 & ~pi0331;
  assign po0497 = ~n6951 | n6952;
  assign n6954 = ~po0637 & ~pi0341;
  assign n6955 = ~n6877 & ~n6954;
  assign po0498 = ~n6955 & n6920;
  assign n6957 = n6870 & pi1049;
  assign n6958 = ~n6870 & pi0342;
  assign po0499 = n6957 | n6958;
  assign n6960 = n6870 & pi1062;
  assign n6961 = ~n6870 & pi0343;
  assign po0500 = n6960 | n6961;
  assign n6963 = n6870 & pi1069;
  assign n6964 = ~n6870 & pi0344;
  assign po0501 = n6963 | n6964;
  assign n6966 = n6870 & pi1039;
  assign n6967 = ~n6870 & pi0345;
  assign po0502 = n6966 | n6967;
  assign n6969 = n6870 & pi1067;
  assign n6970 = ~n6870 & pi0346;
  assign po0503 = n6969 | n6970;
  assign n6972 = n6870 & pi1055;
  assign n6973 = ~n6870 & pi0347;
  assign po0504 = n6972 | n6973;
  assign n6975 = n6870 & pi1087;
  assign n6976 = ~n6870 & pi0348;
  assign po0505 = n6975 | n6976;
  assign n6978 = n6870 & pi1043;
  assign n6979 = ~n6870 & pi0349;
  assign po0506 = n6978 | n6979;
  assign n6981 = n6870 & pi1035;
  assign n6982 = ~n6870 & pi0350;
  assign po0507 = n6981 | n6982;
  assign n6984 = n6870 & pi1079;
  assign n6985 = ~n6870 & pi0351;
  assign po0508 = n6984 | n6985;
  assign n6987 = n6870 & pi1078;
  assign n6988 = ~n6870 & pi0352;
  assign po0509 = n6987 | n6988;
  assign n6990 = n6870 & pi1063;
  assign n6991 = ~n6870 & pi0353;
  assign po0510 = n6990 | n6991;
  assign n6993 = n6870 & pi1045;
  assign n6994 = ~n6870 & pi0354;
  assign po0511 = n6993 | n6994;
  assign n6996 = n6870 & pi1084;
  assign n6997 = ~n6870 & pi0355;
  assign po0512 = n6996 | n6997;
  assign n6999 = n6870 & pi1081;
  assign n7000 = ~n6870 & pi0356;
  assign po0513 = n6999 | n7000;
  assign n7002 = n6870 & pi1076;
  assign n7003 = ~n6870 & pi0357;
  assign po0514 = n7002 | n7003;
  assign n7005 = n6870 & pi1071;
  assign n7006 = ~n6870 & pi0358;
  assign po0515 = n7005 | n7006;
  assign n7008 = n6870 & pi1068;
  assign n7009 = ~n6870 & pi0359;
  assign po0516 = n7008 | n7009;
  assign n7011 = n6870 & pi1042;
  assign n7012 = ~n6870 & pi0360;
  assign po0517 = n7011 | n7012;
  assign n7014 = n6870 & pi1059;
  assign n7015 = ~n6870 & pi0361;
  assign po0518 = n7014 | n7015;
  assign n7017 = n6870 & pi1070;
  assign n7018 = ~n6870 & pi0362;
  assign po0519 = n7017 | n7018;
  assign n7020 = n6877 & pi1049;
  assign n7021 = ~n6877 & pi0363;
  assign po0520 = n7020 | n7021;
  assign n7023 = n6877 & pi1062;
  assign n7024 = ~n6877 & pi0364;
  assign po0521 = n7023 | n7024;
  assign n7026 = n6877 & pi1065;
  assign n7027 = ~n6877 & pi0365;
  assign po0522 = n7026 | n7027;
  assign n7029 = n6877 & pi1069;
  assign n7030 = ~n6877 & pi0366;
  assign po0523 = n7029 | n7030;
  assign n7032 = n6877 & pi1039;
  assign n7033 = ~n6877 & pi0367;
  assign po0524 = n7032 | n7033;
  assign n7035 = n6877 & pi1067;
  assign n7036 = ~n6877 & pi0368;
  assign po0525 = n7035 | n7036;
  assign n7038 = n6877 & pi1080;
  assign n7039 = ~n6877 & pi0369;
  assign po0526 = n7038 | n7039;
  assign n7041 = n6877 & pi1055;
  assign n7042 = ~n6877 & pi0370;
  assign po0527 = n7041 | n7042;
  assign n7044 = n6877 & pi1051;
  assign n7045 = ~n6877 & pi0371;
  assign po0528 = n7044 | n7045;
  assign n7047 = n6877 & pi1048;
  assign n7048 = ~n6877 & pi0372;
  assign po0529 = n7047 | n7048;
  assign n7050 = n6877 & pi1087;
  assign n7051 = ~n6877 & pi0373;
  assign po0530 = n7050 | n7051;
  assign n7053 = n6877 & pi1035;
  assign n7054 = ~n6877 & pi0374;
  assign po0531 = n7053 | n7054;
  assign n7056 = n6877 & pi1047;
  assign n7057 = ~n6877 & pi0375;
  assign po0532 = n7056 | n7057;
  assign n7059 = n6877 & pi1079;
  assign n7060 = ~n6877 & pi0376;
  assign po0533 = n7059 | n7060;
  assign n7062 = n6877 & pi1074;
  assign n7063 = ~n6877 & pi0377;
  assign po0534 = n7062 | n7063;
  assign n7065 = n6877 & pi1063;
  assign n7066 = ~n6877 & pi0378;
  assign po0535 = n7065 | n7066;
  assign n7068 = n6877 & pi1045;
  assign n7069 = ~n6877 & pi0379;
  assign po0536 = n7068 | n7069;
  assign n7071 = n6877 & pi1084;
  assign n7072 = ~n6877 & pi0380;
  assign po0537 = n7071 | n7072;
  assign n7074 = n6877 & pi1081;
  assign n7075 = ~n6877 & pi0381;
  assign po0538 = n7074 | n7075;
  assign n7077 = n6877 & pi1076;
  assign n7078 = ~n6877 & pi0382;
  assign po0539 = n7077 | n7078;
  assign n7080 = n6877 & pi1071;
  assign n7081 = ~n6877 & pi0383;
  assign po0540 = n7080 | n7081;
  assign n7083 = n6877 & pi1068;
  assign n7084 = ~n6877 & pi0384;
  assign po0541 = n7083 | n7084;
  assign n7086 = n6877 & pi1042;
  assign n7087 = ~n6877 & pi0385;
  assign po0542 = n7086 | n7087;
  assign n7089 = n6877 & pi1059;
  assign n7090 = ~n6877 & pi0386;
  assign po0543 = n7089 | n7090;
  assign n7092 = n6877 & pi1053;
  assign n7093 = ~n6877 & pi0387;
  assign po0544 = n7092 | n7093;
  assign n7095 = n6877 & pi1037;
  assign n7096 = ~n6877 & pi0388;
  assign po0545 = n7095 | n7096;
  assign n7098 = n6877 & pi1036;
  assign n7099 = ~n6877 & pi0389;
  assign po0546 = n7098 | n7099;
  assign n7101 = n6881 & pi1049;
  assign n7102 = ~n6881 & pi0390;
  assign po0547 = n7101 | n7102;
  assign n7104 = n6881 & pi1062;
  assign n7105 = ~n6881 & pi0391;
  assign po0548 = n7104 | n7105;
  assign n7107 = n6881 & pi1039;
  assign n7108 = ~n6881 & pi0392;
  assign po0549 = n7107 | n7108;
  assign n7110 = n6881 & pi1067;
  assign n7111 = ~n6881 & pi0393;
  assign po0550 = n7110 | n7111;
  assign n7113 = n6881 & pi1080;
  assign n7114 = ~n6881 & pi0394;
  assign po0551 = n7113 | n7114;
  assign n7116 = n6881 & pi1055;
  assign n7117 = ~n6881 & pi0395;
  assign po0552 = n7116 | n7117;
  assign n7119 = n6881 & pi1051;
  assign n7120 = ~n6881 & pi0396;
  assign po0553 = n7119 | n7120;
  assign n7122 = n6881 & pi1048;
  assign n7123 = ~n6881 & pi0397;
  assign po0554 = n7122 | n7123;
  assign n7125 = n6881 & pi1087;
  assign n7126 = ~n6881 & pi0398;
  assign po0555 = n7125 | n7126;
  assign n7128 = n6881 & pi1047;
  assign n7129 = ~n6881 & pi0399;
  assign po0556 = n7128 | n7129;
  assign n7131 = n6881 & pi1035;
  assign n7132 = ~n6881 & pi0400;
  assign po0557 = n7131 | n7132;
  assign n7134 = n6881 & pi1079;
  assign n7135 = ~n6881 & pi0401;
  assign po0558 = n7134 | n7135;
  assign n7137 = n6881 & pi1078;
  assign n7138 = ~n6881 & pi0402;
  assign po0559 = n7137 | n7138;
  assign n7140 = n6881 & pi1045;
  assign n7141 = ~n6881 & pi0403;
  assign po0560 = n7140 | n7141;
  assign n7143 = n6881 & pi1084;
  assign n7144 = ~n6881 & pi0404;
  assign po0561 = n7143 | n7144;
  assign n7146 = n6881 & pi1081;
  assign n7147 = ~n6881 & pi0405;
  assign po0562 = n7146 | n7147;
  assign n7149 = n6881 & pi1076;
  assign n7150 = ~n6881 & pi0406;
  assign po0563 = n7149 | n7150;
  assign n7152 = n6881 & pi1071;
  assign n7153 = ~n6881 & pi0407;
  assign po0564 = n7152 | n7153;
  assign n7155 = n6881 & pi1068;
  assign n7156 = ~n6881 & pi0408;
  assign po0565 = n7155 | n7156;
  assign n7158 = n6881 & pi1042;
  assign n7159 = ~n6881 & pi0409;
  assign po0566 = n7158 | n7159;
  assign n7161 = n6881 & pi1059;
  assign n7162 = ~n6881 & pi0410;
  assign po0567 = n7161 | n7162;
  assign n7164 = n6881 & pi1053;
  assign n7165 = ~n6881 & pi0411;
  assign po0568 = n7164 | n7165;
  assign n7167 = n6881 & pi1037;
  assign n7168 = ~n6881 & pi0412;
  assign po0569 = n7167 | n7168;
  assign n7170 = n6881 & pi1036;
  assign n7171 = ~n6881 & pi0413;
  assign po0570 = n7170 | n7171;
  assign n7173 = n6952 & pi1049;
  assign n7174 = ~n6952 & pi0414;
  assign po0571 = n7173 | n7174;
  assign n7176 = n6952 & pi1062;
  assign n7177 = ~n6952 & pi0415;
  assign po0572 = n7176 | n7177;
  assign n7179 = n6952 & pi1069;
  assign n7180 = ~n6952 & pi0416;
  assign po0573 = n7179 | n7180;
  assign n7182 = n6952 & pi1039;
  assign n7183 = ~n6952 & pi0417;
  assign po0574 = n7182 | n7183;
  assign n7185 = n6952 & pi1067;
  assign n7186 = ~n6952 & pi0418;
  assign po0575 = n7185 | n7186;
  assign n7188 = n6952 & pi1080;
  assign n7189 = ~n6952 & pi0419;
  assign po0576 = n7188 | n7189;
  assign n7191 = n6952 & pi1055;
  assign n7192 = ~n6952 & pi0420;
  assign po0577 = n7191 | n7192;
  assign n7194 = n6952 & pi1051;
  assign n7195 = ~n6952 & pi0421;
  assign po0578 = n7194 | n7195;
  assign n7197 = n6952 & pi1048;
  assign n7198 = ~n6952 & pi0422;
  assign po0579 = n7197 | n7198;
  assign n7200 = n6952 & pi1087;
  assign n7201 = ~n6952 & pi0423;
  assign po0580 = n7200 | n7201;
  assign n7203 = n6952 & pi1047;
  assign n7204 = ~n6952 & pi0424;
  assign po0581 = n7203 | n7204;
  assign n7206 = n6952 & pi1035;
  assign n7207 = ~n6952 & pi0425;
  assign po0582 = n7206 | n7207;
  assign n7209 = n6952 & pi1079;
  assign n7210 = ~n6952 & pi0426;
  assign po0583 = n7209 | n7210;
  assign n7212 = n6952 & pi1078;
  assign n7213 = ~n6952 & pi0427;
  assign po0584 = n7212 | n7213;
  assign n7215 = n6952 & pi1045;
  assign n7216 = ~n6952 & pi0428;
  assign po0585 = n7215 | n7216;
  assign n7218 = n6952 & pi1084;
  assign n7219 = ~n6952 & pi0429;
  assign po0586 = n7218 | n7219;
  assign n7221 = n6952 & pi1076;
  assign n7222 = ~n6952 & pi0430;
  assign po0587 = n7221 | n7222;
  assign n7224 = n6952 & pi1071;
  assign n7225 = ~n6952 & pi0431;
  assign po0588 = n7224 | n7225;
  assign n7227 = n6952 & pi1068;
  assign n7228 = ~n6952 & pi0432;
  assign po0589 = n7227 | n7228;
  assign n7230 = n6952 & pi1042;
  assign n7231 = ~n6952 & pi0433;
  assign po0590 = n7230 | n7231;
  assign n7233 = n6952 & pi1059;
  assign n7234 = ~n6952 & pi0434;
  assign po0591 = n7233 | n7234;
  assign n7236 = n6952 & pi1053;
  assign n7237 = ~n6952 & pi0435;
  assign po0592 = n7236 | n7237;
  assign n7239 = n6952 & pi1037;
  assign n7240 = ~n6952 & pi0436;
  assign po0593 = n7239 | n7240;
  assign n7242 = n6952 & pi1070;
  assign n7243 = ~n6952 & pi0437;
  assign po0594 = n7242 | n7243;
  assign n7245 = n6952 & pi1036;
  assign n7246 = ~n6952 & pi0438;
  assign po0595 = n7245 | n7246;
  assign n7248 = n6877 & pi1057;
  assign n7249 = ~n6877 & pi0439;
  assign po0596 = n7248 | n7249;
  assign n7251 = n6877 & pi1043;
  assign n7252 = ~n6877 & pi0440;
  assign po0597 = n7251 | n7252;
  assign n7254 = n6870 & pi1044;
  assign n7255 = ~n6870 & pi0441;
  assign po0598 = n7254 | n7255;
  assign n7257 = n6877 & pi1058;
  assign n7258 = ~n6877 & pi0442;
  assign po0599 = n7257 | n7258;
  assign n7260 = n6952 & pi1044;
  assign n7261 = ~n6952 & pi0443;
  assign po0600 = n7260 | n7261;
  assign n7263 = n6952 & pi1072;
  assign n7264 = ~n6952 & pi0444;
  assign po0601 = n7263 | n7264;
  assign n7266 = n6952 & pi1081;
  assign n7267 = ~n6952 & pi0445;
  assign po0602 = n7266 | n7267;
  assign n7269 = n6952 & pi1086;
  assign n7270 = ~n6952 & pi0446;
  assign po0603 = n7269 | n7270;
  assign n7272 = n6877 & pi1040;
  assign n7273 = ~n6877 & pi0447;
  assign po0604 = n7272 | n7273;
  assign n7275 = n6952 & pi1074;
  assign n7276 = ~n6952 & pi0448;
  assign po0605 = n7275 | n7276;
  assign n7278 = n6952 & pi1057;
  assign n7279 = ~n6952 & pi0449;
  assign po0606 = n7278 | n7279;
  assign n7281 = n6870 & pi1036;
  assign n7282 = ~n6870 & pi0450;
  assign po0607 = n7281 | n7282;
  assign n7284 = n6952 & pi1063;
  assign n7285 = ~n6952 & pi0451;
  assign po0608 = n7284 | n7285;
  assign n7287 = n6870 & pi1053;
  assign n7288 = ~n6870 & pi0452;
  assign po0609 = n7287 | n7288;
  assign n7290 = n6952 & pi1040;
  assign n7291 = ~n6952 & pi0453;
  assign po0610 = n7290 | n7291;
  assign n7293 = n6952 & pi1043;
  assign n7294 = ~n6952 & pi0454;
  assign po0611 = n7293 | n7294;
  assign n7296 = n6870 & pi1037;
  assign n7297 = ~n6870 & pi0455;
  assign po0612 = n7296 | n7297;
  assign n7299 = n6881 & pi1044;
  assign n7300 = ~n6881 & pi0456;
  assign po0613 = n7299 | n7300;
  assign n7302 = pi0599 & pi0815;
  assign n7303 = ~n7302 & pi0810;
  assign n7304 = ~n7303 & pi0596;
  assign n7305 = ~n7304 & pi0804;
  assign n7306 = pi0594 & pi0600;
  assign n7307 = pi0597 & pi0601;
  assign n7308 = n7306 & n7307;
  assign n7309 = ~pi0804 & ~pi0810;
  assign n7310 = ~n7309 & ~pi0595;
  assign n7311 = n7308 & ~n7310;
  assign n7312 = ~n7305 & n7311;
  assign n7313 = ~n7309 & ~pi0601;
  assign n7314 = ~n7313 & ~pi0815;
  assign n7315 = pi0600 & ~pi0810;
  assign n7316 = ~n7315 & pi0804;
  assign n7317 = n7314 & ~n7316;
  assign n7318 = ~n7312 & ~n7317;
  assign n7319 = ~n7318 & pi0605;
  assign n7320 = ~pi0815 & pi0990;
  assign n7321 = n7306 & n7320;
  assign n7322 = n7316 & n7321;
  assign n7323 = ~n7319 & ~n7322;
  assign po0614 = ~n7323 & pi0821;
  assign n7325 = n6870 & pi1072;
  assign n7326 = ~n6870 & pi0458;
  assign po0615 = n7325 | n7326;
  assign n7328 = n6952 & pi1058;
  assign n7329 = ~n6952 & pi0459;
  assign po0616 = n7328 | n7329;
  assign n7331 = n6870 & pi1086;
  assign n7332 = ~n6870 & pi0460;
  assign po0617 = n7331 | n7332;
  assign n7334 = n6870 & pi1057;
  assign n7335 = ~n6870 & pi0461;
  assign po0618 = n7334 | n7335;
  assign n7337 = n6870 & pi1074;
  assign n7338 = ~n6870 & pi0462;
  assign po0619 = n7337 | n7338;
  assign n7340 = n6881 & pi1070;
  assign n7341 = ~n6881 & pi0463;
  assign po0620 = n7340 | n7341;
  assign n7343 = n6952 & pi1065;
  assign n7344 = ~n6952 & pi0464;
  assign po0621 = n7343 | n7344;
  assign n7346 = ~n6823 & ~pi0243;
  assign n7347 = ~n6815 & pi0926;
  assign n7348 = ~n7346 & ~n7347;
  assign n7349 = n3369 & pi1157;
  assign po0622 = ~n7348 | n7349;
  assign n7351 = ~n6823 & pi0275;
  assign n7352 = ~n6815 & pi0943;
  assign n7353 = ~n7351 & ~n7352;
  assign n7354 = n3369 & pi1151;
  assign po0623 = ~n7353 | n7354;
  assign n7356 = n4536 & n6048;
  assign n7357 = pi0040 & pi1001;
  assign n7358 = n3416 & n7357;
  assign n7359 = po0950 & n7358;
  assign po0624 = n7356 | n7359;
  assign n7361 = n2763 & ~pi0024;
  assign n7362 = ~n7361 & pi0468;
  assign po0625 = n7362 | n4515;
  assign n7364 = ~n6815 & pi0942;
  assign n7365 = ~n6823 & ~pi0263;
  assign n7366 = ~n7364 & ~n7365;
  assign n7367 = n3369 & pi1156;
  assign po0626 = ~n7366 | n7367;
  assign n7369 = ~n6815 & pi0925;
  assign n7370 = ~n6823 & pi0267;
  assign n7371 = ~n7369 & ~n7370;
  assign n7372 = n3369 & pi1155;
  assign po0627 = ~n7371 | n7372;
  assign n7374 = ~n6815 & pi0941;
  assign n7375 = ~n6823 & pi0253;
  assign n7376 = ~n7374 & ~n7375;
  assign n7377 = n3369 & pi1153;
  assign po0628 = ~n7376 | n7377;
  assign n7379 = ~n6823 & pi0254;
  assign n7380 = ~n6815 & pi0923;
  assign n7381 = ~n7379 & ~n7380;
  assign n7382 = n3369 & pi1154;
  assign po0629 = ~n7381 | n7382;
  assign n7384 = ~n6815 & pi0922;
  assign n7385 = ~n6823 & pi0268;
  assign n7386 = ~n7384 & ~n7385;
  assign n7387 = n3369 & pi1152;
  assign po0630 = ~n7386 | n7387;
  assign n7389 = ~n6815 & pi0931;
  assign n7390 = ~n6823 & pi0272;
  assign n7391 = ~n7389 & ~n7390;
  assign n7392 = n3369 & pi1150;
  assign po0631 = ~n7391 | n7392;
  assign n7394 = ~n6815 & pi0936;
  assign n7395 = ~n6823 & pi0283;
  assign n7396 = ~n7394 & ~n7395;
  assign n7397 = n3369 & pi1149;
  assign po0632 = ~n7396 | n7397;
  assign n7399 = n6376 & pi0071;
  assign po0633 = n4761 | n7399;
  assign po0635 = n6372 & pi0071;
  assign n7402 = n5861 & pi0248;
  assign n7403 = ~n5861 & pi0481;
  assign po0638 = n7402 | n7403;
  assign n7405 = n5876 & pi0249;
  assign n7406 = ~n5876 & pi0482;
  assign po0639 = n7405 | n7406;
  assign n7408 = n5898 & pi0242;
  assign n7409 = ~n5898 & pi0483;
  assign po0640 = n7408 | n7409;
  assign n7411 = n5898 & pi0249;
  assign n7412 = ~n5898 & pi0484;
  assign po0641 = n7411 | n7412;
  assign n7414 = n5968 & pi0234;
  assign n7415 = ~n5968 & pi0485;
  assign po0642 = n7414 | n7415;
  assign n7417 = n5968 & pi0244;
  assign n7418 = ~n5968 & pi0486;
  assign po0643 = n7417 | n7418;
  assign n7420 = n5861 & pi0246;
  assign n7421 = ~n5861 & pi0487;
  assign po0644 = n7420 | n7421;
  assign n7423 = ~n5861 & pi0488;
  assign n7424 = n5861 & ~pi0239;
  assign po0645 = ~n7423 & ~n7424;
  assign n7426 = n5968 & pi0242;
  assign n7427 = ~n5968 & pi0489;
  assign po0646 = n7426 | n7427;
  assign n7429 = n5898 & pi0241;
  assign n7430 = ~n5898 & pi0490;
  assign po0647 = n7429 | n7430;
  assign n7432 = n5898 & pi0238;
  assign n7433 = ~n5898 & pi0491;
  assign po0648 = n7432 | n7433;
  assign n7435 = n5898 & pi0240;
  assign n7436 = ~n5898 & pi0492;
  assign po0649 = n7435 | n7436;
  assign n7438 = n5898 & pi0244;
  assign n7439 = ~n5898 & pi0493;
  assign po0650 = n7438 | n7439;
  assign n7441 = ~n5898 & pi0494;
  assign n7442 = n5898 & ~pi0239;
  assign po0651 = ~n7441 & ~n7442;
  assign n7444 = n5898 & pi0235;
  assign n7445 = ~n5898 & pi0495;
  assign po0652 = n7444 | n7445;
  assign n7447 = n5891 & pi0249;
  assign n7448 = ~n5891 & pi0496;
  assign po0653 = n7447 | n7448;
  assign n7450 = ~n5891 & pi0497;
  assign n7451 = n5891 & ~pi0239;
  assign po0654 = ~n7450 & ~n7451;
  assign n7453 = n5876 & pi0238;
  assign n7454 = ~n5876 & pi0498;
  assign po0655 = n7453 | n7454;
  assign n7456 = n5891 & pi0246;
  assign n7457 = ~n5891 & pi0499;
  assign po0656 = n7456 | n7457;
  assign n7459 = n5891 & pi0241;
  assign n7460 = ~n5891 & pi0500;
  assign po0657 = n7459 | n7460;
  assign n7462 = n5891 & pi0248;
  assign n7463 = ~n5891 & pi0501;
  assign po0658 = n7462 | n7463;
  assign n7465 = n5891 & pi0247;
  assign n7466 = ~n5891 & pi0502;
  assign po0659 = n7465 | n7466;
  assign n7468 = n5891 & pi0245;
  assign n7469 = ~n5891 & pi0503;
  assign po0660 = n7468 | n7469;
  assign n7471 = n5887 & pi0242;
  assign n7472 = ~n5887 & pi0504;
  assign po0661 = n7471 | n7472;
  assign n7474 = n5891 & pi0234;
  assign n7475 = ~n5891 & pi0505;
  assign po0662 = n7474 | n7475;
  assign n7477 = n5887 & pi0241;
  assign n7478 = ~n5887 & pi0506;
  assign po0663 = n7477 | n7478;
  assign n7480 = n5887 & pi0238;
  assign n7481 = ~n5887 & pi0507;
  assign po0664 = n7480 | n7481;
  assign n7483 = n5887 & pi0247;
  assign n7484 = ~n5887 & pi0508;
  assign po0665 = n7483 | n7484;
  assign n7486 = n5887 & pi0245;
  assign n7487 = ~n5887 & pi0509;
  assign po0666 = n7486 | n7487;
  assign n7489 = n5861 & pi0242;
  assign n7490 = ~n5861 & pi0510;
  assign po0667 = n7489 | n7490;
  assign n7492 = n5861 & pi0234;
  assign n7493 = ~n5861 & pi0511;
  assign po0668 = n7492 | n7493;
  assign n7495 = n5861 & pi0235;
  assign n7496 = ~n5861 & pi0512;
  assign po0669 = n7495 | n7496;
  assign n7498 = n5861 & pi0244;
  assign n7499 = ~n5861 & pi0513;
  assign po0670 = n7498 | n7499;
  assign n7501 = n5861 & pi0245;
  assign n7502 = ~n5861 & pi0514;
  assign po0671 = n7501 | n7502;
  assign n7504 = n5861 & pi0240;
  assign n7505 = ~n5861 & pi0515;
  assign po0672 = n7504 | n7505;
  assign n7507 = n5861 & pi0247;
  assign n7508 = ~n5861 & pi0516;
  assign po0673 = n7507 | n7508;
  assign n7510 = n5861 & pi0238;
  assign n7511 = ~n5861 & pi0517;
  assign po0674 = n7510 | n7511;
  assign n7513 = n5869 & pi0234;
  assign n7514 = ~n5869 & pi0518;
  assign po0675 = n7513 | n7514;
  assign n7516 = ~n5869 & pi0519;
  assign n7517 = n5869 & ~pi0239;
  assign po0676 = ~n7516 & ~n7517;
  assign n7519 = n5869 & pi0246;
  assign n7520 = ~n5869 & pi0520;
  assign po0677 = n7519 | n7520;
  assign n7522 = n5869 & pi0248;
  assign n7523 = ~n5869 & pi0521;
  assign po0678 = n7522 | n7523;
  assign n7525 = n5869 & pi0238;
  assign n7526 = ~n5869 & pi0522;
  assign po0679 = n7525 | n7526;
  assign n7528 = n5978 & pi0234;
  assign n7529 = ~n5978 & pi0523;
  assign po0680 = n7528 | n7529;
  assign n7531 = ~n5978 & pi0524;
  assign n7532 = n5978 & ~pi0239;
  assign po0681 = ~n7531 & ~n7532;
  assign n7534 = n5978 & pi0245;
  assign n7535 = ~n5978 & pi0525;
  assign po0682 = n7534 | n7535;
  assign n7537 = n5978 & pi0246;
  assign n7538 = ~n5978 & pi0526;
  assign po0683 = n7537 | n7538;
  assign n7540 = n5978 & pi0247;
  assign n7541 = ~n5978 & pi0527;
  assign po0684 = n7540 | n7541;
  assign n7543 = n5978 & pi0249;
  assign n7544 = ~n5978 & pi0528;
  assign po0685 = n7543 | n7544;
  assign n7546 = n5978 & pi0238;
  assign n7547 = ~n5978 & pi0529;
  assign po0686 = n7546 | n7547;
  assign n7549 = n5978 & pi0240;
  assign n7550 = ~n5978 & pi0530;
  assign po0687 = n7549 | n7550;
  assign n7552 = n5876 & pi0235;
  assign n7553 = ~n5876 & pi0531;
  assign po0688 = n7552 | n7553;
  assign n7555 = n5876 & pi0247;
  assign n7556 = ~n5876 & pi0532;
  assign po0689 = n7555 | n7556;
  assign n7558 = n5887 & pi0235;
  assign n7559 = ~n5887 & pi0533;
  assign po0690 = n7558 | n7559;
  assign n7561 = ~n5887 & pi0534;
  assign n7562 = n5887 & ~pi0239;
  assign po0691 = ~n7561 & ~n7562;
  assign n7564 = n5887 & pi0240;
  assign n7565 = ~n5887 & pi0535;
  assign po0692 = n7564 | n7565;
  assign n7567 = n5887 & pi0246;
  assign n7568 = ~n5887 & pi0536;
  assign po0693 = n7567 | n7568;
  assign n7570 = n5887 & pi0248;
  assign n7571 = ~n5887 & pi0537;
  assign po0694 = n7570 | n7571;
  assign n7573 = n5887 & pi0249;
  assign n7574 = ~n5887 & pi0538;
  assign po0695 = n7573 | n7574;
  assign n7576 = n5891 & pi0242;
  assign n7577 = ~n5891 & pi0539;
  assign po0696 = n7576 | n7577;
  assign n7579 = n5891 & pi0235;
  assign n7580 = ~n5891 & pi0540;
  assign po0697 = n7579 | n7580;
  assign n7582 = n5891 & pi0244;
  assign n7583 = ~n5891 & pi0541;
  assign po0698 = n7582 | n7583;
  assign n7585 = n5891 & pi0240;
  assign n7586 = ~n5891 & pi0542;
  assign po0699 = n7585 | n7586;
  assign n7588 = n5891 & pi0238;
  assign n7589 = ~n5891 & pi0543;
  assign po0700 = n7588 | n7589;
  assign n7591 = n5898 & pi0234;
  assign n7592 = ~n5898 & pi0544;
  assign po0701 = n7591 | n7592;
  assign n7594 = n5898 & pi0245;
  assign n7595 = ~n5898 & pi0545;
  assign po0702 = n7594 | n7595;
  assign n7597 = n5898 & pi0246;
  assign n7598 = ~n5898 & pi0546;
  assign po0703 = n7597 | n7598;
  assign n7600 = n5898 & pi0247;
  assign n7601 = ~n5898 & pi0547;
  assign po0704 = n7600 | n7601;
  assign n7603 = n5898 & pi0248;
  assign n7604 = ~n5898 & pi0548;
  assign po0705 = n7603 | n7604;
  assign n7606 = n5968 & pi0235;
  assign n7607 = ~n5968 & pi0549;
  assign po0706 = n7606 | n7607;
  assign n7609 = ~n5968 & pi0550;
  assign n7610 = n5968 & ~pi0239;
  assign po0707 = ~n7609 & ~n7610;
  assign n7612 = n5968 & pi0240;
  assign n7613 = ~n5968 & pi0551;
  assign po0708 = n7612 | n7613;
  assign n7615 = n5968 & pi0247;
  assign n7616 = ~n5968 & pi0552;
  assign po0709 = n7615 | n7616;
  assign n7618 = n5968 & pi0241;
  assign n7619 = ~n5968 & pi0553;
  assign po0710 = n7618 | n7619;
  assign n7621 = n5968 & pi0248;
  assign n7622 = ~n5968 & pi0554;
  assign po0711 = n7621 | n7622;
  assign n7624 = n5968 & pi0249;
  assign n7625 = ~n5968 & pi0555;
  assign po0712 = n7624 | n7625;
  assign n7627 = n5876 & pi0242;
  assign n7628 = ~n5876 & pi0556;
  assign po0713 = n7627 | n7628;
  assign n7630 = n5887 & pi0234;
  assign n7631 = ~n5887 & pi0557;
  assign po0714 = n7630 | n7631;
  assign n7633 = n5887 & pi0244;
  assign n7634 = ~n5887 & pi0558;
  assign po0715 = n7633 | n7634;
  assign n7636 = n5861 & pi0241;
  assign n7637 = ~n5861 & pi0559;
  assign po0716 = n7636 | n7637;
  assign n7639 = n5876 & pi0240;
  assign n7640 = ~n5876 & pi0560;
  assign po0717 = n7639 | n7640;
  assign n7642 = n5869 & pi0247;
  assign n7643 = ~n5869 & pi0561;
  assign po0718 = n7642 | n7643;
  assign n7645 = n5876 & pi0241;
  assign n7646 = ~n5876 & pi0562;
  assign po0719 = n7645 | n7646;
  assign n7648 = n5968 & pi0246;
  assign n7649 = ~n5968 & pi0563;
  assign po0720 = n7648 | n7649;
  assign n7651 = n5876 & pi0246;
  assign n7652 = ~n5876 & pi0564;
  assign po0721 = n7651 | n7652;
  assign n7654 = n5876 & pi0248;
  assign n7655 = ~n5876 & pi0565;
  assign po0722 = n7654 | n7655;
  assign n7657 = n5876 & pi0244;
  assign n7658 = ~n5876 & pi0566;
  assign po0723 = n7657 | n7658;
  assign n7660 = n5450 & pi0665;
  assign n7661 = n5424 & pi0621;
  assign n7662 = ~n7660 & ~n7661;
  assign n7663 = pi0230 & pi1093;
  assign n7664 = n7663 & pi1091;
  assign n7665 = ~n7662 & n7664;
  assign n7666 = ~n7663 & ~pi0567;
  assign n7667 = ~n7665 & ~n7666;
  assign po0724 = ~n7667 & pi1092;
  assign n7669 = n5876 & pi0245;
  assign n7670 = ~n5876 & pi0568;
  assign po0725 = n7669 | n7670;
  assign n7672 = ~n5876 & pi0569;
  assign n7673 = n5876 & ~pi0239;
  assign po0726 = ~n7672 & ~n7673;
  assign n7675 = n5876 & pi0234;
  assign n7676 = ~n5876 & pi0570;
  assign po0727 = n7675 | n7676;
  assign n7678 = n5978 & pi0241;
  assign n7679 = ~n5978 & pi0571;
  assign po0728 = n7678 | n7679;
  assign n7681 = n5978 & pi0244;
  assign n7682 = ~n5978 & pi0572;
  assign po0729 = n7681 | n7682;
  assign n7684 = n5978 & pi0242;
  assign n7685 = ~n5978 & pi0573;
  assign po0730 = n7684 | n7685;
  assign n7687 = n5869 & pi0241;
  assign n7688 = ~n5869 & pi0574;
  assign po0731 = n7687 | n7688;
  assign n7690 = n5978 & pi0235;
  assign n7691 = ~n5978 & pi0575;
  assign po0732 = n7690 | n7691;
  assign n7693 = n5978 & pi0248;
  assign n7694 = ~n5978 & pi0576;
  assign po0733 = n7693 | n7694;
  assign n7696 = n5968 & pi0238;
  assign n7697 = ~n5968 & pi0577;
  assign po0734 = n7696 | n7697;
  assign n7699 = n5869 & pi0249;
  assign n7700 = ~n5869 & pi0578;
  assign po0735 = n7699 | n7700;
  assign n7702 = n5861 & pi0249;
  assign n7703 = ~n5861 & pi0579;
  assign po0736 = n7702 | n7703;
  assign n7705 = n5968 & pi0245;
  assign n7706 = ~n5968 & pi0580;
  assign po0737 = n7705 | n7706;
  assign n7708 = n5869 & pi0235;
  assign n7709 = ~n5869 & pi0581;
  assign po0738 = n7708 | n7709;
  assign n7711 = n5869 & pi0240;
  assign n7712 = ~n5869 & pi0582;
  assign po0739 = n7711 | n7712;
  assign n7714 = n5869 & pi0245;
  assign n7715 = ~n5869 & pi0584;
  assign po0741 = n7714 | n7715;
  assign n7717 = n5869 & pi0244;
  assign n7718 = ~n5869 & pi0585;
  assign po0742 = n7717 | n7718;
  assign n7720 = n5869 & pi0242;
  assign n7721 = ~n5869 & pi0586;
  assign po0743 = n7720 | n7721;
  assign n7723 = n5426 & pi0230;
  assign n7724 = ~pi0230 & pi0587;
  assign po0744 = n7723 | n7724;
  assign n7726 = ~pi0123 & pi0824;
  assign n7727 = n7726 & pi0950;
  assign n7728 = ~n7727 & ~pi0588;
  assign n7729 = ~n7728 & n6920;
  assign n7730 = n7727 & ~pi0591;
  assign po0745 = n7729 & ~n7730;
  assign n7732 = pi0204 & pi0237;
  assign n7733 = ~n7732 & pi0233;
  assign n7734 = pi0206 & ~pi0237;
  assign n7735 = n7733 & ~n7734;
  assign n7736 = pi0218 & ~pi0237;
  assign n7737 = pi0205 & pi0237;
  assign n7738 = ~n7736 & ~n7737;
  assign n7739 = n7738 & ~pi0233;
  assign n7740 = ~n7735 & ~n7739;
  assign n7741 = ~n5882 & ~n7740;
  assign n7742 = pi0201 & pi0237;
  assign n7743 = ~n7742 & pi0233;
  assign n7744 = pi0220 & ~pi0237;
  assign n7745 = n7743 & ~n7744;
  assign n7746 = pi0203 & ~pi0237;
  assign n7747 = pi0202 & pi0237;
  assign n7748 = ~n7746 & ~n7747;
  assign n7749 = n7748 & ~pi0233;
  assign n7750 = ~n7745 & ~n7749;
  assign n7751 = n5855 & ~n7750;
  assign po0746 = n7741 | n7751;
  assign n7753 = n7727 & pi0588;
  assign n7754 = ~n7753 & n6920;
  assign n7755 = ~n7727 & pi0590;
  assign po0747 = ~n7754 | n7755;
  assign n7757 = ~n7727 & ~pi0591;
  assign n7758 = ~n7757 & n6920;
  assign n7759 = n7727 & ~pi0592;
  assign po0748 = n7758 & ~n7759;
  assign n7761 = ~n7727 & ~pi0592;
  assign n7762 = ~n7761 & n6920;
  assign n7763 = n7727 & ~pi0590;
  assign po0749 = n7762 & ~n7763;
  assign n7765 = ~pi0238 & pi0507;
  assign n7766 = ~n7765 & pi0233;
  assign n7767 = pi0249 ^ ~pi0538;
  assign n7768 = n7766 & n7767;
  assign n7769 = pi0242 ^ ~pi0504;
  assign n7770 = pi0235 ^ ~pi0533;
  assign n7771 = n7769 & n7770;
  assign n7772 = n7768 & n7771;
  assign n7773 = pi0238 & ~pi0507;
  assign n7774 = pi0247 ^ ~pi0508;
  assign n7775 = ~n7773 & n7774;
  assign n7776 = n7772 & n7775;
  assign n7777 = ~pi0240 ^ ~pi0535;
  assign n7778 = pi0234 ^ ~pi0557;
  assign n7779 = ~n7777 & n7778;
  assign n7780 = ~pi0244 ^ ~pi0558;
  assign n7781 = pi0241 ^ ~pi0506;
  assign n7782 = ~n7780 & n7781;
  assign n7783 = n7779 & n7782;
  assign n7784 = ~pi0248 ^ ~pi0537;
  assign n7785 = pi0245 ^ ~pi0509;
  assign n7786 = ~n7784 & n7785;
  assign n7787 = ~pi0246 ^ ~pi0536;
  assign n7788 = ~pi0239 ^ ~pi0534;
  assign n7789 = ~n7787 & n7788;
  assign n7790 = n7786 & n7789;
  assign n7791 = n7783 & n7790;
  assign n7792 = n7776 & n7791;
  assign n7793 = ~pi0245 & pi0503;
  assign n7794 = ~pi0246 & pi0499;
  assign n7795 = ~n7793 & ~n7794;
  assign n7796 = pi0241 & ~pi0500;
  assign n7797 = pi0242 ^ ~pi0539;
  assign n7798 = ~n7796 & n7797;
  assign n7799 = n7795 & n7798;
  assign n7800 = pi0249 ^ ~pi0496;
  assign n7801 = n7800 & ~pi0233;
  assign n7802 = n7799 & n7801;
  assign n7803 = pi0246 & ~pi0499;
  assign n7804 = ~pi0241 & pi0500;
  assign n7805 = ~n7803 & ~n7804;
  assign n7806 = pi0245 & ~pi0503;
  assign n7807 = n7805 & ~n7806;
  assign n7808 = n7802 & n7807;
  assign n7809 = ~pi0238 ^ ~pi0543;
  assign n7810 = pi0248 ^ ~pi0501;
  assign n7811 = ~n7809 & n7810;
  assign n7812 = ~pi0235 ^ ~pi0540;
  assign n7813 = pi0247 ^ ~pi0502;
  assign n7814 = ~n7812 & n7813;
  assign n7815 = n7811 & n7814;
  assign n7816 = ~pi0244 ^ ~pi0541;
  assign n7817 = pi0234 ^ ~pi0505;
  assign n7818 = ~n7816 & n7817;
  assign n7819 = ~pi0239 ^ ~pi0497;
  assign n7820 = pi0240 ^ ~pi0542;
  assign n7821 = n7819 & n7820;
  assign n7822 = n7818 & n7821;
  assign n7823 = n7815 & n7822;
  assign n7824 = n7808 & n7823;
  assign n7825 = ~n7792 & ~n7824;
  assign n7826 = n7825 & pi0237;
  assign n7827 = pi0248 & ~pi0554;
  assign n7828 = ~pi0247 & pi0552;
  assign n7829 = ~n7827 & ~n7828;
  assign n7830 = ~pi0240 & pi0551;
  assign n7831 = pi0242 ^ ~pi0489;
  assign n7832 = ~n7830 & n7831;
  assign n7833 = n7829 & n7832;
  assign n7834 = pi0244 ^ ~pi0486;
  assign n7835 = n7834 & ~pi0233;
  assign n7836 = n7833 & n7835;
  assign n7837 = pi0240 & ~pi0551;
  assign n7838 = ~pi0248 & pi0554;
  assign n7839 = ~n7837 & ~n7838;
  assign n7840 = pi0247 & ~pi0552;
  assign n7841 = n7839 & ~n7840;
  assign n7842 = n7836 & n7841;
  assign n7843 = ~pi0238 ^ ~pi0577;
  assign n7844 = pi0246 ^ ~pi0563;
  assign n7845 = ~n7843 & n7844;
  assign n7846 = ~pi0245 ^ ~pi0580;
  assign n7847 = pi0234 ^ ~pi0485;
  assign n7848 = ~n7846 & n7847;
  assign n7849 = n7845 & n7848;
  assign n7850 = ~pi0235 ^ ~pi0549;
  assign n7851 = pi0249 ^ ~pi0555;
  assign n7852 = ~n7850 & n7851;
  assign n7853 = pi0239 ^ ~pi0550;
  assign n7854 = pi0241 ^ ~pi0553;
  assign n7855 = ~n7853 & n7854;
  assign n7856 = n7852 & n7855;
  assign n7857 = n7849 & n7856;
  assign n7858 = n7842 & n7857;
  assign n7859 = ~pi0241 & pi0490;
  assign n7860 = ~n7859 & pi0233;
  assign n7861 = pi0247 ^ ~pi0547;
  assign n7862 = n7860 & n7861;
  assign n7863 = pi0242 ^ ~pi0483;
  assign n7864 = pi0245 ^ ~pi0545;
  assign n7865 = n7863 & n7864;
  assign n7866 = n7862 & n7865;
  assign n7867 = pi0241 & ~pi0490;
  assign n7868 = pi0238 ^ ~pi0491;
  assign n7869 = ~n7867 & n7868;
  assign n7870 = n7866 & n7869;
  assign n7871 = ~pi0246 ^ ~pi0546;
  assign n7872 = pi0249 ^ ~pi0484;
  assign n7873 = ~n7871 & n7872;
  assign n7874 = pi0248 ^ ~pi0548;
  assign n7875 = pi0244 ^ ~pi0493;
  assign n7876 = n7874 & n7875;
  assign n7877 = n7873 & n7876;
  assign n7878 = ~pi0234 ^ ~pi0544;
  assign n7879 = pi0240 ^ ~pi0492;
  assign n7880 = ~n7878 & n7879;
  assign n7881 = ~pi0239 ^ ~pi0494;
  assign n7882 = pi0235 ^ ~pi0495;
  assign n7883 = n7881 & n7882;
  assign n7884 = n7880 & n7883;
  assign n7885 = n7877 & n7884;
  assign n7886 = n7870 & n7885;
  assign n7887 = ~n7858 & ~n7886;
  assign n7888 = n7887 & ~pi0237;
  assign n7889 = ~n7826 & ~n7888;
  assign n7890 = n7889 & ~n5882;
  assign n7891 = ~pi0245 & pi0514;
  assign n7892 = pi0249 ^ ~pi0579;
  assign n7893 = ~n7891 & n7892;
  assign n7894 = n7893 & pi0233;
  assign n7895 = pi0247 ^ ~pi0516;
  assign n7896 = pi0241 ^ ~pi0559;
  assign n7897 = n7895 & n7896;
  assign n7898 = n7894 & n7897;
  assign n7899 = pi0245 & ~pi0514;
  assign n7900 = pi0248 ^ ~pi0481;
  assign n7901 = ~n7899 & n7900;
  assign n7902 = n7898 & n7901;
  assign n7903 = ~pi0244 ^ ~pi0513;
  assign n7904 = pi0234 ^ ~pi0511;
  assign n7905 = ~n7903 & n7904;
  assign n7906 = pi0242 ^ ~pi0510;
  assign n7907 = pi0240 ^ ~pi0515;
  assign n7908 = n7906 & n7907;
  assign n7909 = n7905 & n7908;
  assign n7910 = pi0239 ^ ~pi0488;
  assign n7911 = ~pi0235 ^ ~pi0512;
  assign n7912 = ~n7910 & ~n7911;
  assign n7913 = pi0238 ^ ~pi0517;
  assign n7914 = pi0246 ^ ~pi0487;
  assign n7915 = n7913 & n7914;
  assign n7916 = n7912 & n7915;
  assign n7917 = n7909 & n7916;
  assign n7918 = n7902 & n7917;
  assign n7919 = ~n7918 & pi0237;
  assign n7920 = ~pi0248 & pi0521;
  assign n7921 = ~n7920 & ~pi0233;
  assign n7922 = ~pi0241 ^ ~pi0574;
  assign n7923 = n7921 & ~n7922;
  assign n7924 = pi0238 ^ ~pi0522;
  assign n7925 = pi0249 ^ ~pi0578;
  assign n7926 = n7924 & n7925;
  assign n7927 = n7923 & n7926;
  assign n7928 = pi0248 & ~pi0521;
  assign n7929 = pi0244 ^ ~pi0585;
  assign n7930 = ~n7928 & n7929;
  assign n7931 = n7927 & n7930;
  assign n7932 = ~pi0245 ^ ~pi0584;
  assign n7933 = ~pi0239 ^ ~pi0519;
  assign n7934 = ~n7932 & n7933;
  assign n7935 = ~pi0246 ^ ~pi0520;
  assign n7936 = pi0234 ^ ~pi0518;
  assign n7937 = ~n7935 & n7936;
  assign n7938 = n7934 & n7937;
  assign n7939 = ~pi0242 ^ ~pi0586;
  assign n7940 = pi0247 ^ ~pi0561;
  assign n7941 = ~n7939 & n7940;
  assign n7942 = pi0240 ^ ~pi0582;
  assign n7943 = pi0235 ^ ~pi0581;
  assign n7944 = n7942 & n7943;
  assign n7945 = n7941 & n7944;
  assign n7946 = n7938 & n7945;
  assign n7947 = n7931 & n7946;
  assign n7948 = n7919 & ~n7947;
  assign n7949 = ~n7948 & n5855;
  assign n7950 = ~pi0239 ^ ~pi0524;
  assign n7951 = pi0245 ^ ~pi0525;
  assign n7952 = n7950 & n7951;
  assign n7953 = ~pi0238 ^ ~pi0529;
  assign n7954 = pi0249 ^ ~pi0528;
  assign n7955 = ~n7953 & n7954;
  assign n7956 = n7952 & n7955;
  assign n7957 = ~pi0235 ^ ~pi0575;
  assign n7958 = pi0246 ^ ~pi0526;
  assign n7959 = ~n7957 & n7958;
  assign n7960 = pi0234 ^ ~pi0523;
  assign n7961 = pi0242 ^ ~pi0573;
  assign n7962 = n7960 & n7961;
  assign n7963 = n7959 & n7962;
  assign n7964 = n7956 & n7963;
  assign n7965 = ~pi0244 & pi0572;
  assign n7966 = ~pi0247 & pi0527;
  assign n7967 = ~n7965 & ~n7966;
  assign n7968 = pi0248 ^ ~pi0576;
  assign n7969 = n7967 & n7968;
  assign n7970 = pi0247 & ~pi0527;
  assign n7971 = ~n7970 & pi0233;
  assign n7972 = ~pi0241 ^ ~pi0571;
  assign n7973 = n7971 & ~n7972;
  assign n7974 = n7969 & n7973;
  assign n7975 = n7964 & n7974;
  assign n7976 = pi0244 & ~pi0572;
  assign n7977 = pi0240 ^ ~pi0530;
  assign n7978 = ~n7976 & n7977;
  assign n7979 = n7975 & n7978;
  assign n7980 = ~pi0248 ^ ~pi0565;
  assign n7981 = pi0234 ^ ~pi0570;
  assign n7982 = ~n7980 & n7981;
  assign n7983 = ~pi0246 ^ ~pi0564;
  assign n7984 = pi0240 ^ ~pi0560;
  assign n7985 = ~n7983 & n7984;
  assign n7986 = n7982 & n7985;
  assign n7987 = ~pi0245 ^ ~pi0568;
  assign n7988 = pi0247 ^ ~pi0532;
  assign n7989 = ~n7987 & n7988;
  assign n7990 = ~pi0239 ^ ~pi0569;
  assign n7991 = pi0238 ^ ~pi0498;
  assign n7992 = n7990 & n7991;
  assign n7993 = n7989 & n7992;
  assign n7994 = n7986 & n7993;
  assign n7995 = ~pi0249 & pi0482;
  assign n7996 = ~n7995 & ~pi0233;
  assign n7997 = pi0241 ^ ~pi0562;
  assign n7998 = n7996 & n7997;
  assign n7999 = pi0235 ^ ~pi0531;
  assign n8000 = ~pi0244 ^ ~pi0566;
  assign n8001 = n7999 & ~n8000;
  assign n8002 = n7998 & n8001;
  assign n8003 = n7994 & n8002;
  assign n8004 = pi0242 ^ ~pi0556;
  assign n8005 = pi0249 & ~pi0482;
  assign n8006 = n8004 & ~n8005;
  assign n8007 = n8003 & n8006;
  assign n8008 = ~n7979 & ~n8007;
  assign n8009 = n8008 & ~pi0237;
  assign n8010 = n7949 & ~n8009;
  assign po0750 = n7890 | n8010;
  assign n8012 = ~pi0806 & pi0990;
  assign n8013 = n8012 & pi0600;
  assign n8014 = ~n8013 ^ ~pi0594;
  assign po0751 = n8014 & ~pi0332;
  assign n8016 = pi0605 & ~pi0806;
  assign n8017 = n7308 & n8016;
  assign n8018 = n8017 ^ ~pi0595;
  assign po0752 = ~n8018 & ~pi0332;
  assign n8020 = n7306 & n8012;
  assign n8021 = pi0595 & pi0597;
  assign n8022 = n8020 & n8021;
  assign n8023 = n8022 ^ ~pi0596;
  assign po0753 = ~n8023 & ~pi0332;
  assign n8025 = ~n8020 ^ ~pi0597;
  assign po0754 = n8025 & ~pi0332;
  assign n8027 = ~po1038 & ~pi0882;
  assign n8028 = n8027 & pi0947;
  assign n8029 = ~n8028 & pi0598;
  assign n8030 = pi0740 & pi0780;
  assign n8031 = n3393 & n8030;
  assign po0755 = n8029 | n8031;
  assign n8033 = n8022 & pi0596;
  assign n8034 = ~n8033 ^ ~pi0599;
  assign po0756 = n8034 & ~pi0332;
  assign n8036 = n8012 ^ ~pi0600;
  assign po0757 = ~n8036 & ~pi0332;
  assign n8038 = ~pi0601 & pi0806;
  assign n8039 = ~n8038 & ~pi0332;
  assign n8040 = ~pi0806 & ~pi0989;
  assign po0758 = n8039 & ~n8040;
  assign n8042 = n5452 & pi0230;
  assign n8043 = ~pi0230 & pi0602;
  assign po0759 = n8042 | n8043;
  assign n8045 = pi0832 & ~pi0980;
  assign n8046 = n8045 & pi1060;
  assign n8047 = pi1038 & ~pi1061;
  assign n8048 = n8046 & n8047;
  assign po0897 = n8048 & pi0952;
  assign n8050 = ~po0897 & pi0603;
  assign n8051 = ~n8050 & ~pi0966;
  assign n8052 = po0897 & pi1100;
  assign n8053 = n8051 & ~n8052;
  assign n8054 = ~pi0871 & pi0966;
  assign n8055 = n8054 & ~pi0872;
  assign po0760 = ~n8053 & ~n8055;
  assign n8057 = n3395 & pi0823;
  assign n8058 = n8057 & ~pi0779;
  assign n8059 = ~pi0299 & pi0983;
  assign n8060 = n8059 & pi0907;
  assign n8061 = ~n8060 & pi0604;
  assign n8062 = ~n8057 & n8061;
  assign po0761 = n8058 | n8062;
  assign n8064 = pi0605 ^ ~pi0806;
  assign po0762 = n8064 & ~pi0332;
  assign n8066 = ~po0897 & ~pi0606;
  assign n8067 = ~n8066 & ~pi0966;
  assign n8068 = po0897 & ~pi1104;
  assign n8069 = n8067 & ~n8068;
  assign n8070 = pi0837 & pi0966;
  assign po0763 = n8069 | n8070;
  assign n8072 = po0897 & ~pi1107;
  assign n8073 = ~n8072 & ~pi0966;
  assign n8074 = ~po0897 & ~pi0607;
  assign po0764 = n8073 & ~n8074;
  assign n8076 = po0897 & ~pi1116;
  assign n8077 = ~n8076 & ~pi0966;
  assign n8078 = ~po0897 & ~pi0608;
  assign po0765 = n8077 & ~n8078;
  assign n8080 = po0897 & ~pi1118;
  assign n8081 = ~n8080 & ~pi0966;
  assign n8082 = ~po0897 & ~pi0609;
  assign po0766 = n8081 & ~n8082;
  assign n8084 = po0897 & ~pi1113;
  assign n8085 = ~n8084 & ~pi0966;
  assign n8086 = ~po0897 & ~pi0610;
  assign po0767 = n8085 & ~n8086;
  assign n8088 = po0897 & ~pi1114;
  assign n8089 = ~n8088 & ~pi0966;
  assign n8090 = ~po0897 & ~pi0611;
  assign po0768 = n8089 & ~n8090;
  assign n8092 = po0897 & ~pi1111;
  assign n8093 = ~n8092 & ~pi0966;
  assign n8094 = ~po0897 & ~pi0612;
  assign po0769 = n8093 & ~n8094;
  assign n8096 = po0897 & ~pi1115;
  assign n8097 = ~n8096 & ~pi0966;
  assign n8098 = ~po0897 & ~pi0613;
  assign po0770 = n8097 & ~n8098;
  assign n8100 = ~po0897 & pi0614;
  assign n8101 = po0897 & pi1102;
  assign n8102 = ~n8100 & ~n8101;
  assign n8103 = n8102 & ~pi0966;
  assign po0771 = ~n8103 & ~n8054;
  assign n8105 = n8027 & pi0907;
  assign n8106 = ~n8105 & ~pi0615;
  assign n8107 = pi0779 & pi0797;
  assign n8108 = n3396 & n8107;
  assign po0772 = n8106 | n8108;
  assign n8110 = ~po0897 & ~pi0616;
  assign n8111 = ~n8110 & ~pi0966;
  assign n8112 = po0897 & ~pi1101;
  assign n8113 = n8111 & ~n8112;
  assign n8114 = pi0872 & pi0966;
  assign po0773 = n8113 | n8114;
  assign n8116 = ~po0897 & ~pi0617;
  assign n8117 = ~n8116 & ~pi0966;
  assign n8118 = po0897 & ~pi1105;
  assign n8119 = n8117 & ~n8118;
  assign n8120 = pi0850 & pi0966;
  assign po0774 = n8119 | n8120;
  assign n8122 = po0897 & ~pi1117;
  assign n8123 = ~n8122 & ~pi0966;
  assign n8124 = ~po0897 & ~pi0618;
  assign po0775 = n8123 & ~n8124;
  assign n8126 = po0897 & ~pi1122;
  assign n8127 = ~n8126 & ~pi0966;
  assign n8128 = ~po0897 & ~pi0619;
  assign po0776 = n8127 & ~n8128;
  assign n8130 = po0897 & ~pi1112;
  assign n8131 = ~n8130 & ~pi0966;
  assign n8132 = ~po0897 & ~pi0620;
  assign po0777 = n8131 & ~n8132;
  assign n8134 = po0897 & ~pi1108;
  assign n8135 = ~n8134 & ~pi0966;
  assign n8136 = ~po0897 & ~pi0621;
  assign po0778 = n8135 & ~n8136;
  assign n8138 = po0897 & ~pi1109;
  assign n8139 = ~n8138 & ~pi0966;
  assign n8140 = ~po0897 & ~pi0622;
  assign po0779 = n8139 & ~n8140;
  assign n8142 = po0897 & ~pi1106;
  assign n8143 = ~n8142 & ~pi0966;
  assign n8144 = ~po0897 & ~pi0623;
  assign po0780 = n8143 & ~n8144;
  assign n8146 = n3392 & pi0831;
  assign n8147 = n8146 & ~pi0780;
  assign n8148 = n8059 & pi0947;
  assign n8149 = ~n8148 & pi0624;
  assign n8150 = ~n8146 & n8149;
  assign po0781 = n8147 | n8150;
  assign n8152 = pi1066 & pi1088;
  assign n8153 = ~pi0973 & ~pi1054;
  assign n8154 = n8152 & n8153;
  assign n8155 = n8154 & pi0832;
  assign po0954 = n8155 & ~pi0953;
  assign n8157 = po0954 & ~pi1116;
  assign n8158 = ~n8157 & ~pi0962;
  assign n8159 = ~po0954 & ~pi0625;
  assign po0782 = n8158 & ~n8159;
  assign n8161 = po0897 & ~pi1121;
  assign n8162 = ~n8161 & ~pi0966;
  assign n8163 = ~po0897 & ~pi0626;
  assign po0783 = n8162 & ~n8163;
  assign n8165 = po0954 & ~pi1117;
  assign n8166 = ~n8165 & ~pi0962;
  assign n8167 = ~po0954 & ~pi0627;
  assign po0784 = n8166 & ~n8167;
  assign n8169 = po0954 & ~pi1119;
  assign n8170 = ~n8169 & ~pi0962;
  assign n8171 = ~po0954 & ~pi0628;
  assign po0785 = n8170 & ~n8171;
  assign n8173 = po0897 & ~pi1119;
  assign n8174 = ~n8173 & ~pi0966;
  assign n8175 = ~po0897 & ~pi0629;
  assign po0786 = n8174 & ~n8175;
  assign n8177 = po0897 & ~pi1120;
  assign n8178 = ~n8177 & ~pi0966;
  assign n8179 = ~po0897 & ~pi0630;
  assign po0787 = n8178 & ~n8179;
  assign n8181 = po0954 & ~pi1113;
  assign n8182 = ~n8181 & ~pi0962;
  assign n8183 = ~po0954 & pi0631;
  assign po0788 = n8182 & ~n8183;
  assign n8185 = po0954 & ~pi1115;
  assign n8186 = ~n8185 & ~pi0962;
  assign n8187 = ~po0954 & pi0632;
  assign po0789 = n8186 & ~n8187;
  assign n8189 = po0897 & ~pi1110;
  assign n8190 = ~n8189 & ~pi0966;
  assign n8191 = ~po0897 & ~pi0633;
  assign po0790 = n8190 & ~n8191;
  assign n8193 = po0954 & ~pi1110;
  assign n8194 = ~n8193 & ~pi0962;
  assign n8195 = ~po0954 & ~pi0634;
  assign po0791 = n8194 & ~n8195;
  assign n8197 = po0954 & ~pi1112;
  assign n8198 = ~n8197 & ~pi0962;
  assign n8199 = ~po0954 & pi0635;
  assign po0792 = n8198 & ~n8199;
  assign n8201 = po0897 & ~pi1127;
  assign n8202 = ~n8201 & ~pi0966;
  assign n8203 = ~po0897 & ~pi0636;
  assign po0793 = n8202 & ~n8203;
  assign n8205 = po0954 & ~pi1105;
  assign n8206 = ~n8205 & ~pi0962;
  assign n8207 = ~po0954 & ~pi0637;
  assign po0794 = n8206 & ~n8207;
  assign n8209 = po0954 & ~pi1107;
  assign n8210 = ~n8209 & ~pi0962;
  assign n8211 = ~po0954 & ~pi0638;
  assign po0795 = n8210 & ~n8211;
  assign n8213 = po0954 & ~pi1109;
  assign n8214 = ~n8213 & ~pi0962;
  assign n8215 = ~po0954 & ~pi0639;
  assign po0796 = n8214 & ~n8215;
  assign n8217 = po0897 & ~pi1128;
  assign n8218 = ~n8217 & ~pi0966;
  assign n8219 = ~po0897 & ~pi0640;
  assign po0797 = n8218 & ~n8219;
  assign n8221 = po0954 & ~pi1121;
  assign n8222 = ~n8221 & ~pi0962;
  assign n8223 = ~po0954 & ~pi0641;
  assign po0798 = n8222 & ~n8223;
  assign n8225 = po0897 & ~pi1103;
  assign n8226 = ~n8225 & ~pi0966;
  assign n8227 = ~po0897 & ~pi0642;
  assign po0799 = n8226 & ~n8227;
  assign n8229 = po0954 & ~pi1104;
  assign n8230 = ~n8229 & ~pi0962;
  assign n8231 = ~po0954 & ~pi0643;
  assign po0800 = n8230 & ~n8231;
  assign n8233 = po0897 & ~pi1123;
  assign n8234 = ~n8233 & ~pi0966;
  assign n8235 = ~po0897 & ~pi0644;
  assign po0801 = n8234 & ~n8235;
  assign n8237 = po0897 & ~pi1125;
  assign n8238 = ~n8237 & ~pi0966;
  assign n8239 = ~po0897 & ~pi0645;
  assign po0802 = n8238 & ~n8239;
  assign n8241 = po0954 & ~pi1114;
  assign n8242 = ~n8241 & ~pi0962;
  assign n8243 = ~po0954 & pi0646;
  assign po0803 = n8242 & ~n8243;
  assign n8245 = po0954 & ~pi1120;
  assign n8246 = ~n8245 & ~pi0962;
  assign n8247 = ~po0954 & ~pi0647;
  assign po0804 = n8246 & ~n8247;
  assign n8249 = po0954 & ~pi1122;
  assign n8250 = ~n8249 & ~pi0962;
  assign n8251 = ~po0954 & ~pi0648;
  assign po0805 = n8250 & ~n8251;
  assign n8253 = po0954 & ~pi1126;
  assign n8254 = ~n8253 & ~pi0962;
  assign n8255 = ~po0954 & pi0649;
  assign po0806 = n8254 & ~n8255;
  assign n8257 = po0954 & ~pi1127;
  assign n8258 = ~n8257 & ~pi0962;
  assign n8259 = ~po0954 & pi0650;
  assign po0807 = n8258 & ~n8259;
  assign n8261 = po0897 & ~pi1130;
  assign n8262 = ~n8261 & ~pi0966;
  assign n8263 = ~po0897 & ~pi0651;
  assign po0808 = n8262 & ~n8263;
  assign n8265 = po0897 & ~pi1131;
  assign n8266 = ~n8265 & ~pi0966;
  assign n8267 = ~po0897 & ~pi0652;
  assign po0809 = n8266 & ~n8267;
  assign n8269 = po0897 & ~pi1129;
  assign n8270 = ~n8269 & ~pi0966;
  assign n8271 = ~po0897 & ~pi0653;
  assign po0810 = n8270 & ~n8271;
  assign n8273 = po0954 & ~pi1130;
  assign n8274 = ~n8273 & ~pi0962;
  assign n8275 = ~po0954 & pi0654;
  assign po0811 = n8274 & ~n8275;
  assign n8277 = po0954 & ~pi1124;
  assign n8278 = ~n8277 & ~pi0962;
  assign n8279 = ~po0954 & pi0655;
  assign po0812 = n8278 & ~n8279;
  assign n8281 = po0897 & ~pi1126;
  assign n8282 = ~n8281 & ~pi0966;
  assign n8283 = ~po0897 & ~pi0656;
  assign po0813 = n8282 & ~n8283;
  assign n8285 = po0954 & ~pi1131;
  assign n8286 = ~n8285 & ~pi0962;
  assign n8287 = ~po0954 & pi0657;
  assign po0814 = n8286 & ~n8287;
  assign n8289 = po0897 & ~pi1124;
  assign n8290 = ~n8289 & ~pi0966;
  assign n8291 = ~po0897 & ~pi0658;
  assign po0815 = n8290 & ~n8291;
  assign n8293 = pi0266 & pi0992;
  assign n8294 = n8293 & ~pi0280;
  assign n8295 = n8294 & ~pi0269;
  assign n8296 = ~pi0281 & ~pi0282;
  assign n8297 = n8295 & n8296;
  assign n8298 = ~pi0270 & ~pi0277;
  assign n8299 = n8298 & ~pi0264;
  assign n8300 = n8297 & n8299;
  assign n8301 = n8300 & ~pi0265;
  assign po0816 = n8301 ^ ~pi0274;
  assign n8303 = po0954 & ~pi1118;
  assign n8304 = ~n8303 & ~pi0962;
  assign n8305 = ~po0954 & ~pi0660;
  assign po0817 = n8304 & ~n8305;
  assign n8307 = po0954 & ~pi1101;
  assign n8308 = ~n8307 & ~pi0962;
  assign n8309 = ~po0954 & ~pi0661;
  assign po0818 = n8308 & ~n8309;
  assign n8311 = po0954 & ~pi1102;
  assign n8312 = ~n8311 & ~pi0962;
  assign n8313 = ~po0954 & ~pi0662;
  assign po0819 = n8312 & ~n8313;
  assign n8315 = pi0591 & ~pi0592;
  assign n8316 = n8315 & pi0334;
  assign n8317 = ~pi0591 & pi0592;
  assign n8318 = n8317 & pi0365;
  assign n8319 = ~n8316 & ~n8318;
  assign n8320 = ~n8319 & n4732;
  assign n8321 = n3823 & pi0588;
  assign n8322 = n8321 & pi0464;
  assign n8323 = ~n8320 & ~n8322;
  assign n8324 = n8323 & n2712;
  assign n8325 = ~n3823 & ~pi0588;
  assign n8326 = n8325 & n3819;
  assign n8327 = n8326 & pi0323;
  assign n8328 = n8324 & ~n8327;
  assign n8329 = ~pi0199 & pi0257;
  assign n8330 = pi0199 & pi1065;
  assign n8331 = ~n8329 & ~n8330;
  assign n8332 = n8331 & ~n2712;
  assign n8333 = ~n8332 & n3927;
  assign n8334 = ~n8328 & n8333;
  assign n8335 = ~pi0633 & pi1136;
  assign n8336 = ~pi0815 & ~pi1136;
  assign n8337 = ~n8335 & ~n8336;
  assign n8338 = n8337 & ~pi1134;
  assign n8339 = ~pi0766 & pi1136;
  assign n8340 = ~pi0855 & ~pi1136;
  assign n8341 = ~n8339 & ~n8340;
  assign n8342 = n8341 & pi1134;
  assign n8343 = ~n8338 & ~n8342;
  assign n8344 = n8343 & ~pi1135;
  assign n8345 = ~pi0634 & pi1136;
  assign n8346 = ~pi0784 & ~pi1136;
  assign n8347 = ~n8345 & ~n8346;
  assign n8348 = n8347 & ~pi1134;
  assign n8349 = pi1134 & pi1136;
  assign n8350 = n8349 & pi0700;
  assign n8351 = ~n8350 & pi1135;
  assign n8352 = ~n8348 & n8351;
  assign n8353 = ~pi1137 & ~pi1138;
  assign n8354 = ~n3927 & n8353;
  assign n8355 = ~n8352 & n8354;
  assign n8356 = ~n8344 & n8355;
  assign po0820 = n8334 | n8356;
  assign n8358 = n8315 & pi0404;
  assign n8359 = n8317 & pi0380;
  assign n8360 = ~n8358 & ~n8359;
  assign n8361 = ~n8360 & n4732;
  assign n8362 = n8321 & pi0429;
  assign n8363 = ~n8361 & ~n8362;
  assign n8364 = n8363 & n2712;
  assign n8365 = n8326 & pi0355;
  assign n8366 = n8364 & ~n8365;
  assign n8367 = ~pi0199 & pi0292;
  assign n8368 = pi0199 & pi1084;
  assign n8369 = ~n8367 & ~n8368;
  assign n8370 = n8369 & ~n2712;
  assign n8371 = ~n8370 & n3927;
  assign n8372 = ~n8366 & n8371;
  assign n8373 = pi0614 & pi1136;
  assign n8374 = pi0811 & ~pi1136;
  assign n8375 = ~n8373 & ~n8374;
  assign n8376 = n8375 & ~pi1134;
  assign n8377 = ~pi0772 & pi1136;
  assign n8378 = ~pi0872 & ~pi1136;
  assign n8379 = ~n8377 & ~n8378;
  assign n8380 = ~n8379 & pi1134;
  assign n8381 = ~n8376 & ~n8380;
  assign n8382 = ~n8381 & ~pi1135;
  assign n8383 = ~pi0662 & pi1136;
  assign n8384 = ~pi0785 & ~pi1136;
  assign n8385 = ~n8383 & ~n8384;
  assign n8386 = n8385 & ~pi1134;
  assign n8387 = n8349 & pi0727;
  assign n8388 = ~n8387 & pi1135;
  assign n8389 = ~n8386 & n8388;
  assign n8390 = ~n8389 & n8354;
  assign n8391 = ~n8382 & n8390;
  assign po0821 = n8372 | n8391;
  assign n8393 = po0954 & ~pi1108;
  assign n8394 = ~n8393 & ~pi0962;
  assign n8395 = ~po0954 & ~pi0665;
  assign po0822 = n8394 & ~n8395;
  assign n8397 = n8315 & pi0456;
  assign n8398 = n8317 & pi0337;
  assign n8399 = ~n8397 & ~n8398;
  assign n8400 = ~n8399 & n4732;
  assign n8401 = n8321 & pi0443;
  assign n8402 = ~n8400 & ~n8401;
  assign n8403 = n8402 & n2712;
  assign n8404 = n8326 & pi0441;
  assign n8405 = n8403 & ~n8404;
  assign n8406 = ~pi0199 & pi0297;
  assign n8407 = pi0199 & pi1044;
  assign n8408 = ~n8406 & ~n8407;
  assign n8409 = n8408 & ~n2712;
  assign n8410 = ~n8409 & n3927;
  assign n8411 = ~n8405 & n8410;
  assign n8412 = ~pi0607 & pi1136;
  assign n8413 = pi0799 & ~pi1136;
  assign n8414 = ~n8412 & ~n8413;
  assign n8415 = n8414 & ~pi1134;
  assign n8416 = ~pi0764 & pi1136;
  assign n8417 = ~n8416 & pi1134;
  assign n8418 = ~pi0873 & ~pi1136;
  assign n8419 = n8417 & ~n8418;
  assign n8420 = ~n8415 & ~n8419;
  assign n8421 = n8420 & ~pi1135;
  assign n8422 = ~pi0638 & pi1136;
  assign n8423 = ~pi0790 & ~pi1136;
  assign n8424 = ~n8422 & ~n8423;
  assign n8425 = n8424 & ~pi1134;
  assign n8426 = n8349 & pi0691;
  assign n8427 = ~n8426 & pi1135;
  assign n8428 = ~n8425 & n8427;
  assign n8429 = ~n8428 & n8354;
  assign n8430 = ~n8421 & n8429;
  assign po0823 = n8411 | n8430;
  assign n8432 = n8326 & pi0458;
  assign n8433 = n8315 & pi0319;
  assign n8434 = n8317 & pi0338;
  assign n8435 = ~n8433 & ~n8434;
  assign n8436 = ~n8435 & n4732;
  assign n8437 = n8321 & pi0444;
  assign n8438 = ~n8436 & ~n8437;
  assign n8439 = ~n8432 & n8438;
  assign n8440 = n8439 & n2712;
  assign n8441 = ~pi0199 & pi0294;
  assign n8442 = pi0199 & pi1072;
  assign n8443 = ~n8441 & ~n8442;
  assign n8444 = n8443 & ~n2712;
  assign n8445 = ~n8444 & n3927;
  assign n8446 = ~n8440 & n8445;
  assign n8447 = ~pi0642 & pi1136;
  assign n8448 = pi0809 & ~pi1136;
  assign n8449 = ~n8447 & ~n8448;
  assign n8450 = n8449 & ~pi1134;
  assign n8451 = ~pi0763 & pi1136;
  assign n8452 = ~n8451 & pi1134;
  assign n8453 = ~pi0871 & ~pi1136;
  assign n8454 = n8452 & ~n8453;
  assign n8455 = ~n8450 & ~n8454;
  assign n8456 = n8455 & ~pi1135;
  assign n8457 = ~pi0681 & pi1136;
  assign n8458 = ~pi0792 & ~pi1136;
  assign n8459 = ~n8457 & ~n8458;
  assign n8460 = n8459 & ~pi1134;
  assign n8461 = n8349 & pi0699;
  assign n8462 = ~n8461 & pi1135;
  assign n8463 = ~n8460 & n8462;
  assign n8464 = ~n8463 & n8354;
  assign n8465 = ~n8456 & n8464;
  assign po0824 = n8446 | n8465;
  assign n8467 = n8326 & pi0342;
  assign n8468 = n8315 & pi0390;
  assign n8469 = n8317 & pi0363;
  assign n8470 = ~n8468 & ~n8469;
  assign n8471 = ~n8470 & n4732;
  assign n8472 = n8321 & pi0414;
  assign n8473 = ~n8471 & ~n8472;
  assign n8474 = ~n8467 & n8473;
  assign n8475 = n8474 & n2712;
  assign n8476 = ~pi0199 & pi0291;
  assign n8477 = pi0199 & pi1049;
  assign n8478 = ~n8476 & ~n8477;
  assign n8479 = n8478 & ~n2712;
  assign n8480 = ~n8479 & n3927;
  assign n8481 = ~n8475 & n8480;
  assign n8482 = ~pi0603 & pi1136;
  assign n8483 = ~pi0981 & ~pi1136;
  assign n8484 = ~n8482 & ~n8483;
  assign n8485 = n8484 & ~pi1134;
  assign n8486 = ~pi0759 & pi1136;
  assign n8487 = ~pi0837 & ~pi1136;
  assign n8488 = ~n8486 & ~n8487;
  assign n8489 = n8488 & pi1134;
  assign n8490 = ~n8485 & ~n8489;
  assign n8491 = n8490 & ~pi1135;
  assign n8492 = ~pi0680 & pi1136;
  assign n8493 = ~pi0778 & ~pi1136;
  assign n8494 = ~n8492 & ~n8493;
  assign n8495 = n8494 & ~pi1134;
  assign n8496 = n8349 & pi0696;
  assign n8497 = ~n8496 & pi1135;
  assign n8498 = ~n8495 & n8497;
  assign n8499 = ~n8498 & n8354;
  assign n8500 = ~n8491 & n8499;
  assign po0825 = n8481 | n8500;
  assign n8502 = po0954 & ~pi1125;
  assign n8503 = ~n8502 & ~pi0962;
  assign n8504 = ~po0954 & pi0669;
  assign po0826 = n8503 & ~n8504;
  assign n8506 = pi0723 & pi1135;
  assign n8507 = ~n8506 & pi1134;
  assign n8508 = pi0745 & ~pi1135;
  assign n8509 = n8507 & ~n8508;
  assign n8510 = ~pi0612 & ~pi1135;
  assign n8511 = ~n8510 & ~pi1134;
  assign n8512 = pi0695 & pi1135;
  assign n8513 = n8511 & ~n8512;
  assign n8514 = ~n8509 & ~n8513;
  assign n8515 = ~n8514 & pi1136;
  assign n8516 = ~pi1135 & ~pi1136;
  assign n8517 = n8516 & pi1134;
  assign n8518 = n8517 & pi0852;
  assign n8519 = ~n8515 & ~n8518;
  assign n8520 = ~n8519 & n8354;
  assign n8521 = n8321 & pi0415;
  assign n8522 = ~n8521 & n2712;
  assign n8523 = n3822 & pi0391;
  assign n8524 = pi0364 & ~pi0590;
  assign n8525 = n8524 & ~pi0591;
  assign n8526 = ~n8523 & ~n8525;
  assign n8527 = n3819 & pi0343;
  assign n8528 = n8526 & ~n8527;
  assign n8529 = ~n8528 & n8325;
  assign n8530 = n8522 & ~n8529;
  assign n8531 = ~pi0199 & pi0258;
  assign n8532 = pi0199 & pi1062;
  assign n8533 = ~n8531 & ~n8532;
  assign n8534 = n8533 & ~n2712;
  assign n8535 = ~n8534 & n3927;
  assign n8536 = ~n8530 & n8535;
  assign po0827 = n8520 | n8536;
  assign n8538 = n8315 & pi0333;
  assign n8539 = n8317 & pi0447;
  assign n8540 = ~n8538 & ~n8539;
  assign n8541 = ~n8540 & n4732;
  assign n8542 = n8321 & pi0453;
  assign n8543 = ~n8541 & ~n8542;
  assign n8544 = n8543 & n2712;
  assign n8545 = n8326 & pi0327;
  assign n8546 = n8544 & ~n8545;
  assign n8547 = ~pi0199 & pi0261;
  assign n8548 = pi0199 & pi1040;
  assign n8549 = ~n8547 & ~n8548;
  assign n8550 = n8549 & ~n2712;
  assign n8551 = ~n8550 & n3927;
  assign n8552 = ~n8546 & n8551;
  assign n8553 = pi0724 & pi1135;
  assign n8554 = ~n8553 & pi1134;
  assign n8555 = pi0741 & ~pi1135;
  assign n8556 = n8554 & ~n8555;
  assign n8557 = ~pi0611 & ~pi1135;
  assign n8558 = ~n8557 & ~pi1134;
  assign n8559 = pi0646 & pi1135;
  assign n8560 = n8558 & ~n8559;
  assign n8561 = ~n8556 & ~n8560;
  assign n8562 = ~n8561 & pi1136;
  assign n8563 = n8517 & pi0865;
  assign n8564 = ~n8562 & ~n8563;
  assign n8565 = ~n8564 & n8354;
  assign po0828 = n8552 | n8565;
  assign n8567 = n8326 & pi0320;
  assign n8568 = n8315 & pi0397;
  assign n8569 = n8317 & pi0372;
  assign n8570 = ~n8568 & ~n8569;
  assign n8571 = ~n8570 & n4732;
  assign n8572 = n8321 & pi0422;
  assign n8573 = ~n8571 & ~n8572;
  assign n8574 = ~n8567 & n8573;
  assign n8575 = n8574 & n2712;
  assign n8576 = ~pi0199 & pi0290;
  assign n8577 = pi0199 & pi1048;
  assign n8578 = ~n8576 & ~n8577;
  assign n8579 = n8578 & ~n2712;
  assign n8580 = ~n8579 & n3927;
  assign n8581 = ~n8575 & n8580;
  assign n8582 = pi0616 & pi1136;
  assign n8583 = pi0808 & ~pi1136;
  assign n8584 = ~n8582 & ~n8583;
  assign n8585 = n8584 & ~pi1134;
  assign n8586 = ~pi0758 & pi1136;
  assign n8587 = ~pi0850 & ~pi1136;
  assign n8588 = ~n8586 & ~n8587;
  assign n8589 = ~n8588 & pi1134;
  assign n8590 = ~n8585 & ~n8589;
  assign n8591 = ~n8590 & ~pi1135;
  assign n8592 = ~pi0661 & pi1136;
  assign n8593 = ~pi0781 & ~pi1136;
  assign n8594 = ~n8592 & ~n8593;
  assign n8595 = n8594 & ~pi1134;
  assign n8596 = n8349 & pi0736;
  assign n8597 = ~n8596 & pi1135;
  assign n8598 = ~n8595 & n8597;
  assign n8599 = ~n8598 & n8354;
  assign n8600 = ~n8591 & n8599;
  assign po0829 = n8581 | n8600;
  assign n8602 = n8315 & pi0411;
  assign n8603 = n8317 & pi0387;
  assign n8604 = ~n8602 & ~n8603;
  assign n8605 = ~n8604 & n4732;
  assign n8606 = n8321 & pi0435;
  assign n8607 = ~n8605 & ~n8606;
  assign n8608 = n8607 & n2712;
  assign n8609 = n8326 & pi0452;
  assign n8610 = n8608 & ~n8609;
  assign n8611 = ~pi0199 & pi0295;
  assign n8612 = pi0199 & pi1053;
  assign n8613 = ~n8611 & ~n8612;
  assign n8614 = n8613 & ~n2712;
  assign n8615 = ~n8614 & n3927;
  assign n8616 = ~n8610 & n8615;
  assign n8617 = pi0749 & pi1136;
  assign n8618 = pi0866 & ~pi1136;
  assign n8619 = ~n8617 & ~n8618;
  assign n8620 = n8619 & pi1134;
  assign n8621 = ~pi0617 & pi1136;
  assign n8622 = pi0814 & ~pi1136;
  assign n8623 = ~n8621 & ~n8622;
  assign n8624 = ~n8623 & ~pi1134;
  assign n8625 = ~n8620 & ~n8624;
  assign n8626 = ~n8625 & ~pi1135;
  assign n8627 = ~pi0637 & pi1136;
  assign n8628 = ~pi0788 & ~pi1136;
  assign n8629 = ~n8627 & ~n8628;
  assign n8630 = n8629 & ~pi1134;
  assign n8631 = n8349 & pi0706;
  assign n8632 = ~n8631 & pi1135;
  assign n8633 = ~n8630 & n8632;
  assign n8634 = ~n8633 & n8354;
  assign n8635 = ~n8626 & n8634;
  assign po0830 = n8616 | n8635;
  assign n8637 = n8326 & pi0362;
  assign n8638 = n8315 & pi0463;
  assign n8639 = n8317 & pi0336;
  assign n8640 = ~n8638 & ~n8639;
  assign n8641 = ~n8640 & n4732;
  assign n8642 = n8321 & pi0437;
  assign n8643 = ~n8641 & ~n8642;
  assign n8644 = ~n8637 & n8643;
  assign n8645 = n8644 & n2712;
  assign n8646 = ~pi0199 & pi0256;
  assign n8647 = pi0199 & pi1070;
  assign n8648 = ~n8646 & ~n8647;
  assign n8649 = n8648 & ~n2712;
  assign n8650 = ~n8649 & n3927;
  assign n8651 = ~n8645 & n8650;
  assign n8652 = pi0622 & pi1136;
  assign n8653 = pi0804 & ~pi1136;
  assign n8654 = ~n8652 & ~n8653;
  assign n8655 = n8654 & ~pi1134;
  assign n8656 = ~pi0743 & pi1136;
  assign n8657 = ~pi0859 & ~pi1136;
  assign n8658 = ~n8656 & ~n8657;
  assign n8659 = ~n8658 & pi1134;
  assign n8660 = ~n8655 & ~n8659;
  assign n8661 = ~n8660 & ~pi1135;
  assign n8662 = ~pi0639 & pi1136;
  assign n8663 = ~pi0783 & ~pi1136;
  assign n8664 = ~n8662 & ~n8663;
  assign n8665 = n8664 & ~pi1134;
  assign n8666 = n8349 & pi0735;
  assign n8667 = ~n8666 & pi1135;
  assign n8668 = ~n8665 & n8667;
  assign n8669 = ~n8668 & n8354;
  assign n8670 = ~n8661 & n8669;
  assign po0831 = n8651 | n8670;
  assign n8672 = n8315 & pi0412;
  assign n8673 = n8317 & pi0388;
  assign n8674 = ~n8672 & ~n8673;
  assign n8675 = ~n8674 & n4732;
  assign n8676 = n8321 & pi0436;
  assign n8677 = ~n8675 & ~n8676;
  assign n8678 = n8677 & n2712;
  assign n8679 = n8326 & pi0455;
  assign n8680 = n8678 & ~n8679;
  assign n8681 = ~pi0199 & pi0296;
  assign n8682 = pi0199 & pi1037;
  assign n8683 = ~n8681 & ~n8682;
  assign n8684 = n8683 & ~n2712;
  assign n8685 = ~n8684 & n3927;
  assign n8686 = ~n8680 & n8685;
  assign n8687 = ~pi0623 & pi1136;
  assign n8688 = pi0803 & ~pi1136;
  assign n8689 = ~n8687 & ~n8688;
  assign n8690 = n8689 & ~pi1134;
  assign n8691 = ~pi0748 & pi1136;
  assign n8692 = ~n8691 & pi1134;
  assign n8693 = ~pi0876 & ~pi1136;
  assign n8694 = n8692 & ~n8693;
  assign n8695 = ~n8690 & ~n8694;
  assign n8696 = n8695 & ~pi1135;
  assign n8697 = ~pi0710 & pi1136;
  assign n8698 = ~pi0789 & ~pi1136;
  assign n8699 = ~n8697 & ~n8698;
  assign n8700 = n8699 & ~pi1134;
  assign n8701 = n8349 & pi0730;
  assign n8702 = ~n8701 & pi1135;
  assign n8703 = ~n8700 & n8702;
  assign n8704 = ~n8703 & n8354;
  assign n8705 = ~n8696 & n8704;
  assign po0832 = n8686 | n8705;
  assign n8707 = n8326 & pi0361;
  assign n8708 = n8315 & pi0410;
  assign n8709 = n8317 & pi0386;
  assign n8710 = ~n8708 & ~n8709;
  assign n8711 = ~n8710 & n4732;
  assign n8712 = n8321 & pi0434;
  assign n8713 = ~n8711 & ~n8712;
  assign n8714 = ~n8707 & n8713;
  assign n8715 = n8714 & n2712;
  assign n8716 = ~pi0199 & pi0293;
  assign n8717 = pi0199 & pi1059;
  assign n8718 = ~n8716 & ~n8717;
  assign n8719 = n8718 & ~n2712;
  assign n8720 = ~n8719 & n3927;
  assign n8721 = ~n8715 & n8720;
  assign n8722 = pi0746 & pi1136;
  assign n8723 = pi0881 & ~pi1136;
  assign n8724 = ~n8722 & ~n8723;
  assign n8725 = n8724 & pi1134;
  assign n8726 = ~pi0606 & pi1136;
  assign n8727 = pi0812 & ~pi1136;
  assign n8728 = ~n8726 & ~n8727;
  assign n8729 = ~n8728 & ~pi1134;
  assign n8730 = ~n8725 & ~n8729;
  assign n8731 = ~n8730 & ~pi1135;
  assign n8732 = ~pi0643 & pi1136;
  assign n8733 = ~pi0787 & ~pi1136;
  assign n8734 = ~n8732 & ~n8733;
  assign n8735 = n8734 & ~pi1134;
  assign n8736 = n8349 & pi0729;
  assign n8737 = ~n8736 & pi1135;
  assign n8738 = ~n8735 & n8737;
  assign n8739 = ~n8738 & n8354;
  assign n8740 = ~n8731 & n8739;
  assign po0833 = n8721 | n8740;
  assign n8742 = n8326 & pi0344;
  assign n8743 = n8315 & pi0335;
  assign n8744 = n8317 & pi0366;
  assign n8745 = ~n8743 & ~n8744;
  assign n8746 = ~n8745 & n4732;
  assign n8747 = n8321 & pi0416;
  assign n8748 = ~n8746 & ~n8747;
  assign n8749 = ~n8742 & n8748;
  assign n8750 = n8749 & n2712;
  assign n8751 = ~pi0199 & pi0259;
  assign n8752 = pi0199 & pi1069;
  assign n8753 = ~n8751 & ~n8752;
  assign n8754 = n8753 & ~n2712;
  assign n8755 = ~n8754 & n3927;
  assign n8756 = ~n8750 & n8755;
  assign n8757 = pi0742 & ~pi1135;
  assign n8758 = pi0704 & pi1135;
  assign n8759 = ~n8757 & ~n8758;
  assign n8760 = ~n8759 & pi1134;
  assign n8761 = ~n8760 & pi1136;
  assign n8762 = ~pi0635 & pi1135;
  assign n8763 = pi0620 & ~pi1135;
  assign n8764 = ~n8762 & ~n8763;
  assign n8765 = n8764 & ~pi1134;
  assign n8766 = n8761 & ~n8765;
  assign n8767 = n8517 & pi0870;
  assign n8768 = ~n8766 & ~n8767;
  assign n8769 = ~n8768 & n8354;
  assign po0834 = n8756 | n8769;
  assign n8771 = pi0688 & pi1135;
  assign n8772 = ~n8771 & pi1134;
  assign n8773 = pi0760 & ~pi1135;
  assign n8774 = n8772 & ~n8773;
  assign n8775 = ~pi0613 & ~pi1135;
  assign n8776 = ~n8775 & ~pi1134;
  assign n8777 = pi0632 & pi1135;
  assign n8778 = n8776 & ~n8777;
  assign n8779 = ~n8774 & ~n8778;
  assign n8780 = ~n8779 & pi1136;
  assign n8781 = n8517 & pi0856;
  assign n8782 = ~n8780 & ~n8781;
  assign n8783 = ~n8782 & n8354;
  assign n8784 = n3822 & pi0393;
  assign n8785 = n3819 & pi0346;
  assign n8786 = ~n8784 & ~n8785;
  assign n8787 = pi0368 & ~pi0590;
  assign n8788 = n8787 & ~pi0591;
  assign n8789 = n8786 & ~n8788;
  assign n8790 = ~n8789 & n8325;
  assign n8791 = n8321 & pi0418;
  assign n8792 = ~n8791 & n2712;
  assign n8793 = ~n8790 & n8792;
  assign n8794 = ~pi0199 & pi0260;
  assign n8795 = pi0199 & pi1067;
  assign n8796 = ~n8794 & ~n8795;
  assign n8797 = n8796 & ~n2712;
  assign n8798 = ~n8797 & n3927;
  assign n8799 = ~n8793 & n8798;
  assign po0835 = n8783 | n8799;
  assign n8801 = n8315 & pi0413;
  assign n8802 = n8317 & pi0389;
  assign n8803 = ~n8801 & ~n8802;
  assign n8804 = ~n8803 & n4732;
  assign n8805 = n8321 & pi0438;
  assign n8806 = ~n8804 & ~n8805;
  assign n8807 = n8806 & n2712;
  assign n8808 = n8326 & pi0450;
  assign n8809 = n8807 & ~n8808;
  assign n8810 = ~pi0199 & pi0255;
  assign n8811 = pi0199 & pi1036;
  assign n8812 = ~n8810 & ~n8811;
  assign n8813 = n8812 & ~n2712;
  assign n8814 = ~n8813 & n3927;
  assign n8815 = ~n8809 & n8814;
  assign n8816 = pi0621 & pi1136;
  assign n8817 = pi0810 & ~pi1136;
  assign n8818 = ~n8816 & ~n8817;
  assign n8819 = n8818 & ~pi1134;
  assign n8820 = ~pi0739 & pi1136;
  assign n8821 = ~pi0874 & ~pi1136;
  assign n8822 = ~n8820 & ~n8821;
  assign n8823 = ~n8822 & pi1134;
  assign n8824 = ~n8819 & ~n8823;
  assign n8825 = ~n8824 & ~pi1135;
  assign n8826 = ~pi0665 & pi1136;
  assign n8827 = ~pi0791 & ~pi1136;
  assign n8828 = ~n8826 & ~n8827;
  assign n8829 = n8828 & ~pi1134;
  assign n8830 = n8349 & pi0690;
  assign n8831 = ~n8830 & pi1135;
  assign n8832 = ~n8829 & n8831;
  assign n8833 = ~n8832 & n8354;
  assign n8834 = ~n8825 & n8833;
  assign po0836 = n8815 | n8834;
  assign n8836 = po0954 & ~pi1100;
  assign n8837 = ~n8836 & ~pi0962;
  assign n8838 = ~po0954 & ~pi0680;
  assign po0837 = n8837 & ~n8838;
  assign n8840 = po0954 & ~pi1103;
  assign n8841 = ~n8840 & ~pi0962;
  assign n8842 = ~po0954 & ~pi0681;
  assign po0838 = n8841 & ~n8842;
  assign n8844 = n8315 & pi0392;
  assign n8845 = n8317 & pi0367;
  assign n8846 = ~n8844 & ~n8845;
  assign n8847 = ~n8846 & n4732;
  assign n8848 = n8321 & pi0417;
  assign n8849 = ~n8847 & ~n8848;
  assign n8850 = n8849 & n2712;
  assign n8851 = n8326 & pi0345;
  assign n8852 = n8850 & ~n8851;
  assign n8853 = ~pi0199 & pi0251;
  assign n8854 = pi0199 & pi1039;
  assign n8855 = ~n8853 & ~n8854;
  assign n8856 = n8855 & ~n2712;
  assign n8857 = ~n8856 & n3927;
  assign n8858 = ~n8852 & n8857;
  assign n8859 = pi0686 & pi1135;
  assign n8860 = ~n8859 & pi1134;
  assign n8861 = pi0757 & ~pi1135;
  assign n8862 = n8860 & ~n8861;
  assign n8863 = ~pi0610 & ~pi1135;
  assign n8864 = ~n8863 & ~pi1134;
  assign n8865 = pi0631 & pi1135;
  assign n8866 = n8864 & ~n8865;
  assign n8867 = ~n8862 & ~n8866;
  assign n8868 = ~n8867 & pi1136;
  assign n8869 = n8517 & pi0848;
  assign n8870 = ~n8868 & ~n8869;
  assign n8871 = ~n8870 & n8354;
  assign po0839 = n8858 | n8871;
  assign po0980 = n8155 & pi0953;
  assign n8874 = po0980 & ~pi1130;
  assign n8875 = ~n8874 & ~pi0962;
  assign n8876 = ~po0980 & pi0684;
  assign po0841 = n8875 & ~n8876;
  assign n8878 = n8315 & pi0406;
  assign n8879 = n8317 & pi0382;
  assign n8880 = ~n8878 & ~n8879;
  assign n8881 = ~n8880 & n4732;
  assign n8882 = n8321 & pi0430;
  assign n8883 = ~n8881 & ~n8882;
  assign n8884 = n8883 & n2712;
  assign n8885 = n8326 & pi0357;
  assign n8886 = n8884 & ~n8885;
  assign n8887 = ~n6505 & ~pi0199;
  assign n8888 = pi0199 & pi1076;
  assign n8889 = ~n2712 & ~n8888;
  assign n8890 = ~n8887 & n8889;
  assign n8891 = ~n8890 & n3927;
  assign n8892 = ~n8886 & n8891;
  assign n8893 = pi0728 & pi1135;
  assign n8894 = ~n8893 & pi1134;
  assign n8895 = pi0744 & ~pi1135;
  assign n8896 = n8894 & ~n8895;
  assign n8897 = ~pi0652 & ~pi1135;
  assign n8898 = ~n8897 & ~pi1134;
  assign n8899 = pi0657 & pi1135;
  assign n8900 = n8898 & ~n8899;
  assign n8901 = ~n8896 & ~n8900;
  assign n8902 = ~n8901 & pi1136;
  assign n8903 = ~pi0813 & ~pi1134;
  assign n8904 = n8516 & ~n8903;
  assign n8905 = ~pi0860 & pi1134;
  assign n8906 = n8904 & ~n8905;
  assign n8907 = ~n8902 & ~n8906;
  assign n8908 = ~n8907 & n8354;
  assign po0842 = n8892 | n8908;
  assign n8910 = po0980 & ~pi1113;
  assign n8911 = ~n8910 & ~pi0962;
  assign n8912 = ~po0980 & pi0686;
  assign po0843 = n8911 & ~n8912;
  assign n8914 = po0980 & ~pi1127;
  assign n8915 = ~n8914 & ~pi0962;
  assign n8916 = ~po0980 & ~pi0687;
  assign po0844 = n8915 & ~n8916;
  assign n8918 = po0980 & ~pi1115;
  assign n8919 = ~n8918 & ~pi0962;
  assign n8920 = ~po0980 & pi0688;
  assign po0845 = n8919 & ~n8920;
  assign n8922 = n8326 & pi0351;
  assign n8923 = n8315 & pi0401;
  assign n8924 = n8317 & pi0376;
  assign n8925 = ~n8923 & ~n8924;
  assign n8926 = ~n8925 & n4732;
  assign n8927 = n8321 & pi0426;
  assign n8928 = ~n8926 & ~n8927;
  assign n8929 = ~n8922 & n8928;
  assign n8930 = n8929 & n2712;
  assign n8931 = ~n6475 & ~pi0199;
  assign n8932 = pi0199 & pi1079;
  assign n8933 = ~n2712 & ~n8932;
  assign n8934 = ~n8931 & n8933;
  assign n8935 = ~n8934 & n3927;
  assign n8936 = ~n8930 & n8935;
  assign n8937 = ~pi0703 & pi1135;
  assign n8938 = pi0752 & ~pi1135;
  assign n8939 = ~n8937 & ~n8938;
  assign n8940 = n8939 & pi1134;
  assign n8941 = ~pi0658 & ~pi1135;
  assign n8942 = pi0655 & pi1135;
  assign n8943 = ~n8941 & ~n8942;
  assign n8944 = n8943 & ~pi1134;
  assign n8945 = ~n8940 & ~n8944;
  assign n8946 = ~n8945 & pi1136;
  assign n8947 = ~pi0798 & ~pi1134;
  assign n8948 = n8516 & ~n8947;
  assign n8949 = ~pi0843 & pi1134;
  assign n8950 = n8948 & ~n8949;
  assign n8951 = ~n8946 & ~n8950;
  assign n8952 = ~n8951 & n8354;
  assign po0846 = n8936 | n8952;
  assign n8954 = po0980 & ~pi1108;
  assign n8955 = ~n8954 & ~pi0962;
  assign n8956 = ~po0980 & ~pi0690;
  assign po0847 = n8955 & ~n8956;
  assign n8958 = po0980 & ~pi1107;
  assign n8959 = ~n8958 & ~pi0962;
  assign n8960 = ~po0980 & ~pi0691;
  assign po0848 = n8959 & ~n8960;
  assign n8962 = n8315 & pi0402;
  assign n8963 = n8317 & pi0317;
  assign n8964 = ~n8962 & ~n8963;
  assign n8965 = ~n8964 & n4732;
  assign n8966 = n8321 & pi0427;
  assign n8967 = ~n8965 & ~n8966;
  assign n8968 = n8967 & n2712;
  assign n8969 = n8326 & pi0352;
  assign n8970 = n8968 & ~n8969;
  assign n8971 = ~n6487 & ~pi0199;
  assign n8972 = pi0199 & pi1078;
  assign n8973 = ~n2712 & ~n8972;
  assign n8974 = ~n8971 & n8973;
  assign n8975 = ~n8974 & n3927;
  assign n8976 = ~n8970 & n8975;
  assign n8977 = ~pi0726 & pi1135;
  assign n8978 = pi0770 & ~pi1135;
  assign n8979 = ~n8977 & ~n8978;
  assign n8980 = n8979 & pi1134;
  assign n8981 = ~pi0656 & ~pi1135;
  assign n8982 = pi0649 & pi1135;
  assign n8983 = ~n8981 & ~n8982;
  assign n8984 = n8983 & ~pi1134;
  assign n8985 = ~n8980 & ~n8984;
  assign n8986 = ~n8985 & pi1136;
  assign n8987 = ~pi0801 & ~pi1134;
  assign n8988 = n8516 & ~n8987;
  assign n8989 = ~pi0844 & pi1134;
  assign n8990 = n8988 & ~n8989;
  assign n8991 = ~n8986 & ~n8990;
  assign n8992 = ~n8991 & n8354;
  assign po0849 = n8976 | n8992;
  assign n8994 = po0954 & ~pi1129;
  assign n8995 = ~n8994 & ~pi0962;
  assign n8996 = ~po0954 & pi0693;
  assign po0850 = n8995 & ~n8996;
  assign n8998 = po0980 & ~pi1128;
  assign n8999 = ~n8998 & ~pi0962;
  assign n9000 = ~po0980 & pi0694;
  assign po0851 = n8999 & ~n9000;
  assign n9002 = po0954 & ~pi1111;
  assign n9003 = ~n9002 & ~pi0962;
  assign n9004 = ~po0954 & pi0695;
  assign po0852 = n9003 & ~n9004;
  assign n9006 = po0980 & ~pi1100;
  assign n9007 = ~n9006 & ~pi0962;
  assign n9008 = ~po0980 & ~pi0696;
  assign po0853 = n9007 & ~n9008;
  assign n9010 = po0980 & ~pi1129;
  assign n9011 = ~n9010 & ~pi0962;
  assign n9012 = ~po0980 & pi0697;
  assign po0854 = n9011 & ~n9012;
  assign n9014 = po0980 & ~pi1116;
  assign n9015 = ~n9014 & ~pi0962;
  assign n9016 = ~po0980 & pi0698;
  assign po0855 = n9015 & ~n9016;
  assign n9018 = po0980 & ~pi1103;
  assign n9019 = ~n9018 & ~pi0962;
  assign n9020 = ~po0980 & ~pi0699;
  assign po0856 = n9019 & ~n9020;
  assign n9022 = po0980 & ~pi1110;
  assign n9023 = ~n9022 & ~pi0962;
  assign n9024 = ~po0980 & ~pi0700;
  assign po0857 = n9023 & ~n9024;
  assign n9026 = po0980 & ~pi1123;
  assign n9027 = ~n9026 & ~pi0962;
  assign n9028 = ~po0980 & pi0701;
  assign po0858 = n9027 & ~n9028;
  assign n9030 = po0980 & ~pi1117;
  assign n9031 = ~n9030 & ~pi0962;
  assign n9032 = ~po0980 & pi0702;
  assign po0859 = n9031 & ~n9032;
  assign n9034 = po0980 & ~pi1124;
  assign n9035 = ~n9034 & ~pi0962;
  assign n9036 = ~po0980 & ~pi0703;
  assign po0860 = n9035 & ~n9036;
  assign n9038 = po0980 & ~pi1112;
  assign n9039 = ~n9038 & ~pi0962;
  assign n9040 = ~po0980 & pi0704;
  assign po0861 = n9039 & ~n9040;
  assign n9042 = po0980 & ~pi1125;
  assign n9043 = ~n9042 & ~pi0962;
  assign n9044 = ~po0980 & ~pi0705;
  assign po0862 = n9043 & ~n9044;
  assign n9046 = po0980 & ~pi1105;
  assign n9047 = ~n9046 & ~pi0962;
  assign n9048 = ~po0980 & ~pi0706;
  assign po0863 = n9047 & ~n9048;
  assign n9050 = n8315 & pi0395;
  assign n9051 = n8317 & pi0370;
  assign n9052 = ~n9050 & ~n9051;
  assign n9053 = ~n9052 & n4732;
  assign n9054 = n8321 & pi0420;
  assign n9055 = ~n9053 & ~n9054;
  assign n9056 = n9055 & n2712;
  assign n9057 = n8326 & pi0347;
  assign n9058 = n9056 & ~n9057;
  assign n9059 = n4379 & ~pi0304;
  assign n9060 = pi0199 & ~pi1055;
  assign n9061 = ~n9059 & ~n9060;
  assign n9062 = n4471 & ~pi1048;
  assign n9063 = n9061 & ~n9062;
  assign n9064 = ~n9063 & ~n2712;
  assign n9065 = ~n9064 & n3927;
  assign n9066 = ~n9058 & n9065;
  assign n9067 = pi0753 & ~pi1135;
  assign n9068 = pi0702 & pi1135;
  assign n9069 = ~n9067 & ~n9068;
  assign n9070 = ~n9069 & pi1134;
  assign n9071 = ~n9070 & pi1136;
  assign n9072 = pi0627 & pi1135;
  assign n9073 = pi0618 & ~pi1135;
  assign n9074 = ~n9072 & ~n9073;
  assign n9075 = n9074 & ~pi1134;
  assign n9076 = n9071 & ~n9075;
  assign n9077 = n8517 & pi0847;
  assign n9078 = ~n9076 & ~n9077;
  assign n9079 = ~n9078 & n8354;
  assign po0864 = n9066 | n9079;
  assign n9081 = n8326 & pi0321;
  assign n9082 = n8315 & pi0328;
  assign n9083 = n8317 & pi0442;
  assign n9084 = ~n9082 & ~n9083;
  assign n9085 = ~n9084 & n4732;
  assign n9086 = n8321 & pi0459;
  assign n9087 = ~n9085 & ~n9086;
  assign n9088 = ~n9081 & n9087;
  assign n9089 = n9088 & n2712;
  assign n9090 = n4379 & ~pi0305;
  assign n9091 = pi0199 & ~pi1058;
  assign n9092 = ~n9090 & ~n9091;
  assign n9093 = n4471 & ~pi1084;
  assign n9094 = n9092 & ~n9093;
  assign n9095 = ~n9094 & ~n2712;
  assign n9096 = ~n9095 & n3927;
  assign n9097 = ~n9089 & n9096;
  assign n9098 = pi0754 & ~pi1135;
  assign n9099 = pi0709 & pi1135;
  assign n9100 = ~n9098 & ~n9099;
  assign n9101 = ~n9100 & pi1134;
  assign n9102 = ~n9101 & pi1136;
  assign n9103 = pi0660 & pi1135;
  assign n9104 = pi0609 & ~pi1135;
  assign n9105 = ~n9103 & ~n9104;
  assign n9106 = n9105 & ~pi1134;
  assign n9107 = n9102 & ~n9106;
  assign n9108 = n8517 & pi0857;
  assign n9109 = ~n9107 & ~n9108;
  assign n9110 = ~n9109 & n8354;
  assign po0865 = n9097 | n9110;
  assign n9112 = po0980 & ~pi1118;
  assign n9113 = ~n9112 & ~pi0962;
  assign n9114 = ~po0980 & pi0709;
  assign po0866 = n9113 & ~n9114;
  assign n9116 = po0954 & ~pi1106;
  assign n9117 = ~n9116 & ~pi0962;
  assign n9118 = ~po0954 & ~pi0710;
  assign po0867 = n9117 & ~n9118;
  assign n9120 = n8315 & pi0398;
  assign n9121 = n8317 & pi0373;
  assign n9122 = ~n9120 & ~n9121;
  assign n9123 = ~n9122 & n4732;
  assign n9124 = n8321 & pi0423;
  assign n9125 = ~n9123 & ~n9124;
  assign n9126 = n9125 & n2712;
  assign n9127 = n8326 & pi0348;
  assign n9128 = n9126 & ~n9127;
  assign n9129 = n4379 & ~pi0306;
  assign n9130 = pi0199 & ~pi1087;
  assign n9131 = ~n9129 & ~n9130;
  assign n9132 = n4471 & ~pi1059;
  assign n9133 = n9131 & ~n9132;
  assign n9134 = ~n9133 & ~n2712;
  assign n9135 = ~n9134 & n3927;
  assign n9136 = ~n9128 & n9135;
  assign n9137 = pi0755 & ~pi1135;
  assign n9138 = pi0725 & pi1135;
  assign n9139 = ~n9137 & ~n9138;
  assign n9140 = ~n9139 & pi1134;
  assign n9141 = ~n9140 & pi1136;
  assign n9142 = pi0647 & pi1135;
  assign n9143 = pi0630 & ~pi1135;
  assign n9144 = ~n9142 & ~n9143;
  assign n9145 = n9144 & ~pi1134;
  assign n9146 = n9141 & ~n9145;
  assign n9147 = n8517 & pi0858;
  assign n9148 = ~n9146 & ~n9147;
  assign n9149 = ~n9148 & n8354;
  assign po0868 = n9136 | n9149;
  assign n9151 = n8315 & pi0400;
  assign n9152 = n8317 & pi0374;
  assign n9153 = ~n9151 & ~n9152;
  assign n9154 = ~n9153 & n4732;
  assign n9155 = n8321 & pi0425;
  assign n9156 = ~n9154 & ~n9155;
  assign n9157 = n9156 & n2712;
  assign n9158 = n8326 & pi0350;
  assign n9159 = n9157 & ~n9158;
  assign n9160 = n4379 & ~pi0298;
  assign n9161 = pi0199 & ~pi1035;
  assign n9162 = ~n9160 & ~n9161;
  assign n9163 = n4471 & ~pi1044;
  assign n9164 = n9162 & ~n9163;
  assign n9165 = ~n9164 & ~n2712;
  assign n9166 = ~n9165 & n3927;
  assign n9167 = ~n9159 & n9166;
  assign n9168 = pi0751 & ~pi1135;
  assign n9169 = pi0701 & pi1135;
  assign n9170 = ~n9168 & ~n9169;
  assign n9171 = ~n9170 & pi1134;
  assign n9172 = ~n9171 & pi1136;
  assign n9173 = pi0715 & pi1135;
  assign n9174 = pi0644 & ~pi1135;
  assign n9175 = ~n9173 & ~n9174;
  assign n9176 = n9175 & ~pi1134;
  assign n9177 = n9172 & ~n9176;
  assign n9178 = n8517 & pi0842;
  assign n9179 = ~n9177 & ~n9178;
  assign n9180 = ~n9179 & n8354;
  assign po0869 = n9167 | n9180;
  assign n9182 = n8315 & pi0396;
  assign n9183 = n8317 & pi0371;
  assign n9184 = ~n9182 & ~n9183;
  assign n9185 = ~n9184 & n4732;
  assign n9186 = n8321 & pi0421;
  assign n9187 = ~n9185 & ~n9186;
  assign n9188 = n9187 & n2712;
  assign n9189 = n8326 & pi0322;
  assign n9190 = n9188 & ~n9189;
  assign n9191 = n4379 & ~pi0309;
  assign n9192 = pi0199 & ~pi1051;
  assign n9193 = ~n9191 & ~n9192;
  assign n9194 = n4471 & ~pi1072;
  assign n9195 = n9193 & ~n9194;
  assign n9196 = ~n9195 & ~n2712;
  assign n9197 = ~n9196 & n3927;
  assign n9198 = ~n9190 & n9197;
  assign n9199 = pi0756 & ~pi1135;
  assign n9200 = pi0734 & pi1135;
  assign n9201 = ~n9199 & ~n9200;
  assign n9202 = ~n9201 & pi1134;
  assign n9203 = ~n9202 & pi1136;
  assign n9204 = pi0628 & pi1135;
  assign n9205 = pi0629 & ~pi1135;
  assign n9206 = ~n9204 & ~n9205;
  assign n9207 = n9206 & ~pi1134;
  assign n9208 = n9203 & ~n9207;
  assign n9209 = n8517 & pi0854;
  assign n9210 = ~n9208 & ~n9209;
  assign n9211 = ~n9210 & n8354;
  assign po0870 = n9198 | n9211;
  assign n9213 = n8326 & pi0461;
  assign n9214 = n8315 & pi0326;
  assign n9215 = n8317 & pi0439;
  assign n9216 = ~n9214 & ~n9215;
  assign n9217 = ~n9216 & n4732;
  assign n9218 = n8321 & pi0449;
  assign n9219 = ~n9217 & ~n9218;
  assign n9220 = ~n9213 & n9219;
  assign n9221 = n9220 & n2712;
  assign n9222 = ~n6445 & ~pi0199;
  assign n9223 = pi0199 & pi1057;
  assign n9224 = ~n2712 & ~n9223;
  assign n9225 = ~n9222 & n9224;
  assign n9226 = ~n9225 & n3927;
  assign n9227 = ~n9221 & n9226;
  assign n9228 = pi0697 & pi1135;
  assign n9229 = ~n9228 & pi1134;
  assign n9230 = pi0762 & ~pi1135;
  assign n9231 = n9229 & ~n9230;
  assign n9232 = ~pi0653 & ~pi1135;
  assign n9233 = ~n9232 & ~pi1134;
  assign n9234 = pi0693 & pi1135;
  assign n9235 = n9233 & ~n9234;
  assign n9236 = ~n9231 & ~n9235;
  assign n9237 = ~n9236 & pi1136;
  assign n9238 = ~pi0816 & ~pi1134;
  assign n9239 = n8516 & ~n9238;
  assign n9240 = ~pi0867 & pi1134;
  assign n9241 = n9239 & ~n9240;
  assign n9242 = ~n9237 & ~n9241;
  assign n9243 = ~n9242 & n8354;
  assign po0871 = n9227 | n9243;
  assign n9245 = po0954 & ~pi1123;
  assign n9246 = ~n9245 & ~pi0962;
  assign n9247 = ~po0954 & ~pi0715;
  assign po0872 = n9246 & ~n9247;
  assign n9249 = n8326 & pi0349;
  assign n9250 = n8315 & pi0329;
  assign n9251 = n8317 & pi0440;
  assign n9252 = ~n9250 & ~n9251;
  assign n9253 = ~n9252 & n4732;
  assign n9254 = ~n9249 & ~n9253;
  assign n9255 = n8321 & pi0454;
  assign n9256 = ~n9255 & n2712;
  assign n9257 = n9254 & n9256;
  assign n9258 = n4471 & ~pi1053;
  assign n9259 = n4379 & ~pi0307;
  assign n9260 = ~n9258 & ~n9259;
  assign n9261 = pi0199 & ~pi1043;
  assign n9262 = n9260 & ~n9261;
  assign n9263 = ~n9262 & ~n2712;
  assign n9264 = ~n9263 & n3927;
  assign n9265 = ~n9257 & n9264;
  assign n9266 = pi0761 & ~pi1135;
  assign n9267 = pi0738 & pi1135;
  assign n9268 = ~n9266 & ~n9267;
  assign n9269 = ~n9268 & pi1134;
  assign n9270 = ~n9269 & pi1136;
  assign n9271 = pi0641 & pi1135;
  assign n9272 = pi0626 & ~pi1135;
  assign n9273 = ~n9271 & ~n9272;
  assign n9274 = n9273 & ~pi1134;
  assign n9275 = n9270 & ~n9274;
  assign n9276 = n8517 & pi0845;
  assign n9277 = ~n9275 & ~n9276;
  assign n9278 = ~n9277 & n8354;
  assign po0873 = n9265 | n9278;
  assign n9280 = n8326 & pi0462;
  assign n9281 = n8315 & pi0318;
  assign n9282 = n8317 & pi0377;
  assign n9283 = ~n9281 & ~n9282;
  assign n9284 = ~n9283 & n4732;
  assign n9285 = n8321 & pi0448;
  assign n9286 = ~n9284 & ~n9285;
  assign n9287 = ~n9280 & n9286;
  assign n9288 = n9287 & n2712;
  assign n9289 = ~n6481 & ~pi0199;
  assign n9290 = pi0199 & pi1074;
  assign n9291 = ~n2712 & ~n9290;
  assign n9292 = ~n9289 & n9291;
  assign n9293 = ~n9292 & n3927;
  assign n9294 = ~n9288 & n9293;
  assign n9295 = ~pi0705 & pi1135;
  assign n9296 = pi0768 & ~pi1135;
  assign n9297 = ~n9295 & ~n9296;
  assign n9298 = ~n9297 & pi1134;
  assign n9299 = ~n9298 & pi1136;
  assign n9300 = ~pi0669 & pi1135;
  assign n9301 = pi0645 & ~pi1135;
  assign n9302 = ~n9300 & ~n9301;
  assign n9303 = n9302 & ~pi1134;
  assign n9304 = n9299 & ~n9303;
  assign n9305 = ~pi0800 & ~pi1134;
  assign n9306 = n8516 & ~n9305;
  assign n9307 = ~pi0839 & pi1134;
  assign n9308 = n9306 & ~n9307;
  assign n9309 = ~n9304 & ~n9308;
  assign n9310 = ~n9309 & n8354;
  assign po0874 = n9294 | n9310;
  assign n9312 = n8326 & pi0315;
  assign n9313 = n8321 & pi0419;
  assign n9314 = ~n9312 & ~n9313;
  assign n9315 = n8315 & pi0394;
  assign n9316 = n8317 & pi0369;
  assign n9317 = ~n9315 & ~n9316;
  assign n9318 = ~n9317 & n4732;
  assign n9319 = ~n9318 & n2712;
  assign n9320 = n9314 & n9319;
  assign n9321 = n4379 & ~pi0303;
  assign n9322 = pi0199 & ~pi1080;
  assign n9323 = ~n9321 & ~n9322;
  assign n9324 = n4471 & ~pi1049;
  assign n9325 = n9323 & ~n9324;
  assign n9326 = ~n9325 & ~n2712;
  assign n9327 = ~n9326 & n3927;
  assign n9328 = ~n9320 & n9327;
  assign n9329 = pi0767 & ~pi1135;
  assign n9330 = pi0698 & pi1135;
  assign n9331 = ~n9329 & ~n9330;
  assign n9332 = ~n9331 & pi1134;
  assign n9333 = ~n9332 & pi1136;
  assign n9334 = pi0625 & pi1135;
  assign n9335 = pi0608 & ~pi1135;
  assign n9336 = ~n9334 & ~n9335;
  assign n9337 = n9336 & ~pi1134;
  assign n9338 = n9333 & ~n9337;
  assign n9339 = n8517 & pi0853;
  assign n9340 = ~n9338 & ~n9339;
  assign n9341 = ~n9340 & n8354;
  assign po0875 = n9328 | n9341;
  assign n9343 = n8326 & pi0353;
  assign n9344 = n8315 & pi0325;
  assign n9345 = n8317 & pi0378;
  assign n9346 = ~n9344 & ~n9345;
  assign n9347 = ~n9346 & n4732;
  assign n9348 = n8321 & pi0451;
  assign n9349 = ~n9347 & ~n9348;
  assign n9350 = ~n9343 & n9349;
  assign n9351 = n9350 & n2712;
  assign n9352 = ~n6493 & ~pi0199;
  assign n9353 = pi0199 & pi1063;
  assign n9354 = ~n2712 & ~n9353;
  assign n9355 = ~n9352 & n9354;
  assign n9356 = ~n9355 & n3927;
  assign n9357 = ~n9351 & n9356;
  assign n9358 = pi0774 & ~pi1135;
  assign n9359 = ~n9358 & pi1134;
  assign n9360 = ~pi0687 & pi1135;
  assign n9361 = n9359 & ~n9360;
  assign n9362 = ~pi0636 & ~pi1135;
  assign n9363 = ~n9362 & ~pi1134;
  assign n9364 = pi0650 & pi1135;
  assign n9365 = n9363 & ~n9364;
  assign n9366 = ~n9361 & ~n9365;
  assign n9367 = ~n9366 & pi1136;
  assign n9368 = ~pi0807 & ~pi1134;
  assign n9369 = n8516 & ~n9368;
  assign n9370 = ~pi0868 & pi1134;
  assign n9371 = n9369 & ~n9370;
  assign n9372 = ~n9367 & ~n9371;
  assign n9373 = ~n9372 & n8354;
  assign po0876 = n9357 | n9373;
  assign n9375 = n8326 & pi0356;
  assign n9376 = n8315 & pi0405;
  assign n9377 = n8317 & pi0381;
  assign n9378 = ~n9376 & ~n9377;
  assign n9379 = ~n9378 & n4732;
  assign n9380 = n8321 & pi0445;
  assign n9381 = ~n9379 & ~n9380;
  assign n9382 = ~n9375 & n9381;
  assign n9383 = n9382 & n2712;
  assign n9384 = ~n6511 & ~pi0199;
  assign n9385 = pi0199 & pi1081;
  assign n9386 = ~n2712 & ~n9385;
  assign n9387 = ~n9384 & n9386;
  assign n9388 = ~n9387 & n3927;
  assign n9389 = ~n9383 & n9388;
  assign n9390 = pi0684 & pi1135;
  assign n9391 = ~n9390 & pi1134;
  assign n9392 = pi0750 & ~pi1135;
  assign n9393 = n9391 & ~n9392;
  assign n9394 = ~pi0651 & ~pi1135;
  assign n9395 = ~n9394 & ~pi1134;
  assign n9396 = pi0654 & pi1135;
  assign n9397 = n9395 & ~n9396;
  assign n9398 = ~n9393 & ~n9397;
  assign n9399 = ~n9398 & pi1136;
  assign n9400 = ~pi0794 & ~pi1134;
  assign n9401 = n8516 & ~n9400;
  assign n9402 = ~pi0880 & pi1134;
  assign n9403 = n9401 & ~n9402;
  assign n9404 = ~n9399 & ~n9403;
  assign n9405 = ~n9404 & n8354;
  assign po0877 = n9389 | n9405;
  assign n9407 = pi0747 & pi0773;
  assign n9408 = pi0731 & ~pi0945;
  assign n9409 = n9407 & n9408;
  assign n9410 = pi0775 & pi0988;
  assign n9411 = n9409 & n9410;
  assign n9412 = n9411 & pi0769;
  assign n9413 = ~n9412 ^ ~pi0721;
  assign n9414 = pi0765 ^ ~pi0798;
  assign n9415 = pi0771 ^ ~pi0800;
  assign n9416 = n9414 & n9415;
  assign n9417 = pi0747 ^ ~pi0807;
  assign n9418 = ~pi0775 ^ ~pi0816;
  assign n9419 = n9417 & ~n9418;
  assign n9420 = n9416 & n9419;
  assign n9421 = pi0769 ^ ~pi0794;
  assign n9422 = pi0773 ^ ~pi0801;
  assign n9423 = n9421 & n9422;
  assign n9424 = pi0721 ^ ~pi0813;
  assign n9425 = ~pi0731 ^ ~pi0795;
  assign n9426 = n9424 & ~n9425;
  assign n9427 = n9423 & n9426;
  assign po0978 = n9420 & n9427;
  assign po0878 = n9413 & ~po0978;
  assign n9430 = n8315 & pi0403;
  assign n9431 = n8317 & pi0379;
  assign n9432 = ~n9430 & ~n9431;
  assign n9433 = ~n9432 & n4732;
  assign n9434 = n8321 & pi0428;
  assign n9435 = ~n9433 & ~n9434;
  assign n9436 = n9435 & n2712;
  assign n9437 = n8326 & pi0354;
  assign n9438 = n9436 & ~n9437;
  assign n9439 = ~n6499 & ~pi0199;
  assign n9440 = pi0199 & pi1045;
  assign n9441 = ~n2712 & ~n9440;
  assign n9442 = ~n9439 & n9441;
  assign n9443 = ~n9442 & n3927;
  assign n9444 = ~n9438 & n9443;
  assign n9445 = pi0694 & pi1135;
  assign n9446 = ~n9445 & pi1134;
  assign n9447 = pi0776 & ~pi1135;
  assign n9448 = n9446 & ~n9447;
  assign n9449 = ~pi0640 & ~pi1135;
  assign n9450 = ~n9449 & ~pi1134;
  assign n9451 = pi0732 & pi1135;
  assign n9452 = n9450 & ~n9451;
  assign n9453 = ~n9448 & ~n9452;
  assign n9454 = ~n9453 & pi1136;
  assign n9455 = ~pi0795 & ~pi1134;
  assign n9456 = n8516 & ~n9455;
  assign n9457 = ~pi0851 & pi1134;
  assign n9458 = n9456 & ~n9457;
  assign n9459 = ~n9454 & ~n9458;
  assign n9460 = ~n9459 & n8354;
  assign po0879 = n9444 | n9460;
  assign n9462 = po0980 & ~pi1111;
  assign n9463 = ~n9462 & ~pi0962;
  assign n9464 = ~po0980 & pi0723;
  assign po0880 = n9463 & ~n9464;
  assign n9466 = po0980 & ~pi1114;
  assign n9467 = ~n9466 & ~pi0962;
  assign n9468 = ~po0980 & pi0724;
  assign po0881 = n9467 & ~n9468;
  assign n9470 = po0980 & ~pi1120;
  assign n9471 = ~n9470 & ~pi0962;
  assign n9472 = ~po0980 & pi0725;
  assign po0882 = n9471 & ~n9472;
  assign n9474 = po0980 & ~pi1126;
  assign n9475 = ~n9474 & ~pi0962;
  assign n9476 = ~po0980 & ~pi0726;
  assign po0883 = n9475 & ~n9476;
  assign n9478 = po0980 & ~pi1102;
  assign n9479 = ~n9478 & ~pi0962;
  assign n9480 = ~po0980 & ~pi0727;
  assign po0884 = n9479 & ~n9480;
  assign n9482 = po0980 & ~pi1131;
  assign n9483 = ~n9482 & ~pi0962;
  assign n9484 = ~po0980 & pi0728;
  assign po0885 = n9483 & ~n9484;
  assign n9486 = po0980 & ~pi1104;
  assign n9487 = ~n9486 & ~pi0962;
  assign n9488 = ~po0980 & ~pi0729;
  assign po0886 = n9487 & ~n9488;
  assign n9490 = po0980 & ~pi1106;
  assign n9491 = ~n9490 & ~pi0962;
  assign n9492 = ~po0980 & ~pi0730;
  assign po0887 = n9491 & ~n9492;
  assign n9494 = ~pi0945 & pi0988;
  assign n9495 = n9407 & n9494;
  assign n9496 = ~n9495 ^ ~pi0731;
  assign po0888 = ~po0978 & n9496;
  assign n9498 = po0954 & ~pi1128;
  assign n9499 = ~n9498 & ~pi0962;
  assign n9500 = ~po0954 & pi0732;
  assign po0889 = n9499 & ~n9500;
  assign n9502 = n8326 & pi0316;
  assign n9503 = n8315 & pi0399;
  assign n9504 = n8317 & pi0375;
  assign n9505 = ~n9503 & ~n9504;
  assign n9506 = ~n9505 & n4732;
  assign n9507 = n8321 & pi0424;
  assign n9508 = ~n9506 & ~n9507;
  assign n9509 = ~n9502 & n9508;
  assign n9510 = n9509 & n2712;
  assign n9511 = n4379 & ~pi0308;
  assign n9512 = pi0199 & ~pi1047;
  assign n9513 = ~n9511 & ~n9512;
  assign n9514 = n4471 & ~pi1037;
  assign n9515 = n9513 & ~n9514;
  assign n9516 = ~n9515 & ~n2712;
  assign n9517 = ~n9516 & n3927;
  assign n9518 = ~n9510 & n9517;
  assign n9519 = pi0777 & ~pi1135;
  assign n9520 = pi0737 & pi1135;
  assign n9521 = ~n9519 & ~n9520;
  assign n9522 = ~n9521 & pi1134;
  assign n9523 = ~n9522 & pi1136;
  assign n9524 = pi0648 & pi1135;
  assign n9525 = pi0619 & ~pi1135;
  assign n9526 = ~n9524 & ~n9525;
  assign n9527 = n9526 & ~pi1134;
  assign n9528 = n9523 & ~n9527;
  assign n9529 = n8517 & pi0838;
  assign n9530 = ~n9528 & ~n9529;
  assign n9531 = ~n9530 & n8354;
  assign po0890 = n9518 | n9531;
  assign n9533 = po0980 & ~pi1119;
  assign n9534 = ~n9533 & ~pi0962;
  assign n9535 = ~po0980 & pi0734;
  assign po0891 = n9534 & ~n9535;
  assign n9537 = po0980 & ~pi1109;
  assign n9538 = ~n9537 & ~pi0962;
  assign n9539 = ~po0980 & ~pi0735;
  assign po0892 = n9538 & ~n9539;
  assign n9541 = po0980 & ~pi1101;
  assign n9542 = ~n9541 & ~pi0962;
  assign n9543 = ~po0980 & ~pi0736;
  assign po0893 = n9542 & ~n9543;
  assign n9545 = po0980 & ~pi1122;
  assign n9546 = ~n9545 & ~pi0962;
  assign n9547 = ~po0980 & pi0737;
  assign po0894 = n9546 & ~n9547;
  assign n9549 = po0980 & ~pi1121;
  assign n9550 = ~n9549 & ~pi0962;
  assign n9551 = ~po0980 & pi0738;
  assign po0895 = n9550 & ~n9551;
  assign po0988 = n8048 & ~pi0952;
  assign n9554 = ~po0988 & pi0739;
  assign n9555 = ~n9554 & ~pi0966;
  assign n9556 = po0988 & pi1108;
  assign po0896 = ~n9555 | n9556;
  assign n9558 = ~po0988 & ~pi0741;
  assign n9559 = ~n9558 & ~pi0966;
  assign n9560 = po0988 & pi1114;
  assign po0898 = ~n9559 | n9560;
  assign n9562 = ~po0988 & ~pi0742;
  assign n9563 = ~n9562 & ~pi0966;
  assign n9564 = po0988 & pi1112;
  assign po0899 = ~n9563 | n9564;
  assign n9566 = ~po0988 & pi0743;
  assign n9567 = ~n9566 & ~pi0966;
  assign n9568 = po0988 & pi1109;
  assign po0900 = ~n9567 | n9568;
  assign n9570 = ~po0988 & ~pi0744;
  assign n9571 = ~n9570 & ~pi0966;
  assign n9572 = po0988 & pi1131;
  assign po0901 = ~n9571 | n9572;
  assign n9574 = ~po0988 & ~pi0745;
  assign n9575 = ~n9574 & ~pi0966;
  assign n9576 = po0988 & pi1111;
  assign po0902 = ~n9575 | n9576;
  assign n9578 = ~po0988 & pi0746;
  assign n9579 = ~n9578 & ~pi0966;
  assign n9580 = po0988 & pi1104;
  assign po0903 = ~n9579 | n9580;
  assign n9582 = n9494 & pi0773;
  assign n9583 = ~n9582 ^ ~pi0747;
  assign po0904 = ~po0978 & n9583;
  assign n9585 = ~po0988 & pi0748;
  assign n9586 = ~n9585 & ~pi0966;
  assign n9587 = po0988 & pi1106;
  assign po0905 = ~n9586 | n9587;
  assign n9589 = ~po0988 & pi0749;
  assign n9590 = ~n9589 & ~pi0966;
  assign n9591 = po0988 & pi1105;
  assign po0906 = ~n9590 | n9591;
  assign n9593 = ~po0988 & ~pi0750;
  assign n9594 = ~n9593 & ~pi0966;
  assign n9595 = po0988 & pi1130;
  assign po0907 = ~n9594 | n9595;
  assign n9597 = ~po0988 & ~pi0751;
  assign n9598 = ~n9597 & ~pi0966;
  assign n9599 = po0988 & pi1123;
  assign po0908 = ~n9598 | n9599;
  assign n9601 = ~po0988 & ~pi0752;
  assign n9602 = ~n9601 & ~pi0966;
  assign n9603 = po0988 & pi1124;
  assign po0909 = ~n9602 | n9603;
  assign n9605 = ~po0988 & ~pi0753;
  assign n9606 = ~n9605 & ~pi0966;
  assign n9607 = po0988 & pi1117;
  assign po0910 = ~n9606 | n9607;
  assign n9609 = ~po0988 & ~pi0754;
  assign n9610 = ~n9609 & ~pi0966;
  assign n9611 = po0988 & pi1118;
  assign po0911 = ~n9610 | n9611;
  assign n9613 = ~po0988 & ~pi0755;
  assign n9614 = ~n9613 & ~pi0966;
  assign n9615 = po0988 & pi1120;
  assign po0912 = ~n9614 | n9615;
  assign n9617 = ~po0988 & ~pi0756;
  assign n9618 = ~n9617 & ~pi0966;
  assign n9619 = po0988 & pi1119;
  assign po0913 = ~n9618 | n9619;
  assign n9621 = ~po0988 & ~pi0757;
  assign n9622 = ~n9621 & ~pi0966;
  assign n9623 = po0988 & pi1113;
  assign po0914 = ~n9622 | n9623;
  assign n9625 = ~po0988 & pi0758;
  assign n9626 = ~n9625 & ~pi0966;
  assign n9627 = po0988 & pi1101;
  assign po0915 = ~n9626 | n9627;
  assign n9629 = ~po0988 & pi0759;
  assign n9630 = ~n9629 & ~pi0966;
  assign n9631 = po0988 & pi1100;
  assign po0916 = ~n9630 | n9631;
  assign n9633 = ~po0988 & ~pi0760;
  assign n9634 = ~n9633 & ~pi0966;
  assign n9635 = po0988 & pi1115;
  assign po0917 = ~n9634 | n9635;
  assign n9637 = ~po0988 & ~pi0761;
  assign n9638 = ~n9637 & ~pi0966;
  assign n9639 = po0988 & pi1121;
  assign po0918 = ~n9638 | n9639;
  assign n9641 = ~po0988 & ~pi0762;
  assign n9642 = ~n9641 & ~pi0966;
  assign n9643 = po0988 & pi1129;
  assign po0919 = ~n9642 | n9643;
  assign n9645 = ~po0988 & pi0763;
  assign n9646 = ~n9645 & ~pi0966;
  assign n9647 = po0988 & pi1103;
  assign po0920 = ~n9646 | n9647;
  assign n9649 = ~po0988 & pi0764;
  assign n9650 = ~n9649 & ~pi0966;
  assign n9651 = po0988 & pi1107;
  assign po0921 = ~n9650 | n9651;
  assign n9653 = ~pi0773 & ~pi0794;
  assign n9654 = ~pi0795 & ~pi0816;
  assign n9655 = n9653 & n9654;
  assign n9656 = ~pi0721 & ~pi0747;
  assign n9657 = ~pi0765 & ~pi0771;
  assign n9658 = n9656 & n9657;
  assign n9659 = n9655 & n9658;
  assign po0963 = po0978 & ~n9659;
  assign n9661 = pi0765 ^ ~pi0945;
  assign po0922 = ~po0963 & n9661;
  assign n9663 = ~po0988 & pi0766;
  assign n9664 = ~n9663 & ~pi0966;
  assign n9665 = po0988 & pi1110;
  assign po0923 = ~n9664 | n9665;
  assign n9667 = ~po0988 & ~pi0767;
  assign n9668 = ~n9667 & ~pi0966;
  assign n9669 = po0988 & pi1116;
  assign po0924 = ~n9668 | n9669;
  assign n9671 = ~po0988 & ~pi0768;
  assign n9672 = ~n9671 & ~pi0966;
  assign n9673 = po0988 & pi1125;
  assign po0925 = ~n9672 | n9673;
  assign n9675 = ~n9411 ^ ~pi0769;
  assign po0926 = ~po0978 & n9675;
  assign n9677 = ~po0988 & ~pi0770;
  assign n9678 = ~n9677 & ~pi0966;
  assign n9679 = po0988 & pi1126;
  assign po0927 = ~n9678 | n9679;
  assign n9681 = ~pi0945 & pi0987;
  assign n9682 = pi0771 & pi0945;
  assign n9683 = ~n9681 & ~n9682;
  assign po0928 = ~po0963 & ~n9683;
  assign n9685 = ~po0988 & pi0772;
  assign n9686 = ~n9685 & ~pi0966;
  assign n9687 = po0988 & pi1102;
  assign po0929 = ~n9686 | n9687;
  assign n9689 = ~n9494 ^ ~pi0773;
  assign po0930 = ~po0963 & n9689;
  assign n9691 = ~po0988 & ~pi0774;
  assign n9692 = ~n9691 & ~pi0966;
  assign n9693 = po0988 & pi1127;
  assign po0931 = ~n9692 | n9693;
  assign n9695 = pi0765 & pi0771;
  assign n9696 = n9409 & n9695;
  assign n9697 = ~n9696 ^ ~pi0775;
  assign po0932 = ~po0978 & n9697;
  assign n9699 = ~po0988 & ~pi0776;
  assign n9700 = ~n9699 & ~pi0966;
  assign n9701 = po0988 & pi1128;
  assign po0933 = ~n9700 | n9701;
  assign n9703 = ~po0988 & ~pi0777;
  assign n9704 = ~n9703 & ~pi0966;
  assign n9705 = po0988 & pi1122;
  assign po0934 = ~n9704 | n9705;
  assign n9707 = pi0832 & pi0956;
  assign n9708 = ~pi1083 & pi1085;
  assign n9709 = n9707 & n9708;
  assign n9710 = n9709 & ~pi1046;
  assign n9711 = n9710 & ~pi0968;
  assign n9712 = n9711 & pi1100;
  assign n9713 = ~n9711 & pi0778;
  assign po0935 = n9712 | n9713;
  assign po0936 = n8105 | ~pi0779;
  assign po0937 = n8028 | ~pi0780;
  assign n9717 = n9711 & pi1101;
  assign n9718 = ~n9711 & pi0781;
  assign po0938 = n9717 | n9718;
  assign n9720 = ~n3415 & ~n8059;
  assign po0939 = n8027 | ~n9720;
  assign n9722 = n9711 & pi1109;
  assign n9723 = ~n9711 & pi0783;
  assign po0940 = n9722 | n9723;
  assign n9725 = n9711 & pi1110;
  assign n9726 = ~n9711 & pi0784;
  assign po0941 = n9725 | n9726;
  assign n9728 = n9711 & pi1102;
  assign n9729 = ~n9711 & pi0785;
  assign po0942 = n9728 | n9729;
  assign n9731 = pi0786 & pi0954;
  assign n9732 = pi0024 & ~pi0954;
  assign po0943 = ~n9731 & ~n9732;
  assign n9734 = n9711 & pi1104;
  assign n9735 = ~n9711 & pi0787;
  assign po0944 = n9734 | n9735;
  assign n9737 = n9711 & pi1105;
  assign n9738 = ~n9711 & pi0788;
  assign po0945 = n9737 | n9738;
  assign n9740 = n9711 & pi1106;
  assign n9741 = ~n9711 & pi0789;
  assign po0946 = n9740 | n9741;
  assign n9743 = n9711 & pi1107;
  assign n9744 = ~n9711 & pi0790;
  assign po0947 = n9743 | n9744;
  assign n9746 = n9711 & pi1108;
  assign n9747 = ~n9711 & pi0791;
  assign po0948 = n9746 | n9747;
  assign n9749 = n9711 & pi1103;
  assign n9750 = ~n9711 & pi0792;
  assign po0949 = n9749 | n9750;
  assign n9752 = n9710 & pi0968;
  assign n9753 = n9752 & pi1130;
  assign n9754 = ~n9752 & pi0794;
  assign po0951 = n9753 | n9754;
  assign n9756 = n9752 & pi1128;
  assign n9757 = ~n9752 & pi0795;
  assign po0952 = n9756 | n9757;
  assign n9759 = pi0266 & ~pi0269;
  assign n9760 = n9759 & pi0279;
  assign n9761 = pi0278 & ~pi0280;
  assign n9762 = n9760 & n9761;
  assign n9763 = n8296 & n8298;
  assign n9764 = n9762 & n9763;
  assign po0953 = n9764 ^ ~pi0264;
  assign n9766 = n9752 & pi1124;
  assign n9767 = ~n9752 & pi0798;
  assign po0955 = n9766 | n9767;
  assign n9769 = ~n9752 & pi0799;
  assign n9770 = n9752 & ~pi1107;
  assign po0956 = ~n9769 & ~n9770;
  assign n9772 = n9752 & pi1125;
  assign n9773 = ~n9752 & pi0800;
  assign po0957 = n9772 | n9773;
  assign n9775 = n9752 & pi1126;
  assign n9776 = ~n9752 & pi0801;
  assign po0958 = n9775 | n9776;
  assign po0959 = n8301 & ~pi0274;
  assign n9779 = ~n9752 & pi0803;
  assign n9780 = n9752 & ~pi1106;
  assign po0960 = ~n9779 & ~n9780;
  assign n9782 = n9752 & pi1109;
  assign n9783 = ~n9752 & pi0804;
  assign po0961 = n9782 | n9783;
  assign po0962 = n8297 ^ ~pi0270;
  assign n9786 = n9752 & pi1127;
  assign n9787 = ~n9752 & pi0807;
  assign po0964 = n9786 | n9787;
  assign n9789 = n9752 & pi1101;
  assign n9790 = ~n9752 & pi0808;
  assign po0965 = n9789 | n9790;
  assign n9792 = ~n9752 & pi0809;
  assign n9793 = n9752 & ~pi1103;
  assign po0966 = ~n9792 & ~n9793;
  assign n9795 = n9752 & pi1108;
  assign n9796 = ~n9752 & pi0810;
  assign po0967 = n9795 | n9796;
  assign n9798 = n9752 & pi1102;
  assign n9799 = ~n9752 & pi0811;
  assign po0968 = n9798 | n9799;
  assign n9801 = ~n9752 & pi0812;
  assign n9802 = n9752 & ~pi1104;
  assign po0969 = ~n9801 & ~n9802;
  assign n9804 = n9752 & pi1131;
  assign n9805 = ~n9752 & pi0813;
  assign po0970 = n9804 | n9805;
  assign n9807 = ~n9752 & pi0814;
  assign n9808 = n9752 & ~pi1105;
  assign po0971 = ~n9807 & ~n9808;
  assign n9810 = n9752 & pi1110;
  assign n9811 = ~n9752 & pi0815;
  assign po0972 = n9810 | n9811;
  assign n9813 = n9752 & pi1129;
  assign n9814 = ~n9752 & pi0816;
  assign po0973 = n9813 | n9814;
  assign po0974 = n8294 ^ ~pi0269;
  assign po0975 = n5003 | n4999;
  assign po0976 = n8300 ^ ~pi0265;
  assign n9819 = n8297 & ~pi0270;
  assign po0977 = n9819 ^ ~pi0277;
  assign po0979 = ~pi0811 & ~pi0893;
  assign n9822 = n3927 & n2643;
  assign n9823 = ~n2642 & ~pi0982;
  assign n9824 = ~n9822 & ~n9823;
  assign po0981 = ~n9824 & n2645;
  assign n9826 = n2713 & pi0123;
  assign n9827 = n9826 & ~pi0825;
  assign n9828 = ~pi1126 ^ ~pi1127;
  assign n9829 = ~pi1124 ^ ~pi1125;
  assign n9830 = n9828 ^ ~n9829;
  assign n9831 = pi1128 ^ ~pi1129;
  assign n9832 = pi1130 ^ ~pi1131;
  assign n9833 = ~n9831 ^ ~n9832;
  assign n9834 = ~n9830 ^ ~n9833;
  assign n9835 = ~n9826 & ~n9834;
  assign po0982 = n9827 | n9835;
  assign n9837 = n9826 & ~pi0826;
  assign n9838 = ~pi1118 ^ ~pi1119;
  assign n9839 = ~pi1116 ^ ~pi1117;
  assign n9840 = n9838 ^ ~n9839;
  assign n9841 = pi1120 ^ ~pi1121;
  assign n9842 = pi1122 ^ ~pi1123;
  assign n9843 = ~n9841 ^ ~n9842;
  assign n9844 = ~n9840 ^ ~n9843;
  assign n9845 = ~n9826 & ~n9844;
  assign po0983 = n9837 | n9845;
  assign n9847 = n9826 & ~pi0827;
  assign n9848 = ~pi1100 ^ ~pi1101;
  assign n9849 = pi1102 ^ ~pi1103;
  assign n9850 = ~n9848 ^ ~n9849;
  assign n9851 = ~pi1104 ^ ~pi1105;
  assign n9852 = pi1106 ^ ~pi1107;
  assign n9853 = n9851 ^ ~n9852;
  assign n9854 = ~n9850 ^ ~n9853;
  assign n9855 = ~n9826 & ~n9854;
  assign po0984 = n9847 | n9855;
  assign n9857 = n9826 & ~pi0828;
  assign n9858 = pi1114 ^ ~pi1115;
  assign n9859 = ~pi1112 ^ ~pi1113;
  assign n9860 = ~n9858 ^ ~n9859;
  assign n9861 = pi1110 ^ ~pi1111;
  assign n9862 = ~pi1108 ^ ~pi1109;
  assign n9863 = n9861 ^ ~n9862;
  assign n9864 = ~n9860 ^ ~n9863;
  assign n9865 = ~n9826 & ~n9864;
  assign po0985 = n9857 | n9865;
  assign n9867 = n3923 & pi1091;
  assign n9868 = n3927 & n9867;
  assign n9869 = ~pi0951 & pi1092;
  assign po0986 = n9868 | n9869;
  assign po0987 = n9762 ^ ~pi0281;
  assign n9872 = ~pi0832 & ~pi1163;
  assign n9873 = n3962 & n9872;
  assign po0989 = n9867 & n9873;
  assign n9875 = ~n3923 & pi0833;
  assign po0990 = n9867 | n9875;
  assign po0991 = n3923 & pi0946;
  assign n9878 = n8295 & ~pi0281;
  assign po0992 = n9878 ^ ~pi0282;
  assign n9880 = pi0837 & pi0955;
  assign n9881 = ~pi0955 & pi1049;
  assign po0993 = n9880 | n9881;
  assign n9883 = pi0838 & pi0955;
  assign n9884 = ~pi0955 & pi1047;
  assign po0994 = n9883 | n9884;
  assign n9886 = pi0839 & pi0955;
  assign n9887 = ~pi0955 & pi1074;
  assign po0995 = n9886 | n9887;
  assign n9889 = n3923 & pi1196;
  assign n9890 = ~n3923 & pi0840;
  assign po0996 = n9889 | n9890;
  assign n9892 = pi0842 & pi0955;
  assign n9893 = ~pi0955 & pi1035;
  assign po0998 = n9892 | n9893;
  assign n9895 = pi0843 & pi0955;
  assign n9896 = ~pi0955 & pi1079;
  assign po0999 = n9895 | n9896;
  assign n9898 = pi0844 & pi0955;
  assign n9899 = ~pi0955 & pi1078;
  assign po1000 = n9898 | n9899;
  assign n9901 = pi0845 & pi0955;
  assign n9902 = ~pi0955 & pi1043;
  assign po1001 = n9901 | n9902;
  assign n9904 = n6516 & pi0846;
  assign n9905 = ~n6516 & pi1134;
  assign po1002 = n9904 | n9905;
  assign n9907 = pi0847 & pi0955;
  assign n9908 = ~pi0955 & pi1055;
  assign po1003 = n9907 | n9908;
  assign n9910 = pi0848 & pi0955;
  assign n9911 = ~pi0955 & pi1039;
  assign po1004 = n9910 | n9911;
  assign n9913 = n3923 & pi1198;
  assign n9914 = ~n3923 & pi0849;
  assign po1005 = n9913 | n9914;
  assign n9916 = pi0850 & pi0955;
  assign n9917 = ~pi0955 & pi1048;
  assign po1006 = n9916 | n9917;
  assign n9919 = pi0851 & pi0955;
  assign n9920 = ~pi0955 & pi1045;
  assign po1007 = n9919 | n9920;
  assign n9922 = pi0852 & pi0955;
  assign n9923 = ~pi0955 & pi1062;
  assign po1008 = n9922 | n9923;
  assign n9925 = pi0853 & pi0955;
  assign n9926 = ~pi0955 & pi1080;
  assign po1009 = n9925 | n9926;
  assign n9928 = pi0854 & pi0955;
  assign n9929 = ~pi0955 & pi1051;
  assign po1010 = n9928 | n9929;
  assign n9931 = pi0855 & pi0955;
  assign n9932 = ~pi0955 & pi1065;
  assign po1011 = n9931 | n9932;
  assign n9934 = pi0856 & pi0955;
  assign n9935 = ~pi0955 & pi1067;
  assign po1012 = n9934 | n9935;
  assign n9937 = pi0857 & pi0955;
  assign n9938 = ~pi0955 & pi1058;
  assign po1013 = n9937 | n9938;
  assign n9940 = pi0858 & pi0955;
  assign n9941 = ~pi0955 & pi1087;
  assign po1014 = n9940 | n9941;
  assign n9943 = pi0859 & pi0955;
  assign n9944 = ~pi0955 & pi1070;
  assign po1015 = n9943 | n9944;
  assign n9946 = pi0860 & pi0955;
  assign n9947 = ~pi0955 & pi1076;
  assign po1016 = n9946 | n9947;
  assign n9949 = n6516 & pi0861;
  assign n9950 = ~n6516 & pi1141;
  assign po1017 = n9949 | n9950;
  assign n9952 = n6516 & pi0862;
  assign n9953 = ~n6516 & pi1139;
  assign po1018 = n9952 | n9953;
  assign n9955 = n3923 & pi1199;
  assign n9956 = ~n3923 & pi0863;
  assign po1019 = n9955 | n9956;
  assign n9958 = n3923 & pi1197;
  assign n9959 = ~n3923 & pi0864;
  assign po1020 = n9958 | n9959;
  assign n9961 = pi0865 & pi0955;
  assign n9962 = ~pi0955 & pi1040;
  assign po1021 = n9961 | n9962;
  assign n9964 = pi0866 & pi0955;
  assign n9965 = ~pi0955 & pi1053;
  assign po1022 = n9964 | n9965;
  assign n9967 = pi0867 & pi0955;
  assign n9968 = ~pi0955 & pi1057;
  assign po1023 = n9967 | n9968;
  assign n9970 = pi0868 & pi0955;
  assign n9971 = ~pi0955 & pi1063;
  assign po1024 = n9970 | n9971;
  assign n9973 = n6516 & pi0869;
  assign n9974 = ~n6516 & pi1140;
  assign po1025 = n9973 | n9974;
  assign n9976 = pi0870 & pi0955;
  assign n9977 = ~pi0955 & pi1069;
  assign po1026 = n9976 | n9977;
  assign n9979 = pi0871 & pi0955;
  assign n9980 = ~pi0955 & pi1072;
  assign po1027 = n9979 | n9980;
  assign n9982 = pi0872 & pi0955;
  assign n9983 = ~pi0955 & pi1084;
  assign po1028 = n9982 | n9983;
  assign n9985 = pi0873 & pi0955;
  assign n9986 = ~pi0955 & pi1044;
  assign po1029 = n9985 | n9986;
  assign n9988 = pi0874 & pi0955;
  assign n9989 = ~pi0955 & pi1036;
  assign po1030 = n9988 | n9989;
  assign n9991 = n6516 & pi0875;
  assign n9992 = ~n6516 & pi1136;
  assign po1031 = n9991 | n9992;
  assign n9994 = pi0876 & pi0955;
  assign n9995 = ~pi0955 & pi1037;
  assign po1032 = n9994 | n9995;
  assign n9997 = n6516 & pi0877;
  assign n9998 = ~n6516 & pi1138;
  assign po1033 = n9997 | n9998;
  assign n10000 = n6516 & pi0878;
  assign n10001 = ~n6516 & pi1137;
  assign po1034 = n10000 | n10001;
  assign n10003 = n6516 & pi0879;
  assign n10004 = ~n6516 & pi1135;
  assign po1035 = n10003 | n10004;
  assign n10006 = pi0880 & pi0955;
  assign n10007 = ~pi0955 & pi1081;
  assign po1036 = n10006 | n10007;
  assign n10009 = pi0881 & pi0955;
  assign n10010 = ~pi0955 & pi1059;
  assign po1037 = n10009 | n10010;
  assign n10012 = ~n9826 & pi1107;
  assign n10013 = n9826 & ~pi0883;
  assign po1039 = n10012 | n10013;
  assign n10015 = ~n9826 & pi1124;
  assign n10016 = n9826 & ~pi0884;
  assign po1040 = n10015 | n10016;
  assign n10018 = ~n9826 & pi1125;
  assign n10019 = n9826 & ~pi0885;
  assign po1041 = n10018 | n10019;
  assign n10021 = ~n9826 & pi1109;
  assign n10022 = n9826 & ~pi0886;
  assign po1042 = n10021 | n10022;
  assign n10024 = ~n9826 & pi1100;
  assign n10025 = n9826 & ~pi0887;
  assign po1043 = n10024 | n10025;
  assign n10027 = ~n9826 & pi1120;
  assign n10028 = n9826 & ~pi0888;
  assign po1044 = n10027 | n10028;
  assign n10030 = ~n9826 & pi1103;
  assign n10031 = n9826 & ~pi0889;
  assign po1045 = n10030 | n10031;
  assign n10033 = ~n9826 & pi1126;
  assign n10034 = n9826 & ~pi0890;
  assign po1046 = n10033 | n10034;
  assign n10036 = ~n9826 & pi1116;
  assign n10037 = n9826 & ~pi0891;
  assign po1047 = n10036 | n10037;
  assign n10039 = ~n9826 & pi1101;
  assign n10040 = n9826 & ~pi0892;
  assign po1048 = n10039 | n10040;
  assign n10042 = ~n9826 & pi1119;
  assign n10043 = n9826 & ~pi0894;
  assign po1050 = n10042 | n10043;
  assign n10045 = ~n9826 & pi1113;
  assign n10046 = n9826 & ~pi0895;
  assign po1051 = n10045 | n10046;
  assign n10048 = ~n9826 & pi1118;
  assign n10049 = n9826 & ~pi0896;
  assign po1052 = n10048 | n10049;
  assign n10051 = ~n9826 & pi1129;
  assign n10052 = n9826 & ~pi0898;
  assign po1054 = n10051 | n10052;
  assign n10054 = ~n9826 & pi1115;
  assign n10055 = n9826 & ~pi0899;
  assign po1055 = n10054 | n10055;
  assign n10057 = ~n9826 & pi1110;
  assign n10058 = n9826 & ~pi0900;
  assign po1056 = n10057 | n10058;
  assign n10060 = ~n9826 & pi1111;
  assign n10061 = n9826 & ~pi0902;
  assign po1058 = n10060 | n10061;
  assign n10063 = ~n9826 & pi1121;
  assign n10064 = n9826 & ~pi0903;
  assign po1059 = n10063 | n10064;
  assign n10066 = ~n9826 & pi1127;
  assign n10067 = n9826 & ~pi0904;
  assign po1060 = n10066 | n10067;
  assign n10069 = ~n9826 & pi1131;
  assign n10070 = n9826 & ~pi0905;
  assign po1061 = n10069 | n10070;
  assign n10072 = ~n9826 & pi1128;
  assign n10073 = n9826 & ~pi0906;
  assign po1062 = n10072 | n10073;
  assign n10075 = ~pi0624 & ~pi0979;
  assign n10076 = n10075 & pi0604;
  assign n10077 = ~pi0598 & pi0979;
  assign n10078 = n10077 & ~pi0615;
  assign n10079 = ~n10076 & ~n10078;
  assign n10080 = n10079 & pi0782;
  assign n10081 = ~pi0782 & ~pi0907;
  assign po1063 = ~n10080 & ~n10081;
  assign n10083 = ~n9826 & pi1122;
  assign n10084 = n9826 & ~pi0908;
  assign po1064 = n10083 | n10084;
  assign n10086 = ~n9826 & pi1105;
  assign n10087 = n9826 & ~pi0909;
  assign po1065 = n10086 | n10087;
  assign n10089 = ~n9826 & pi1117;
  assign n10090 = n9826 & ~pi0910;
  assign po1066 = n10089 | n10090;
  assign n10092 = ~n9826 & pi1130;
  assign n10093 = n9826 & ~pi0911;
  assign po1067 = n10092 | n10093;
  assign n10095 = ~n9826 & pi1114;
  assign n10096 = n9826 & ~pi0912;
  assign po1068 = n10095 | n10096;
  assign n10098 = ~n9826 & pi1106;
  assign n10099 = n9826 & ~pi0913;
  assign po1069 = n10098 | n10099;
  assign po1070 = n8293 ^ ~pi0280;
  assign n10102 = ~n9826 & pi1108;
  assign n10103 = n9826 & ~pi0915;
  assign po1071 = n10102 | n10103;
  assign n10105 = ~n9826 & pi1123;
  assign n10106 = n9826 & ~pi0916;
  assign po1072 = n10105 | n10106;
  assign n10108 = ~n9826 & pi1112;
  assign n10109 = n9826 & ~pi0917;
  assign po1073 = n10108 | n10109;
  assign n10111 = ~n9826 & pi1104;
  assign n10112 = n9826 & ~pi0918;
  assign po1074 = n10111 | n10112;
  assign n10114 = ~n9826 & pi1102;
  assign n10115 = n9826 & ~pi0919;
  assign po1075 = n10114 | n10115;
  assign n10117 = pi1093 & pi1139;
  assign n10118 = pi0920 & ~pi1093;
  assign po1076 = n10117 | n10118;
  assign n10120 = pi1093 & pi1140;
  assign n10121 = pi0921 & ~pi1093;
  assign po1077 = n10120 | n10121;
  assign n10123 = pi1093 & pi1152;
  assign n10124 = pi0922 & ~pi1093;
  assign po1078 = n10123 | n10124;
  assign n10126 = pi1093 & pi1154;
  assign n10127 = pi0923 & ~pi1093;
  assign po1079 = n10126 | n10127;
  assign po1080 = n6856 & pi0311;
  assign n10130 = pi1093 & pi1155;
  assign n10131 = pi0925 & ~pi1093;
  assign po1081 = n10130 | n10131;
  assign n10133 = pi1093 & pi1157;
  assign n10134 = pi0926 & ~pi1093;
  assign po1082 = n10133 | n10134;
  assign n10136 = pi1093 & pi1145;
  assign n10137 = pi0927 & ~pi1093;
  assign po1083 = n10136 | n10137;
  assign n10139 = pi1093 & pi1136;
  assign n10140 = pi0928 & ~pi1093;
  assign po1084 = n10139 | n10140;
  assign n10142 = pi1093 & pi1144;
  assign n10143 = pi0929 & ~pi1093;
  assign po1085 = n10142 | n10143;
  assign n10145 = pi1093 & pi1134;
  assign n10146 = pi0930 & ~pi1093;
  assign po1086 = n10145 | n10146;
  assign n10148 = pi1093 & pi1150;
  assign n10149 = pi0931 & ~pi1093;
  assign po1087 = n10148 | n10149;
  assign n10151 = pi1093 & pi1142;
  assign n10152 = pi0932 & ~pi1093;
  assign po1088 = n10151 | n10152;
  assign n10154 = pi1093 & pi1137;
  assign n10155 = pi0933 & ~pi1093;
  assign po1089 = n10154 | n10155;
  assign n10157 = pi1093 & pi1147;
  assign n10158 = pi0934 & ~pi1093;
  assign po1090 = n10157 | n10158;
  assign n10160 = pi1093 & pi1141;
  assign n10161 = pi0935 & ~pi1093;
  assign po1091 = n10160 | n10161;
  assign n10163 = pi1093 & pi1149;
  assign n10164 = pi0936 & ~pi1093;
  assign po1092 = n10163 | n10164;
  assign n10166 = pi1093 & pi1148;
  assign n10167 = pi0937 & ~pi1093;
  assign po1093 = n10166 | n10167;
  assign n10169 = pi1093 & pi1135;
  assign n10170 = pi0938 & ~pi1093;
  assign po1094 = n10169 | n10170;
  assign n10172 = pi1093 & pi1146;
  assign n10173 = pi0939 & ~pi1093;
  assign po1095 = n10172 | n10173;
  assign n10175 = pi1093 & pi1138;
  assign n10176 = pi0940 & ~pi1093;
  assign po1096 = n10175 | n10176;
  assign n10178 = pi1093 & pi1153;
  assign n10179 = pi0941 & ~pi1093;
  assign po1097 = n10178 | n10179;
  assign n10181 = pi1093 & pi1156;
  assign n10182 = pi0942 & ~pi1093;
  assign po1098 = n10181 | n10182;
  assign n10184 = pi1093 & pi1151;
  assign n10185 = pi0943 & ~pi1093;
  assign po1099 = n10184 | n10185;
  assign n10187 = pi1093 & pi1143;
  assign n10188 = pi0944 & ~pi1093;
  assign po1100 = n10187 | n10188;
  assign po1102 = n3923 & pi0230;
  assign n10191 = ~n10075 & ~n10077;
  assign n10192 = ~n10191 & pi0782;
  assign n10193 = ~pi0782 & ~pi0947;
  assign po1103 = ~n10192 & ~n10193;
  assign po1104 = ~pi0266 ^ ~pi0992;
  assign n10196 = pi0313 & ~pi0954;
  assign n10197 = ~pi0949 & pi0954;
  assign po1105 = ~n10196 & ~n10197;
  assign po1106 = n2642 & pi1092;
  assign n10200 = pi0957 & pi1092;
  assign po1112 = n10200 | pi0031;
  assign po1115 = ~pi0782 & pi0960;
  assign po1116 = ~pi0230 & pi0961;
  assign po1118 = ~pi0782 & pi0963;
  assign po1122 = ~pi0230 & pi0967;
  assign po1124 = ~pi0230 & pi0969;
  assign po1125 = ~pi0782 & pi0970;
  assign po1126 = ~pi0230 & pi0971;
  assign po1127 = ~pi0782 & pi0972;
  assign po1128 = ~pi0230 & pi0974;
  assign po1129 = ~pi0782 & pi0975;
  assign po1131 = ~pi0230 & pi0977;
  assign po1132 = ~pi0782 & pi0978;
  assign po1133 = pi0598 | ~pi0615;
  assign po1135 = pi0824 & pi1092;
  assign po1137 = pi0604 | pi0624;
  assign po0166 = 1'b1;
  assign po0170 = ~pi1090;
  assign po1110 = ~pi0954;
  assign po1130 = ~pi0278;
  assign po1146 = ~pi0915;
  assign po1147 = ~pi0825;
  assign po1148 = ~pi0826;
  assign po1149 = ~pi0913;
  assign po1150 = ~pi0894;
  assign po1151 = ~pi0905;
  assign po1153 = ~pi0890;
  assign po1155 = ~pi0906;
  assign po1156 = ~pi0896;
  assign po1157 = ~pi0909;
  assign po1158 = ~pi0911;
  assign po1159 = ~pi0908;
  assign po1160 = ~pi0891;
  assign po1161 = ~pi0902;
  assign po1162 = ~pi0903;
  assign po1163 = ~pi0883;
  assign po1164 = ~pi0888;
  assign po1165 = ~pi0919;
  assign po1166 = ~pi0886;
  assign po1167 = ~pi0912;
  assign po1168 = ~pi0895;
  assign po1169 = ~pi0916;
  assign po1170 = ~pi0889;
  assign po1171 = ~pi0900;
  assign po1172 = ~pi0885;
  assign po1173 = ~pi0904;
  assign po1174 = ~pi0899;
  assign po1175 = ~pi0918;
  assign po1176 = ~pi0898;
  assign po1177 = ~pi0917;
  assign po1178 = ~pi0827;
  assign po1179 = ~pi0887;
  assign po1180 = ~pi0884;
  assign po1181 = ~pi0910;
  assign po1182 = ~pi0828;
  assign po1183 = ~pi0892;
  assign po0000 = pi0668;
  assign po0001 = pi0672;
  assign po0002 = pi0664;
  assign po0003 = pi0667;
  assign po0004 = pi0676;
  assign po0005 = pi0673;
  assign po0006 = pi0675;
  assign po0007 = pi0666;
  assign po0008 = pi0679;
  assign po0009 = pi0674;
  assign po0010 = pi0663;
  assign po0011 = pi0670;
  assign po0012 = pi0677;
  assign po0013 = pi0682;
  assign po0014 = pi0671;
  assign po0015 = pi0678;
  assign po0016 = pi0718;
  assign po0017 = pi0707;
  assign po0018 = pi0708;
  assign po0019 = pi0713;
  assign po0020 = pi0711;
  assign po0021 = pi0716;
  assign po0022 = pi0733;
  assign po0023 = pi0712;
  assign po0024 = pi0689;
  assign po0025 = pi0717;
  assign po0026 = pi0692;
  assign po0027 = pi0719;
  assign po0028 = pi0722;
  assign po0029 = pi0714;
  assign po0030 = pi0720;
  assign po0031 = pi0685;
  assign po0032 = pi0837;
  assign po0033 = pi0850;
  assign po0034 = pi0872;
  assign po0035 = pi0871;
  assign po0036 = pi0881;
  assign po0037 = pi0866;
  assign po0038 = pi0876;
  assign po0039 = pi0873;
  assign po0040 = pi0874;
  assign po0041 = pi0859;
  assign po0042 = pi0855;
  assign po0043 = pi0852;
  assign po0044 = pi0870;
  assign po0045 = pi0848;
  assign po0046 = pi0865;
  assign po0047 = pi0856;
  assign po0048 = pi0853;
  assign po0049 = pi0847;
  assign po0050 = pi0857;
  assign po0051 = pi0854;
  assign po0052 = pi0858;
  assign po0053 = pi0845;
  assign po0054 = pi0838;
  assign po0055 = pi0842;
  assign po0056 = pi0843;
  assign po0057 = pi0839;
  assign po0058 = pi0844;
  assign po0059 = pi0868;
  assign po0060 = pi0851;
  assign po0061 = pi0867;
  assign po0062 = pi0880;
  assign po0063 = pi0860;
  assign po0064 = pi1030;
  assign po0065 = pi1034;
  assign po0066 = pi1015;
  assign po0067 = pi1020;
  assign po0068 = pi1025;
  assign po0069 = pi1005;
  assign po0070 = pi0996;
  assign po0071 = pi1012;
  assign po0072 = pi0993;
  assign po0073 = pi1016;
  assign po0074 = pi1021;
  assign po0075 = pi1010;
  assign po0076 = pi1027;
  assign po0077 = pi1018;
  assign po0078 = pi1017;
  assign po0079 = pi1024;
  assign po0080 = pi1009;
  assign po0081 = pi1032;
  assign po0082 = pi1003;
  assign po0083 = pi0997;
  assign po0084 = pi1013;
  assign po0085 = pi1011;
  assign po0086 = pi1008;
  assign po0087 = pi1019;
  assign po0088 = pi1031;
  assign po0089 = pi1022;
  assign po0090 = pi1000;
  assign po0091 = pi1023;
  assign po0092 = pi1002;
  assign po0093 = pi1026;
  assign po0094 = pi1006;
  assign po0095 = pi0998;
  assign po0096 = pi0031;
  assign po0097 = pi0080;
  assign po0098 = pi0893;
  assign po0099 = pi0467;
  assign po0100 = pi0078;
  assign po0101 = pi0112;
  assign po0102 = pi0013;
  assign po0103 = pi0025;
  assign po0104 = pi0226;
  assign po0105 = pi0127;
  assign po0106 = pi0822;
  assign po0107 = pi0808;
  assign po0108 = pi0227;
  assign po0109 = pi0477;
  assign po0110 = pi0834;
  assign po0111 = pi0229;
  assign po0112 = pi0012;
  assign po0113 = pi0011;
  assign po0114 = pi0010;
  assign po0115 = pi0009;
  assign po0116 = pi0008;
  assign po0117 = pi0007;
  assign po0118 = pi0006;
  assign po0119 = pi0005;
  assign po0120 = pi0004;
  assign po0121 = pi0003;
  assign po0122 = pi0000;
  assign po0123 = pi0002;
  assign po0124 = pi0001;
  assign po0125 = pi0310;
  assign po0126 = pi0302;
  assign po0127 = pi0475;
  assign po0128 = pi0474;
  assign po0129 = pi0466;
  assign po0130 = pi0473;
  assign po0131 = pi0471;
  assign po0132 = pi0472;
  assign po0133 = pi0470;
  assign po0134 = pi0469;
  assign po0135 = pi0465;
  assign po0136 = pi1028;
  assign po0137 = pi1033;
  assign po0138 = pi0995;
  assign po0139 = pi0994;
  assign po0140 = pi0028;
  assign po0141 = pi0027;
  assign po0142 = pi0026;
  assign po0143 = pi0029;
  assign po0144 = pi0015;
  assign po0145 = pi0014;
  assign po0146 = pi0021;
  assign po0147 = pi0020;
  assign po0148 = pi0019;
  assign po0149 = pi0018;
  assign po0150 = pi0017;
  assign po0151 = pi0016;
  assign po0152 = pi1096;
  assign po0168 = pi0228;
  assign po0169 = pi0022;
  assign po0179 = pi1089;
  assign po0180 = pi0023;
  assign po0181 = po0167;
  assign po0188 = pi0037;
  assign po0263 = pi0117;
  assign po0285 = pi0131;
  assign po0386 = pi0232;
  assign po0388 = pi0236;
  assign po0636 = pi0583;
  assign po1053 = pi0067;
  assign po1108 = pi1134;
  assign po1109 = pi0964;
  assign po1111 = pi0965;
  assign po1113 = pi0991;
  assign po1114 = pi0985;
  assign po1117 = pi1014;
  assign po1119 = pi1029;
  assign po1120 = pi1004;
  assign po1121 = pi1007;
  assign po1123 = pi1135;
  assign po1134 = pi1064;
  assign po1136 = pi0299;
  assign po1138 = pi1075;
  assign po1139 = pi1052;
  assign po1140 = pi0771;
  assign po1141 = pi0765;
  assign po1142 = pi0605;
  assign po1143 = pi0601;
  assign po1144 = pi0278;
  assign po1145 = pi0279;
  assign po1152 = pi1095;
  assign po1154 = pi1094;
  assign po1184 = pi1187;
  assign po1185 = pi1172;
  assign po1186 = pi1170;
  assign po1187 = pi1138;
  assign po1188 = pi1177;
  assign po1189 = pi1178;
  assign po1190 = pi0863;
  assign po1191 = pi1203;
  assign po1192 = pi1185;
  assign po1193 = pi1171;
  assign po1194 = pi1192;
  assign po1195 = pi1137;
  assign po1196 = pi1186;
  assign po1197 = pi1165;
  assign po1198 = pi1164;
  assign po1199 = pi1098;
  assign po1200 = pi1183;
  assign po1201 = pi0230;
  assign po1202 = pi1169;
  assign po1203 = pi1136;
  assign po1204 = pi1181;
  assign po1205 = pi0849;
  assign po1206 = pi1193;
  assign po1207 = pi1182;
  assign po1208 = pi1168;
  assign po1209 = pi1175;
  assign po1210 = pi1191;
  assign po1211 = pi1099;
  assign po1212 = pi1174;
  assign po1213 = pi1179;
  assign po1214 = pi1202;
  assign po1215 = pi1176;
  assign po1216 = pi1173;
  assign po1217 = pi1201;
  assign po1218 = pi1167;
  assign po1219 = pi0840;
  assign po1220 = pi1189;
  assign po1221 = pi1195;
  assign po1222 = pi0864;
  assign po1223 = pi1190;
  assign po1224 = pi1188;
  assign po1225 = pi1180;
  assign po1226 = pi1194;
  assign po1227 = pi1097;
  assign po1228 = pi1166;
  assign po1229 = pi1200;
  assign po1230 = pi1184;
endmodule


