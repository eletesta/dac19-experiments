module top(x0, x1, x2, x3, x4, x5, x6, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25);
  input x0, x1, x2, x3, x4, x5, x6;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25;
  wire n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95;
  assign n8 = x3 & x4;
  assign n9 = ~x0 & ~x1;
  assign n10 = n8 & ~n9;
  assign n11 = x2 & n8;
  assign n12 = ~n10 & ~n11;
  assign n13 = x2 & ~x3;
  assign n14 = x1 & ~x4;
  assign n15 = n13 & n14;
  assign n16 = n12 & ~n15;
  assign n17 = ~x2 & x3;
  assign n18 = x4 & n17;
  assign n19 = n9 & n18;
  assign n20 = ~n15 & ~n19;
  assign n21 = x1 & ~x3;
  assign n22 = ~x2 & x4;
  assign n23 = n21 & n22;
  assign n24 = n20 & ~n23;
  assign n25 = ~x0 & n22;
  assign n26 = x2 & ~x4;
  assign n27 = ~n25 & ~n26;
  assign n28 = n21 & ~n27;
  assign n29 = ~x1 & x4;
  assign n30 = n17 & n29;
  assign n31 = ~n28 & ~n30;
  assign n32 = n25 & ~n31;
  assign n33 = n14 & n17;
  assign n34 = ~n32 & ~n33;
  assign n35 = ~x1 & n17;
  assign n36 = ~x3 & x4;
  assign n37 = ~n35 & ~n36;
  assign n38 = ~n10 & ~n37;
  assign n39 = x4 & n13;
  assign n40 = ~n33 & ~n39;
  assign n41 = x0 & ~n40;
  assign n42 = n17 & ~n29;
  assign n43 = x5 & n8;
  assign n44 = n42 & n43;
  assign n45 = x0 & x1;
  assign n46 = ~x6 & n45;
  assign n47 = n44 & ~n46;
  assign n48 = ~n41 & ~n47;
  assign n49 = x4 & ~x6;
  assign n50 = n17 & ~n49;
  assign n51 = ~n39 & ~n50;
  assign n52 = x1 & ~n51;
  assign n53 = n18 & ~n45;
  assign n54 = x3 ^ x2;
  assign n55 = ~x4 & ~n54;
  assign n56 = ~n13 & ~n55;
  assign n57 = ~n53 & n56;
  assign n58 = x0 & n11;
  assign n59 = n20 & ~n58;
  assign n60 = x1 & n11;
  assign n61 = ~n28 & ~n60;
  assign n62 = ~n28 & n36;
  assign n63 = ~n42 & ~n62;
  assign n64 = ~x3 & n9;
  assign n65 = n55 & n64;
  assign n66 = ~x1 & ~x3;
  assign n67 = ~n27 & n66;
  assign n68 = ~n55 & ~n67;
  assign n69 = ~x4 & n13;
  assign n70 = x0 & n69;
  assign n71 = ~x0 & n69;
  assign n72 = x3 & n26;
  assign n73 = n9 & n72;
  assign n74 = x0 & ~x1;
  assign n75 = n72 & n74;
  assign n76 = n45 & n72;
  assign n77 = ~x0 & x1;
  assign n78 = n72 & n77;
  assign n79 = x4 & ~x5;
  assign n80 = ~x2 & ~n79;
  assign n81 = x0 & ~n29;
  assign n82 = n80 & n81;
  assign n83 = x2 & x4;
  assign n84 = ~n45 & n83;
  assign n85 = ~n82 & ~n84;
  assign n86 = x3 & ~n85;
  assign n87 = n45 & ~n49;
  assign n88 = n80 & n87;
  assign n89 = ~n84 & ~n88;
  assign n90 = n86 & n89;
  assign n91 = x3 & ~n89;
  assign n92 = ~x2 & n36;
  assign n93 = x1 ^ x0;
  assign n94 = n92 & ~n93;
  assign n95 = n74 & n92;
  assign y0 = ~n16;
  assign y1 = ~n24;
  assign y2 = ~n34;
  assign y3 = n38;
  assign y4 = ~n48;
  assign y5 = n52;
  assign y6 = n57;
  assign y7 = ~n59;
  assign y8 = ~n61;
  assign y9 = ~n31;
  assign y10 = ~n63;
  assign y11 = n65;
  assign y12 = n68;
  assign y13 = n70;
  assign y14 = n71;
  assign y15 = n73;
  assign y16 = n75;
  assign y17 = n76;
  assign y18 = n78;
  assign y19 = n69;
  assign y20 = n86;
  assign y21 = n90;
  assign y22 = n91;
  assign y23 = ~1'b0;
  assign y24 = n94;
  assign y25 = n95;
endmodule
