module top(n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n375);
  input n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63;
  output n375;
  wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374;
  assign n348 = ~n38;
  assign n352 = ~n27;
  assign n361 = ~n49;
  assign n346 = ~n45;
  assign n363 = ~n41;
  assign n354 = ~n50;
  assign n373 = ~n63;
  assign n259 = ~n10;
  assign n350 = ~n44;
  assign n369 = ~n7;
  assign n166 = ~n4;
  assign n345 = ~n54;
  assign n267 = ~n6;
  assign n355 = ~n52;
  assign n276 = ~n28;
  assign n366 = ~n39;
  assign n229 = ~n51;
  assign n347 = ~n20;
  assign n372 = ~n59;
  assign n289 = ~n19;
  assign n336 = ~n9;
  assign n342 = ~n15;
  assign n353 = ~n3;
  assign n367 = ~n17;
  assign n237 = ~n5;
  assign n164 = ~n24;
  assign n281 = ~n14;
  assign n343 = ~n60;
  assign n231 = ~n55;
  assign n371 = ~n31;
  assign n370 = ~n2;
  assign n364 = ~n57;
  assign n365 = ~n16;
  assign n357 = ~n62;
  assign n359 = ~n42;
  assign n341 = ~n58;
  assign n269 = ~n26;
  assign n344 = ~n34;
  assign n252 = ~n12;
  assign n291 = ~n23;
  assign n242 = ~n25;
  assign n275 = ~n30;
  assign n263 = ~n1;
  assign n338 = ~n46;
  assign n337 = ~n48;
  assign n199 = ~n8;
  assign n334 = ~n22;
  assign n333 = ~n32;
  assign n368 = ~n18;
  assign n360 = ~n11;
  assign n339 = ~n21;
  assign n362 = ~n13;
  assign n340 = ~n47;
  assign n335 = ~n61;
  assign n358 = ~n37;
  assign n374 = ~n29;
  assign n351 = ~n35;
  assign n349 = ~n53;
  assign n356 = ~n43;
  assign n292 = n333 & n0;
  assign n290 = n334 & n54;
  assign n293 = n335 & n29;
  assign n220 = n336 & n41;
  assign n294 = n337 & n16;
  assign n299 = n338 & n14;
  assign n298 = n339 & n53;
  assign n297 = n340 & n15;
  assign n301 = n341 & n26;
  assign n295 = n342 & n47;
  assign n302 = n343 & n28;
  assign n303 = n344 & n2;
  assign n304 = n345 & n22;
  assign n305 = n346 & n13;
  assign n296 = n347 & n52;
  assign n306 = n348 & n6;
  assign n307 = n349 & n21;
  assign n308 = n350 & n12;
  assign n309 = n351 & n3;
  assign n310 = n352 & n59;
  assign n311 = n353 & n35;
  assign n312 = n354 & n18;
  assign n313 = n355 & n20;
  assign n314 = n356 & n11;
  assign n316 = n357 & n30;
  assign n317 = n358 & n5;
  assign n318 = n359 & n10;
  assign n319 = n360 & n43;
  assign n320 = n361 & n17;
  assign n300 = n362 & n45;
  assign n321 = n363 & n9;
  assign n322 = n364 & n25;
  assign n323 = n365 & n48;
  assign n324 = n366 & n7;
  assign n325 = n367 & n49;
  assign n288 = n368 & n50;
  assign n315 = n369 & n39;
  assign n326 = n370 & n34;
  assign n328 = n231 & n23;
  assign n329 = n371 & n63;
  assign n330 = n372 & n27;
  assign n331 = n373 & n31;
  assign n332 = n229 & n19;
  assign n327 = n374 & n61;
  assign n284 = n288 & n289;
  assign n286 = n290 & n291;
  assign n287 = n292 & n1;
  assign n285 = ~n290;
  assign n272 = ~n293;
  assign n77 = ~n294;
  assign n186 = ~n295;
  assign n279 = ~n296;
  assign n280 = ~n297;
  assign n278 = ~n298;
  assign n282 = ~n299;
  assign n188 = ~n300;
  assign n257 = ~n301;
  assign n273 = ~n302;
  assign n140 = ~n303;
  assign n233 = ~n304;
  assign n251 = ~n305;
  assign n268 = ~n306;
  assign n254 = ~n307;
  assign n255 = ~n308;
  assign n109 = ~n309;
  assign n133 = ~n310;
  assign n262 = ~n292;
  assign n103 = ~n311;
  assign n239 = ~n312;
  assign n197 = ~n313;
  assign n258 = ~n314;
  assign n135 = ~n315;
  assign n277 = ~n316;
  assign n240 = ~n317;
  assign n261 = ~n318;
  assign n154 = ~n319;
  assign n271 = ~n320;
  assign n260 = ~n321;
  assign n235 = ~n322;
  assign n265 = ~n323;
  assign n266 = ~n324;
  assign n264 = ~n325;
  assign n283 = ~n288;
  assign n126 = ~n326;
  assign n184 = ~n327;
  assign n253 = ~n328;
  assign n274 = ~n329;
  assign n256 = ~n330;
  assign n124 = ~n331;
  assign n270 = ~n332;
  assign n243 = n251 & n252;
  assign n232 = n253 & n254;
  assign n244 = n251 & n255;
  assign n234 = n256 & n257;
  assign n245 = n258 & n259;
  assign n223 = n260 & n199;
  assign n219 = n258 & n261;
  assign n246 = n262 & n263;
  assign n247 = n264 & n265;
  assign n224 = n266 & n267;
  assign n236 = n266 & n268;
  assign n222 = n256 & n269;
  assign n238 = n270 & n271;
  assign n218 = n272 & n273;
  assign n225 = n274 & n275;
  assign n226 = n272 & n276;
  assign n142 = n274 & n277;
  assign n248 = n278 & n279;
  assign n227 = n280 & n281;
  assign n144 = n280 & n282;
  assign n249 = n283 & n19;
  assign n221 = n260 & n40;
  assign n228 = ~n284;
  assign n250 = n285 & n23;
  assign n230 = ~n286;
  assign n241 = ~n287;
  assign n113 = n142 & n218;
  assign n206 = n219 & n220;
  assign n198 = n219 & n221;
  assign n207 = n222 & n58;
  assign n208 = n219 & n223;
  assign n209 = n224 & n38;
  assign n210 = n225 & n62;
  assign n211 = n226 & n60;
  assign n212 = n227 & n46;
  assign n213 = n228 & n229;
  assign n214 = n230 & n231;
  assign n196 = n232 & n233;
  assign n201 = n234 & n235;
  assign n204 = n236 & n237;
  assign n75 = n238 & n239;
  assign n202 = n236 & n240;
  assign n215 = n241 & n33;
  assign n205 = n234 & n242;
  assign n216 = n243 & n44;
  assign n85 = n144 & n244;
  assign n217 = n245 & n42;
  assign n180 = ~n246;
  assign n200 = ~n247;
  assign n203 = ~n248;
  assign n176 = ~n249;
  assign n182 = ~n250;
  assign n73 = n196 & n197;
  assign n189 = n198 & n199;
  assign n190 = n75 & n200;
  assign n191 = n201 & n164;
  assign n192 = n202 & n166;
  assign n193 = n196 & n203;
  assign n163 = n201 & n56;
  assign n194 = n204 & n37;
  assign n165 = n202 & n36;
  assign n195 = n205 & n57;
  assign n173 = ~n206;
  assign n177 = ~n198;
  assign n156 = ~n207;
  assign n178 = ~n208;
  assign n158 = ~n209;
  assign n115 = ~n210;
  assign n183 = ~n211;
  assign n185 = ~n212;
  assign n175 = ~n213;
  assign n181 = ~n214;
  assign n179 = ~n215;
  assign n187 = ~n216;
  assign n174 = ~n217;
  assign n151 = n163 & n164;
  assign n152 = n165 & n166;
  assign n137 = n173 & n174;
  assign n167 = n175 & n176;
  assign n168 = n177 & n178;
  assign n169 = n179 & n180;
  assign n170 = n181 & n182;
  assign n171 = n183 & n184;
  assign n80 = n185 & n186;
  assign n172 = n187 & n188;
  assign n153 = ~n189;
  assign n146 = ~n190;
  assign n160 = ~n191;
  assign n162 = ~n192;
  assign n149 = ~n193;
  assign n159 = ~n163;
  assign n157 = ~n194;
  assign n161 = ~n165;
  assign n155 = ~n195;
  assign n132 = ~n151;
  assign n134 = ~n152;
  assign n136 = n153 & n154;
  assign n120 = n155 & n156;
  assign n122 = n157 & n158;
  assign n147 = n159 & n160;
  assign n150 = n161 & n162;
  assign n145 = ~n167;
  assign n91 = ~n168;
  assign n139 = ~n169;
  assign n148 = ~n170;
  assign n141 = ~n171;
  assign n143 = ~n172;
  assign n119 = n132 & n133;
  assign n121 = n134 & n135;
  assign n88 = n136 & n137;
  assign n129 = n139 & n140;
  assign n130 = n141 & n142;
  assign n131 = n143 & n144;
  assign n138 = n145 & n146;
  assign n128 = ~n147;
  assign n111 = n148 & n149;
  assign n99 = ~n150;
  assign n116 = n119 & n120;
  assign n94 = n121 & n122;
  assign n71 = n128 & n113;
  assign n125 = ~n129;
  assign n123 = ~n130;
  assign n82 = ~n131;
  assign n127 = ~n138;
  assign n112 = ~n116;
  assign n114 = n123 & n124;
  assign n117 = n125 & n126;
  assign n118 = n127 & n73;
  assign n106 = n112 & n113;
  assign n68 = n114 & n115;
  assign n108 = ~n117;
  assign n110 = ~n118;
  assign n97 = ~n106;
  assign n107 = n108 & n109;
  assign n105 = n110 & n111;
  assign n104 = ~n105;
  assign n102 = ~n107;
  assign n100 = n102 & n103;
  assign n101 = n104 & n71;
  assign n98 = ~n100;
  assign n96 = ~n101;
  assign n66 = n96 & n97;
  assign n95 = n98 & n99;
  assign n93 = ~n95;
  assign n92 = n93 & n94;
  assign n90 = ~n92;
  assign n89 = n90 & n91;
  assign n87 = ~n89;
  assign n86 = n87 & n88;
  assign n84 = ~n86;
  assign n83 = n84 & n85;
  assign n81 = ~n83;
  assign n79 = n81 & n82;
  assign n78 = n79 & n80;
  assign n76 = ~n78;
  assign n74 = n76 & n77;
  assign n72 = n74 & n75;
  assign n70 = n72 & n73;
  assign n69 = n70 & n71;
  assign n67 = ~n69;
  assign n65 = n67 & n68;
  assign n64 = n65 & n66;
  assign n375 = ~n64;
endmodule
