module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63;
  output y0;
  wire n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254;
  assign n65 = x29 & ~x61;
  assign n66 = x28 & ~x60;
  assign n67 = ~n65 & ~n66;
  assign n68 = x30 & ~x62;
  assign n69 = x31 & ~x63;
  assign n70 = ~n68 & ~n69;
  assign n71 = n67 & n70;
  assign n72 = ~x27 & x59;
  assign n73 = x25 & ~x57;
  assign n74 = x26 & ~x58;
  assign n75 = x27 & ~x59;
  assign n76 = ~n74 & ~n75;
  assign n77 = ~n73 & n76;
  assign n78 = x56 & n77;
  assign n79 = ~x24 & n78;
  assign n80 = ~n72 & ~n79;
  assign n81 = x58 ^ x26;
  assign n82 = n81 ^ n75;
  assign n83 = x57 ^ x25;
  assign n84 = x57 & ~n83;
  assign n85 = n84 ^ x26;
  assign n86 = n85 ^ x57;
  assign n87 = n82 & ~n86;
  assign n88 = n87 ^ n84;
  assign n89 = n88 ^ x57;
  assign n90 = ~n75 & n89;
  assign n91 = n80 & ~n90;
  assign n92 = n71 & ~n91;
  assign n93 = ~x24 & n77;
  assign n94 = ~n78 & ~n93;
  assign n95 = n71 & ~n94;
  assign n96 = ~x21 & x53;
  assign n97 = ~x20 & x52;
  assign n98 = ~n96 & ~n97;
  assign n99 = x22 & ~x54;
  assign n100 = x21 & ~x53;
  assign n101 = x23 & ~x55;
  assign n102 = ~n100 & ~n101;
  assign n103 = ~n99 & n102;
  assign n104 = ~n98 & n103;
  assign n105 = x55 ^ x23;
  assign n106 = ~x22 & x54;
  assign n107 = n106 ^ x55;
  assign n108 = ~n105 & ~n107;
  assign n109 = n108 ^ x23;
  assign n110 = ~n104 & n109;
  assign n111 = x20 & ~x52;
  assign n112 = n103 & ~n111;
  assign n113 = ~x16 & x48;
  assign n114 = ~x17 & x49;
  assign n115 = ~n113 & ~n114;
  assign n116 = x18 & ~x50;
  assign n117 = x17 & ~x49;
  assign n118 = x19 & ~x51;
  assign n119 = ~n117 & ~n118;
  assign n120 = ~n116 & n119;
  assign n121 = ~n115 & n120;
  assign n122 = x51 ^ x19;
  assign n123 = ~x18 & x50;
  assign n124 = n123 ^ x51;
  assign n125 = ~n122 & ~n124;
  assign n126 = n125 ^ x19;
  assign n127 = ~n121 & n126;
  assign n128 = n112 & ~n127;
  assign n129 = n110 & ~n128;
  assign n130 = n95 & ~n129;
  assign n131 = ~n92 & ~n130;
  assign n132 = ~x30 & ~n69;
  assign n133 = x62 & n132;
  assign n134 = x63 ^ x31;
  assign n135 = x61 ^ x29;
  assign n136 = x61 ^ x28;
  assign n137 = n136 ^ x61;
  assign n138 = x61 ^ x60;
  assign n139 = n138 ^ x61;
  assign n140 = ~n137 & n139;
  assign n141 = n140 ^ x61;
  assign n142 = ~n135 & ~n141;
  assign n143 = n142 ^ x29;
  assign n144 = n143 ^ x63;
  assign n145 = n144 ^ x63;
  assign n146 = n68 ^ x63;
  assign n147 = n146 ^ x63;
  assign n148 = ~n145 & ~n147;
  assign n149 = n148 ^ x63;
  assign n150 = ~n134 & ~n149;
  assign n151 = n150 ^ x31;
  assign n152 = ~n133 & n151;
  assign n153 = x16 & ~x48;
  assign n154 = x47 ^ x15;
  assign n155 = x47 ^ x14;
  assign n156 = n155 ^ x47;
  assign n157 = x47 ^ x46;
  assign n158 = n157 ^ x47;
  assign n159 = ~n156 & n158;
  assign n160 = n159 ^ x47;
  assign n161 = ~n154 & ~n160;
  assign n162 = n161 ^ x15;
  assign n163 = x45 ^ x13;
  assign n164 = x45 ^ x12;
  assign n165 = n164 ^ x45;
  assign n166 = x45 ^ x44;
  assign n167 = n166 ^ x45;
  assign n168 = ~n165 & n167;
  assign n169 = n168 ^ x45;
  assign n170 = ~n163 & ~n169;
  assign n171 = n170 ^ x13;
  assign n232 = x13 & ~x45;
  assign n233 = x12 & ~x44;
  assign n234 = ~n232 & ~n233;
  assign n172 = ~x11 & x43;
  assign n173 = x11 & ~x43;
  assign n174 = x10 & ~x42;
  assign n175 = ~n173 & ~n174;
  assign n176 = x9 & ~x41;
  assign n177 = x40 & ~n176;
  assign n178 = n175 & n177;
  assign n179 = ~x8 & n178;
  assign n180 = ~n172 & ~n179;
  assign n181 = x42 ^ x10;
  assign n182 = ~x9 & x41;
  assign n183 = n182 ^ x42;
  assign n184 = ~n181 & n183;
  assign n185 = n184 ^ x42;
  assign n186 = ~n173 & n185;
  assign n187 = n180 & ~n186;
  assign n188 = ~x8 & ~n176;
  assign n189 = n175 & n188;
  assign n190 = ~n178 & ~n189;
  assign n191 = ~x7 & x39;
  assign n192 = x5 & ~x37;
  assign n193 = x6 & ~x38;
  assign n194 = x7 & ~x39;
  assign n195 = ~n193 & ~n194;
  assign n196 = ~n192 & n195;
  assign n197 = x36 & n196;
  assign n198 = ~x4 & n197;
  assign n199 = ~n191 & ~n198;
  assign n200 = x38 ^ x6;
  assign n201 = n200 ^ n194;
  assign n202 = x37 ^ x5;
  assign n203 = x37 & ~n202;
  assign n204 = n203 ^ x6;
  assign n205 = n204 ^ x37;
  assign n206 = n201 & ~n205;
  assign n207 = n206 ^ n203;
  assign n208 = n207 ^ x37;
  assign n209 = ~n194 & n208;
  assign n210 = n199 & ~n209;
  assign n211 = ~x4 & n196;
  assign n212 = ~n197 & ~n211;
  assign n213 = x35 ^ x3;
  assign n214 = x34 ^ x2;
  assign n217 = x34 ^ x1;
  assign n215 = x0 & ~x32;
  assign n216 = n215 ^ x34;
  assign n218 = n217 ^ n216;
  assign n219 = x34 ^ x33;
  assign n220 = n219 ^ n217;
  assign n221 = n218 & ~n220;
  assign n222 = n221 ^ n217;
  assign n223 = ~n214 & n222;
  assign n224 = n223 ^ x2;
  assign n225 = n224 ^ x35;
  assign n226 = ~n213 & n225;
  assign n227 = n226 ^ x3;
  assign n228 = ~n212 & ~n227;
  assign n229 = n210 & ~n228;
  assign n230 = ~n190 & ~n229;
  assign n231 = n187 & ~n230;
  assign n235 = n234 ^ n231;
  assign n236 = x14 & ~x46;
  assign n237 = x15 & ~x47;
  assign n238 = ~n236 & ~n237;
  assign n239 = n238 ^ n231;
  assign n240 = ~n231 & ~n239;
  assign n241 = n240 ^ n231;
  assign n242 = ~n235 & ~n241;
  assign n243 = n242 ^ n240;
  assign n244 = n243 ^ n231;
  assign n245 = n244 ^ n238;
  assign n246 = n171 & ~n245;
  assign n247 = n246 ^ n238;
  assign n248 = n162 & ~n247;
  assign n249 = ~n153 & ~n248;
  assign n250 = n120 & n249;
  assign n251 = n112 & n250;
  assign n252 = n95 & n251;
  assign n253 = n152 & ~n252;
  assign n254 = n131 & n253;
  assign y0 = ~n254;
endmodule
