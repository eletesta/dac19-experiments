module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700, x701, x702, x703, x704, x705, x706, x707, x708, x709, x710, x711, x712, x713, x714, x715, x716, x717, x718, x719, x720, x721, x722, x723, x724, x725, x726, x727, x728, x729, x730, x731, x732, x733, x734, x735, x736, x737, x738, x739, x740, x741, x742, x743, x744, x745, x746, x747, x748, x749, x750, x751, x752, x753, x754, x755, x756, x757, x758, x759, x760, x761, x762, x763, x764, x765, x766, x767, x768, x769, x770, x771, x772, x773, x774, x775, x776, x777, x778, x779, x780, x781, x782, x783, x784, x785, x786, x787, x788, x789, x790, x791, x792, x793, x794, x795, x796, x797, x798, x799, x800, x801, x802, x803, x804, x805, x806, x807, x808, x809, x810, x811, x812, x813, x814, x815, x816, x817, x818, x819, x820, x821, x822, x823, x824, x825, x826, x827, x828, x829, x830, x831, x832, x833, x834, x835, x836, x837, x838, x839, x840, x841, x842, x843, x844, x845, x846, x847, x848, x849, x850, x851, x852, x853, x854, x855, x856, x857, x858, x859, x860, x861, x862, x863, x864, x865, x866, x867, x868, x869, x870, x871, x872, x873, x874, x875, x876, x877, x878, x879, x880, x881, x882, x883, x884, x885, x886, x887, x888, x889, x890, x891, x892, x893, x894, x895, x896, x897, x898, x899, x900, x901, x902, x903, x904, x905, x906, x907, x908, x909, x910, x911, x912, x913, x914, x915, x916, x917, x918, x919, x920, x921, x922, x923, x924, x925, x926, x927, x928, x929, x930, x931, x932, x933, x934, x935, x936, x937, x938, x939, x940, x941, x942, x943, x944, x945, x946, x947, x948, x949, x950, x951, x952, x953, x954, x955, x956, x957, x958, x959, x960, x961, x962, x963, x964, x965, x966, x967, x968, x969, x970, x971, x972, x973, x974, x975, x976, x977, x978, x979, x980, x981, x982, x983, x984, x985, x986, x987, x988, x989, x990, x991, x992, x993, x994, x995, x996, x997, x998, x999, x1000, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700, x701, x702, x703, x704, x705, x706, x707, x708, x709, x710, x711, x712, x713, x714, x715, x716, x717, x718, x719, x720, x721, x722, x723, x724, x725, x726, x727, x728, x729, x730, x731, x732, x733, x734, x735, x736, x737, x738, x739, x740, x741, x742, x743, x744, x745, x746, x747, x748, x749, x750, x751, x752, x753, x754, x755, x756, x757, x758, x759, x760, x761, x762, x763, x764, x765, x766, x767, x768, x769, x770, x771, x772, x773, x774, x775, x776, x777, x778, x779, x780, x781, x782, x783, x784, x785, x786, x787, x788, x789, x790, x791, x792, x793, x794, x795, x796, x797, x798, x799, x800, x801, x802, x803, x804, x805, x806, x807, x808, x809, x810, x811, x812, x813, x814, x815, x816, x817, x818, x819, x820, x821, x822, x823, x824, x825, x826, x827, x828, x829, x830, x831, x832, x833, x834, x835, x836, x837, x838, x839, x840, x841, x842, x843, x844, x845, x846, x847, x848, x849, x850, x851, x852, x853, x854, x855, x856, x857, x858, x859, x860, x861, x862, x863, x864, x865, x866, x867, x868, x869, x870, x871, x872, x873, x874, x875, x876, x877, x878, x879, x880, x881, x882, x883, x884, x885, x886, x887, x888, x889, x890, x891, x892, x893, x894, x895, x896, x897, x898, x899, x900, x901, x902, x903, x904, x905, x906, x907, x908, x909, x910, x911, x912, x913, x914, x915, x916, x917, x918, x919, x920, x921, x922, x923, x924, x925, x926, x927, x928, x929, x930, x931, x932, x933, x934, x935, x936, x937, x938, x939, x940, x941, x942, x943, x944, x945, x946, x947, x948, x949, x950, x951, x952, x953, x954, x955, x956, x957, x958, x959, x960, x961, x962, x963, x964, x965, x966, x967, x968, x969, x970, x971, x972, x973, x974, x975, x976, x977, x978, x979, x980, x981, x982, x983, x984, x985, x986, x987, x988, x989, x990, x991, x992, x993, x994, x995, x996, x997, x998, x999, x1000;
  output y0;
  wire n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235;
  assign n2014 = x243 & x244;
  assign n2015 = x245 & x246;
  assign n2023 = n2014 & n2015;
  assign n1867 = x242 ^ x241;
  assign n2016 = ~n2014 & ~n2015;
  assign n2017 = n1867 & ~n2016;
  assign n2018 = ~x243 & ~x244;
  assign n2019 = ~x245 & ~x246;
  assign n2020 = ~n2018 & ~n2019;
  assign n2021 = n2017 & n2020;
  assign n2022 = n2016 & ~n2020;
  assign n2024 = x241 & x242;
  assign n2025 = ~n2023 & n2024;
  assign n2026 = ~n2022 & n2025;
  assign n2027 = ~n2021 & ~n2026;
  assign n2120 = ~n2023 & n2027;
  assign n2036 = x239 & x240;
  assign n2037 = x237 & x238;
  assign n2044 = n2036 & n2037;
  assign n2038 = ~n2036 & ~n2037;
  assign n2039 = ~x239 & ~x240;
  assign n2040 = ~x237 & ~x238;
  assign n2041 = ~n2039 & ~n2040;
  assign n2042 = n2038 & ~n2041;
  assign n2048 = x235 & x236;
  assign n2050 = ~n2044 & n2048;
  assign n2051 = ~n2042 & n2050;
  assign n1872 = x236 ^ x235;
  assign n2052 = n1872 & ~n2038;
  assign n2053 = n2041 & n2052;
  assign n2054 = ~n2051 & ~n2053;
  assign n2121 = ~n2044 & n2054;
  assign n2183 = ~n2120 & ~n2121;
  assign n2059 = x231 & x232;
  assign n2060 = x233 & x234;
  assign n2061 = ~n2059 & ~n2060;
  assign n2062 = ~x231 & ~x232;
  assign n2063 = ~x233 & ~x234;
  assign n2064 = ~n2062 & ~n2063;
  assign n2065 = ~n2061 & n2064;
  assign n2066 = x230 & n2065;
  assign n2067 = n2059 & n2060;
  assign n2068 = ~n2066 & ~n2067;
  assign n2069 = n2061 & ~n2064;
  assign n2073 = ~n2067 & ~n2069;
  assign n2074 = x230 & ~n2073;
  assign n2075 = ~x230 & ~n2065;
  assign n2076 = x229 & ~n2075;
  assign n2077 = ~n2074 & n2076;
  assign n2128 = n2068 & ~n2077;
  assign n2082 = x225 & x226;
  assign n2083 = x227 & x228;
  assign n2084 = ~n2082 & ~n2083;
  assign n2085 = ~x225 & ~x226;
  assign n2086 = ~x227 & ~x228;
  assign n2087 = ~n2085 & ~n2086;
  assign n2088 = ~n2084 & n2087;
  assign n2089 = x224 & n2088;
  assign n2090 = n2082 & n2083;
  assign n2091 = ~n2089 & ~n2090;
  assign n2092 = n2084 & ~n2087;
  assign n2096 = ~n2090 & ~n2092;
  assign n2097 = x224 & ~n2096;
  assign n2098 = ~x224 & ~n2088;
  assign n2099 = x223 & ~n2098;
  assign n2100 = ~n2097 & n2099;
  assign n2127 = n2091 & ~n2100;
  assign n2129 = n2128 ^ n2127;
  assign n2093 = ~x224 & n2092;
  assign n2094 = n2091 & ~n2093;
  assign n2095 = ~x223 & ~n2094;
  assign n1861 = x224 ^ x223;
  assign n2101 = n2085 & n2086;
  assign n2102 = n1861 & n2101;
  assign n2103 = ~n2100 & ~n2102;
  assign n2104 = ~n2095 & n2103;
  assign n2070 = ~x230 & n2069;
  assign n2071 = n2068 & ~n2070;
  assign n2072 = ~x229 & ~n2071;
  assign n1856 = x230 ^ x229;
  assign n2078 = n2062 & n2063;
  assign n2079 = n1856 & n2078;
  assign n2080 = ~n2077 & ~n2079;
  assign n2081 = ~n2072 & n2080;
  assign n2105 = n2104 ^ n2081;
  assign n1855 = x234 ^ x233;
  assign n1857 = n1856 ^ n1855;
  assign n1854 = x232 ^ x231;
  assign n1858 = n1857 ^ n1854;
  assign n1860 = x228 ^ x227;
  assign n1862 = n1861 ^ n1860;
  assign n1859 = x226 ^ x225;
  assign n1863 = n1862 ^ n1859;
  assign n2058 = n1858 & n1863;
  assign n2124 = n2081 ^ n2058;
  assign n2125 = n2105 & ~n2124;
  assign n2126 = n2125 ^ n2104;
  assign n2130 = n2129 ^ n2126;
  assign n2122 = n2121 ^ n2120;
  assign n2043 = ~n1872 & n2042;
  assign n2045 = n2039 & n2040;
  assign n2046 = ~n2044 & ~n2045;
  assign n2047 = ~n2043 & n2046;
  assign n2049 = ~n2047 & ~n2048;
  assign n2055 = ~n2049 & n2054;
  assign n2028 = ~x241 & ~x242;
  assign n2029 = n2022 & n2028;
  assign n2030 = ~x241 & n2023;
  assign n2031 = n2018 & n2019;
  assign n2032 = ~n2024 & n2031;
  assign n2033 = ~n2030 & ~n2032;
  assign n2034 = ~n2029 & n2033;
  assign n2035 = n2027 & n2034;
  assign n2056 = n2055 ^ n2035;
  assign n1866 = x246 ^ x245;
  assign n1868 = n1867 ^ n1866;
  assign n1865 = x244 ^ x243;
  assign n1869 = n1868 ^ n1865;
  assign n1871 = x240 ^ x239;
  assign n1873 = n1872 ^ n1871;
  assign n1870 = x238 ^ x237;
  assign n1874 = n1873 ^ n1870;
  assign n2013 = n1869 & n1874;
  assign n2117 = n2035 ^ n2013;
  assign n2118 = n2056 & ~n2117;
  assign n2119 = n2118 ^ n2055;
  assign n2123 = n2122 ^ n2119;
  assign n2131 = n2130 ^ n2123;
  assign n2106 = n2105 ^ n2058;
  assign n2057 = n2056 ^ n2013;
  assign n2107 = n2106 ^ n2057;
  assign n1864 = n1863 ^ n1858;
  assign n1875 = n1874 ^ n1869;
  assign n1901 = n1864 & n1875;
  assign n2114 = n2057 ^ n1901;
  assign n2115 = n2107 & ~n2114;
  assign n2116 = n2115 ^ n2106;
  assign n2132 = n2131 ^ n2116;
  assign n2181 = ~n2119 & ~n2130;
  assign n2182 = ~n2132 & ~n2181;
  assign n2184 = ~n2182 & ~n2183;
  assign n2185 = ~n2116 & ~n2119;
  assign n2186 = n2120 & n2121;
  assign n2189 = ~n2130 & n2186;
  assign n2190 = ~n2185 & ~n2189;
  assign n2187 = n2130 & ~n2186;
  assign n2188 = ~n2185 & n2187;
  assign n2191 = n2190 ^ n2188;
  assign n2192 = ~n2184 & ~n2191;
  assign n2193 = n2192 ^ n2190;
  assign n2178 = n2128 ^ n2126;
  assign n2179 = ~n2129 & ~n2178;
  assign n2180 = n2179 ^ n2126;
  assign n2194 = n2193 ^ n2180;
  assign n2201 = ~n2183 & n2194;
  assign n2202 = ~n2180 & ~n2182;
  assign n2203 = ~n2201 & ~n2202;
  assign n1987 = x251 & x252;
  assign n1988 = x249 & x250;
  assign n1989 = ~n1987 & ~n1988;
  assign n1990 = ~x251 & ~x252;
  assign n1991 = ~x249 & ~x250;
  assign n1992 = ~n1990 & ~n1991;
  assign n1993 = ~n1989 & n1992;
  assign n1994 = x248 & n1993;
  assign n1995 = n1987 & n1988;
  assign n1996 = ~n1994 & ~n1995;
  assign n1997 = n1989 & ~n1992;
  assign n2001 = ~n1995 & ~n1997;
  assign n2002 = x248 & ~n2001;
  assign n2003 = ~x248 & ~n1993;
  assign n2004 = x247 & ~n2003;
  assign n2005 = ~n2002 & n2004;
  assign n2148 = n1996 & ~n2005;
  assign n1964 = x257 & x258;
  assign n1965 = x255 & x256;
  assign n1966 = ~n1964 & ~n1965;
  assign n1967 = ~x257 & ~x258;
  assign n1968 = ~x255 & ~x256;
  assign n1969 = ~n1967 & ~n1968;
  assign n1970 = ~n1966 & n1969;
  assign n1971 = x254 & n1970;
  assign n1972 = n1964 & n1965;
  assign n1973 = ~n1971 & ~n1972;
  assign n1974 = n1966 & ~n1969;
  assign n1978 = ~n1972 & ~n1974;
  assign n1979 = x254 & ~n1978;
  assign n1980 = ~x254 & ~n1970;
  assign n1981 = x253 & ~n1980;
  assign n1982 = ~n1979 & n1981;
  assign n2147 = n1973 & ~n1982;
  assign n2149 = n2148 ^ n2147;
  assign n1998 = ~x248 & n1997;
  assign n1999 = n1996 & ~n1998;
  assign n2000 = ~x247 & ~n1999;
  assign n1895 = x248 ^ x247;
  assign n2006 = n1990 & n1991;
  assign n2007 = n1895 & n2006;
  assign n2008 = ~n2005 & ~n2007;
  assign n2009 = ~n2000 & n2008;
  assign n1975 = ~x254 & n1974;
  assign n1976 = n1973 & ~n1975;
  assign n1977 = ~x253 & ~n1976;
  assign n1890 = x254 ^ x253;
  assign n1983 = n1967 & n1968;
  assign n1984 = n1890 & n1983;
  assign n1985 = ~n1982 & ~n1984;
  assign n1986 = ~n1977 & n1985;
  assign n2010 = n2009 ^ n1986;
  assign n1889 = x256 ^ x255;
  assign n1891 = n1890 ^ n1889;
  assign n1888 = x258 ^ x257;
  assign n1892 = n1891 ^ n1888;
  assign n1894 = x250 ^ x249;
  assign n1896 = n1895 ^ n1894;
  assign n1893 = x252 ^ x251;
  assign n1897 = n1896 ^ n1893;
  assign n2143 = n1892 & n1897;
  assign n2144 = n2143 ^ n1986;
  assign n2145 = n2010 & ~n2144;
  assign n2146 = n2145 ^ n2009;
  assign n2150 = n2149 ^ n2146;
  assign n1929 = ~x269 & ~x270;
  assign n1930 = ~x267 & ~x268;
  assign n1931 = ~n1929 & ~n1930;
  assign n1932 = x269 & x270;
  assign n1933 = x267 & x268;
  assign n1934 = ~n1932 & ~n1933;
  assign n1935 = n1931 & ~n1934;
  assign n1936 = x266 & n1935;
  assign n1937 = n1932 & n1933;
  assign n1938 = ~n1936 & ~n1937;
  assign n1939 = ~n1931 & n1934;
  assign n1940 = ~x266 & n1939;
  assign n1941 = n1929 & n1930;
  assign n1942 = ~n1940 & ~n1941;
  assign n1943 = n1938 & n1942;
  assign n1944 = ~x265 & ~n1943;
  assign n1884 = x266 ^ x265;
  assign n1945 = n1884 & n1935;
  assign n1946 = x265 & x266;
  assign n1947 = n1933 & n1946;
  assign n1948 = x270 & n1947;
  assign n1949 = n1948 ^ n1946;
  assign n1950 = ~n1939 & n1949;
  assign n1951 = ~n1945 & ~n1950;
  assign n1952 = ~x266 & ~x270;
  assign n1953 = n1930 & n1952;
  assign n1954 = ~n1947 & ~n1953;
  assign n1955 = ~x269 & ~n1954;
  assign n1956 = n1951 & ~n1955;
  assign n1957 = ~n1944 & n1956;
  assign n1903 = x263 & x264;
  assign n1904 = ~x261 & ~x262;
  assign n1905 = ~n1903 & n1904;
  assign n1906 = ~x263 & ~x264;
  assign n1907 = x260 & ~n1906;
  assign n1908 = n1905 & ~n1907;
  assign n1909 = x261 & x262;
  assign n1910 = n1903 & n1909;
  assign n1911 = ~n1908 & ~n1910;
  assign n1912 = ~x259 & ~n1911;
  assign n1879 = x260 ^ x259;
  assign n1878 = x262 ^ x261;
  assign n1880 = n1879 ^ n1878;
  assign n1913 = ~x260 & n1906;
  assign n1914 = ~n1909 & n1913;
  assign n1915 = n1880 & n1914;
  assign n1916 = x259 & x260;
  assign n1917 = n1909 & n1916;
  assign n1918 = ~n1903 & n1917;
  assign n1919 = ~n1915 & ~n1918;
  assign n1920 = ~n1912 & n1919;
  assign n1921 = ~n1903 & ~n1909;
  assign n1922 = n1879 & ~n1904;
  assign n1923 = ~n1921 & n1922;
  assign n1924 = ~n1909 & n1916;
  assign n1925 = ~n1905 & n1924;
  assign n1926 = ~n1923 & ~n1925;
  assign n1927 = ~n1906 & ~n1926;
  assign n1928 = n1920 & ~n1927;
  assign n1958 = n1957 ^ n1928;
  assign n1877 = x264 ^ x263;
  assign n1881 = n1880 ^ n1877;
  assign n1883 = x268 ^ x267;
  assign n1885 = n1884 ^ n1883;
  assign n1882 = x270 ^ x269;
  assign n1886 = n1885 ^ n1882;
  assign n2138 = n1881 & n1886;
  assign n2139 = n1958 & n2138;
  assign n2140 = n1928 & n1957;
  assign n2141 = ~n2139 & ~n2140;
  assign n2171 = n2150 ^ n2141;
  assign n1959 = n1892 ^ n1886;
  assign n1961 = n1959 ^ n1881;
  assign n1962 = ~n1897 & n1961;
  assign n1887 = n1886 ^ n1881;
  assign n1960 = ~n1887 & ~n1959;
  assign n1963 = n1962 ^ n1960;
  assign n2011 = n2010 ^ n1963;
  assign n2012 = n2011 ^ n1958;
  assign n2152 = n2010 & ~n2143;
  assign n2153 = ~n2012 & ~n2152;
  assign n1898 = n1897 ^ n1892;
  assign n2154 = ~n1881 & ~n1886;
  assign n2155 = n1898 & ~n2154;
  assign n2156 = ~n2138 & ~n2155;
  assign n2157 = n2156 ^ n2138;
  assign n2158 = ~n1958 & n2157;
  assign n2159 = n2158 ^ n2138;
  assign n2160 = ~n2153 & ~n2159;
  assign n2172 = n2160 ^ n2150;
  assign n2173 = n2171 & n2172;
  assign n2174 = n2173 ^ n2160;
  assign n2168 = n2148 ^ n2146;
  assign n2169 = ~n2149 & ~n2168;
  assign n2170 = n2169 ^ n2146;
  assign n2175 = n2174 ^ n2170;
  assign n2135 = ~n1910 & ~n1917;
  assign n2136 = ~n1927 & n2135;
  assign n2134 = n1938 & n1951;
  assign n2137 = n2136 ^ n2134;
  assign n2142 = n2141 ^ n2137;
  assign n2151 = n2150 ^ n2142;
  assign n2161 = n2160 ^ n2151;
  assign n2165 = n2161 ^ n2134;
  assign n2166 = n2137 & n2165;
  assign n2167 = n2166 ^ n2136;
  assign n2198 = n2170 ^ n2167;
  assign n2199 = n2175 & n2198;
  assign n2200 = n2199 ^ n2174;
  assign n2204 = n2203 ^ n2200;
  assign n2176 = n2175 ^ n2167;
  assign n1876 = n1875 ^ n1864;
  assign n1899 = n1898 ^ n1887;
  assign n1900 = n1876 & n1899;
  assign n2108 = n2107 ^ n2012;
  assign n1902 = ~n1900 & ~n1901;
  assign n2109 = n2108 ^ n1902;
  assign n2110 = ~n1900 & n2109;
  assign n2111 = ~n1901 & n2107;
  assign n2112 = n2012 & ~n2111;
  assign n2113 = ~n2110 & ~n2112;
  assign n2133 = n2132 ^ n2113;
  assign n2162 = n2161 ^ n2113;
  assign n2163 = n2133 & n2162;
  assign n2164 = n2163 ^ n2132;
  assign n2177 = n2176 ^ n2164;
  assign n2195 = n2194 ^ n2164;
  assign n2196 = n2177 & n2195;
  assign n2197 = n2196 ^ n2194;
  assign n2205 = n2204 ^ n2197;
  assign n2453 = ~x189 & ~x190;
  assign n2454 = ~x191 & ~x192;
  assign n2455 = ~n2453 & ~n2454;
  assign n2456 = x189 & x190;
  assign n2457 = x191 & x192;
  assign n2458 = ~n2456 & ~n2457;
  assign n2459 = n2455 & ~n2458;
  assign n2460 = x188 & n2459;
  assign n2461 = n2456 & n2457;
  assign n2462 = ~n2460 & ~n2461;
  assign n2469 = ~x188 & n2459;
  assign n2463 = ~n2455 & n2458;
  assign n2470 = x192 & n2456;
  assign n2471 = x188 & ~n2470;
  assign n2472 = ~n2463 & n2471;
  assign n2473 = ~n2469 & ~n2472;
  assign n2474 = x187 & ~n2473;
  assign n2530 = n2462 & ~n2474;
  assign n2436 = x197 & x198;
  assign n2437 = x195 & x196;
  assign n2441 = n2436 & n2437;
  assign n2433 = ~x197 & ~x198;
  assign n2434 = ~x195 & ~x196;
  assign n2435 = ~n2433 & ~n2434;
  assign n2357 = x194 ^ x193;
  assign n2438 = ~n2436 & ~n2437;
  assign n2447 = n2357 & ~n2438;
  assign n2448 = n2435 & n2447;
  assign n2439 = ~n2435 & n2438;
  assign n2445 = x193 & x194;
  assign n2449 = ~n2441 & n2445;
  assign n2450 = ~n2439 & n2449;
  assign n2451 = ~n2448 & ~n2450;
  assign n2529 = ~n2441 & n2451;
  assign n2531 = n2530 ^ n2529;
  assign n2464 = ~x188 & n2463;
  assign n2465 = n2453 & n2454;
  assign n2466 = ~n2464 & ~n2465;
  assign n2467 = n2462 & n2466;
  assign n2468 = ~x187 & ~n2467;
  assign n2475 = x187 & x188;
  assign n2476 = n2456 & n2475;
  assign n2477 = ~x188 & ~x192;
  assign n2478 = n2453 & n2477;
  assign n2479 = ~n2476 & ~n2478;
  assign n2480 = ~x191 & ~n2479;
  assign n2481 = ~n2474 & ~n2480;
  assign n2482 = ~n2468 & n2481;
  assign n2440 = ~n2357 & n2439;
  assign n2442 = n2433 & n2434;
  assign n2443 = ~n2441 & ~n2442;
  assign n2444 = ~n2440 & n2443;
  assign n2446 = ~n2444 & ~n2445;
  assign n2452 = ~n2446 & n2451;
  assign n2483 = n2482 ^ n2452;
  assign n2352 = x190 ^ x189;
  assign n2351 = x192 ^ x191;
  assign n2353 = n2352 ^ n2351;
  assign n2350 = x188 ^ x187;
  assign n2354 = n2353 ^ n2350;
  assign n2356 = x198 ^ x197;
  assign n2358 = n2357 ^ n2356;
  assign n2355 = x196 ^ x195;
  assign n2359 = n2358 ^ n2355;
  assign n2432 = n2354 & n2359;
  assign n2526 = n2452 ^ n2432;
  assign n2527 = n2483 & ~n2526;
  assign n2528 = n2527 ^ n2482;
  assign n2532 = n2531 ^ n2528;
  assign n2378 = x179 & x180;
  assign n2379 = x177 & x178;
  assign n2380 = ~n2378 & ~n2379;
  assign n2381 = ~x179 & ~x180;
  assign n2382 = ~x177 & ~x178;
  assign n2383 = ~n2381 & ~n2382;
  assign n2384 = ~n2380 & n2383;
  assign n2385 = x176 & n2384;
  assign n2386 = n2378 & n2379;
  assign n2387 = ~n2385 & ~n2386;
  assign n2388 = n2380 & ~n2383;
  assign n2392 = ~n2386 & ~n2388;
  assign n2393 = x176 & ~n2392;
  assign n2394 = ~x176 & ~n2384;
  assign n2395 = x175 & ~n2394;
  assign n2396 = ~n2393 & n2395;
  assign n2523 = n2387 & ~n2396;
  assign n2401 = ~x185 & ~x186;
  assign n2402 = ~x183 & ~x184;
  assign n2403 = ~n2401 & ~n2402;
  assign n2404 = x185 & x186;
  assign n2405 = x183 & x184;
  assign n2406 = ~n2404 & ~n2405;
  assign n2407 = n2403 & ~n2406;
  assign n2408 = x182 & n2407;
  assign n2409 = n2404 & n2405;
  assign n2410 = ~n2408 & ~n2409;
  assign n2368 = x182 ^ x181;
  assign n2417 = n2368 & n2407;
  assign n2411 = ~n2403 & n2406;
  assign n2418 = x181 & x182;
  assign n2419 = n2405 & n2418;
  assign n2420 = x186 & n2419;
  assign n2421 = n2420 ^ n2418;
  assign n2422 = ~n2411 & n2421;
  assign n2423 = ~n2417 & ~n2422;
  assign n2522 = n2410 & n2423;
  assign n2524 = n2523 ^ n2522;
  assign n2412 = ~x182 & n2411;
  assign n2413 = n2401 & n2402;
  assign n2414 = ~n2412 & ~n2413;
  assign n2415 = n2410 & n2414;
  assign n2416 = ~x181 & ~n2415;
  assign n2424 = ~x182 & ~x186;
  assign n2425 = n2402 & n2424;
  assign n2426 = ~n2419 & ~n2425;
  assign n2427 = ~x185 & ~n2426;
  assign n2428 = n2423 & ~n2427;
  assign n2429 = ~n2416 & n2428;
  assign n2389 = ~x176 & n2388;
  assign n2390 = n2387 & ~n2389;
  assign n2391 = ~x175 & ~n2390;
  assign n2363 = x176 ^ x175;
  assign n2397 = n2381 & n2382;
  assign n2398 = n2363 & n2397;
  assign n2399 = ~n2396 & ~n2398;
  assign n2400 = ~n2391 & n2399;
  assign n2430 = n2429 ^ n2400;
  assign n2362 = x178 ^ x177;
  assign n2364 = n2363 ^ n2362;
  assign n2361 = x180 ^ x179;
  assign n2365 = n2364 ^ n2361;
  assign n2367 = x184 ^ x183;
  assign n2369 = n2368 ^ n2367;
  assign n2366 = x186 ^ x185;
  assign n2370 = n2369 ^ n2366;
  assign n2377 = n2365 & n2370;
  assign n2519 = n2400 ^ n2377;
  assign n2520 = n2430 & ~n2519;
  assign n2521 = n2520 ^ n2429;
  assign n2525 = n2524 ^ n2521;
  assign n2533 = n2532 ^ n2525;
  assign n2484 = n2483 ^ n2432;
  assign n2431 = n2430 ^ n2377;
  assign n2485 = n2484 ^ n2431;
  assign n2360 = n2359 ^ n2354;
  assign n2371 = n2370 ^ n2365;
  assign n2488 = n2360 & n2371;
  assign n2516 = n2488 ^ n2431;
  assign n2517 = n2485 & ~n2516;
  assign n2518 = n2517 ^ n2484;
  assign n2534 = n2533 ^ n2518;
  assign n2557 = ~n2518 & n2522;
  assign n2558 = ~n2534 & ~n2557;
  assign n2559 = n2518 & ~n2522;
  assign n2560 = n2523 ^ n2521;
  assign n2561 = n2532 ^ n2521;
  assign n2562 = n2560 & n2561;
  assign n2563 = n2562 ^ n2532;
  assign n2564 = ~n2559 & ~n2563;
  assign n2565 = ~n2558 & n2564;
  assign n2566 = n2558 & n2563;
  assign n2567 = ~n2565 & ~n2566;
  assign n2554 = n2530 ^ n2528;
  assign n2555 = ~n2531 & ~n2554;
  assign n2556 = n2555 ^ n2528;
  assign n2568 = n2567 ^ n2556;
  assign n2273 = x206 ^ x205;
  assign n2297 = ~x209 & ~x210;
  assign n2302 = n2273 & ~n2297;
  assign n2272 = x208 ^ x207;
  assign n2290 = x209 & x210;
  assign n2304 = n2290 ^ x208;
  assign n2305 = n2272 & ~n2304;
  assign n2306 = n2305 ^ x207;
  assign n2307 = n2302 & n2306;
  assign n2292 = x207 & x208;
  assign n2291 = ~x207 & ~x208;
  assign n2293 = n2292 ^ n2291;
  assign n2294 = ~n2290 & n2293;
  assign n2295 = n2294 ^ n2292;
  assign n2298 = ~n2292 & n2297;
  assign n2308 = x205 & x206;
  assign n2309 = ~n2298 & n2308;
  assign n2310 = ~n2295 & n2309;
  assign n2311 = ~n2307 & ~n2310;
  assign n2493 = n2290 & n2292;
  assign n2494 = n2311 & ~n2493;
  assign n2313 = ~x203 & ~x204;
  assign n2314 = x200 & ~n2313;
  assign n2315 = x203 & x204;
  assign n2316 = x201 & x202;
  assign n2317 = n2315 & n2316;
  assign n2318 = ~n2314 & ~n2317;
  assign n2277 = x202 ^ x201;
  assign n2319 = n2315 ^ x202;
  assign n2320 = n2277 & ~n2319;
  assign n2321 = n2320 ^ x201;
  assign n2322 = ~n2318 & n2321;
  assign n2323 = ~x201 & ~x202;
  assign n2324 = ~n2315 & n2323;
  assign n2325 = ~n2314 & n2324;
  assign n2326 = ~n2322 & ~n2325;
  assign n2327 = ~x199 & ~n2326;
  assign n2328 = x199 & ~n2313;
  assign n2329 = n2321 & n2328;
  assign n2330 = x199 & x200;
  assign n2331 = ~n2329 & ~n2330;
  assign n2332 = ~n2313 & ~n2316;
  assign n2333 = ~n2324 & n2332;
  assign n2334 = ~x204 & n2316;
  assign n2335 = x200 & ~n2334;
  assign n2336 = ~n2333 & n2335;
  assign n2337 = ~n2331 & ~n2336;
  assign n2338 = ~n2327 & ~n2337;
  assign n2339 = x199 & ~n2323;
  assign n2340 = ~x200 & ~x204;
  assign n2341 = ~n2316 & n2340;
  assign n2342 = ~n2339 & n2341;
  assign n2343 = n2316 & n2330;
  assign n2344 = ~n2342 & ~n2343;
  assign n2345 = ~x203 & ~n2344;
  assign n2346 = n2338 & ~n2345;
  assign n2296 = ~x205 & n2295;
  assign n2274 = n2273 ^ n2272;
  assign n2299 = ~x206 & n2298;
  assign n2300 = n2274 & n2299;
  assign n2301 = ~n2296 & ~n2300;
  assign n2303 = ~n2301 & ~n2302;
  assign n2312 = ~n2303 & n2311;
  assign n2347 = n2346 ^ n2312;
  assign n2263 = x216 ^ x215;
  assign n2256 = x212 ^ x211;
  assign n2264 = n2263 ^ n2256;
  assign n2262 = x214 ^ x213;
  assign n2265 = n2264 ^ n2262;
  assign n2267 = x222 ^ x221;
  assign n2223 = x218 ^ x217;
  assign n2268 = n2267 ^ n2223;
  assign n2266 = x220 ^ x219;
  assign n2269 = n2268 ^ n2266;
  assign n2270 = n2265 & n2269;
  assign n2271 = x210 ^ x209;
  assign n2275 = n2274 ^ n2271;
  assign n2278 = x204 ^ x203;
  assign n2279 = n2278 ^ n2277;
  assign n2276 = x200 ^ x199;
  assign n2280 = n2279 ^ n2276;
  assign n2286 = n2275 & n2280;
  assign n2281 = n2280 ^ n2275;
  assign n2282 = n2269 ^ n2265;
  assign n2283 = n2282 ^ n2280;
  assign n2284 = ~n2281 & n2283;
  assign n2285 = n2284 ^ n2282;
  assign n2287 = n2286 ^ n2285;
  assign n2288 = ~n2270 & ~n2287;
  assign n2289 = n2288 ^ n2286;
  assign n2348 = n2347 ^ n2289;
  assign n2237 = x213 & x214;
  assign n2238 = x215 & x216;
  assign n2239 = ~n2237 & ~n2238;
  assign n2240 = ~x213 & ~x214;
  assign n2241 = ~x215 & ~x216;
  assign n2242 = ~n2240 & ~n2241;
  assign n2243 = ~n2239 & n2242;
  assign n2244 = x212 & n2243;
  assign n2245 = n2237 & n2238;
  assign n2246 = ~n2244 & ~n2245;
  assign n2247 = n2239 & ~n2242;
  assign n2248 = ~x212 & n2247;
  assign n2249 = n2246 & ~n2248;
  assign n2250 = ~x211 & ~n2249;
  assign n2251 = ~n2245 & ~n2247;
  assign n2252 = x212 & ~n2251;
  assign n2253 = ~x212 & ~n2243;
  assign n2254 = x211 & ~n2253;
  assign n2255 = ~n2252 & n2254;
  assign n2257 = n2240 & n2241;
  assign n2258 = n2256 & n2257;
  assign n2259 = ~n2255 & ~n2258;
  assign n2260 = ~n2250 & n2259;
  assign n2207 = x221 & x222;
  assign n2208 = x219 & x220;
  assign n2209 = ~n2207 & ~n2208;
  assign n2210 = ~x221 & ~x222;
  assign n2211 = ~x219 & ~x220;
  assign n2212 = ~n2210 & ~n2211;
  assign n2213 = ~n2209 & n2212;
  assign n2214 = x218 & n2213;
  assign n2215 = n2207 & n2208;
  assign n2216 = ~n2214 & ~n2215;
  assign n2217 = n2209 & ~n2212;
  assign n2218 = ~x218 & n2217;
  assign n2219 = n2210 & n2211;
  assign n2220 = ~n2218 & ~n2219;
  assign n2221 = n2216 & n2220;
  assign n2222 = ~x217 & ~n2221;
  assign n2224 = n2213 & n2223;
  assign n2225 = x217 & x218;
  assign n2226 = n2208 & n2225;
  assign n2227 = x222 & n2226;
  assign n2228 = n2227 ^ n2225;
  assign n2229 = ~n2217 & n2228;
  assign n2230 = ~n2224 & ~n2229;
  assign n2231 = ~x218 & ~x222;
  assign n2232 = n2211 & n2231;
  assign n2233 = ~n2226 & ~n2232;
  assign n2234 = ~x221 & ~n2233;
  assign n2235 = n2230 & ~n2234;
  assign n2236 = ~n2222 & n2235;
  assign n2261 = n2260 ^ n2236;
  assign n2349 = n2348 ^ n2261;
  assign n2508 = n2261 & ~n2270;
  assign n2509 = ~n2349 & ~n2508;
  assign n2510 = ~n2287 & ~n2347;
  assign n2511 = n2510 ^ n2286;
  assign n2512 = ~n2509 & ~n2511;
  assign n2504 = n2246 & ~n2255;
  assign n2503 = n2216 & n2230;
  assign n2505 = n2504 ^ n2503;
  assign n2500 = n2270 ^ n2260;
  assign n2501 = ~n2261 & n2500;
  assign n2502 = n2501 ^ n2270;
  assign n2506 = n2505 ^ n2502;
  assign n2496 = n2286 & n2347;
  assign n2497 = n2312 & n2346;
  assign n2498 = ~n2496 & ~n2497;
  assign n2495 = ~n2322 & ~n2337;
  assign n2499 = n2498 ^ n2495;
  assign n2507 = n2506 ^ n2499;
  assign n2513 = n2512 ^ n2507;
  assign n2541 = n2494 & n2513;
  assign n2542 = n2512 ^ n2498;
  assign n2543 = ~n2499 & ~n2542;
  assign n2544 = n2543 ^ n2512;
  assign n2545 = n2541 & ~n2544;
  assign n2546 = n2495 & n2498;
  assign n2547 = ~n2506 & n2546;
  assign n2548 = ~n2512 & n2547;
  assign n2549 = ~n2545 & ~n2548;
  assign n2514 = n2513 ^ n2494;
  assign n2550 = n2506 & n2544;
  assign n2551 = n2514 & n2550;
  assign n2552 = n2549 & ~n2551;
  assign n2538 = n2504 ^ n2502;
  assign n2539 = ~n2505 & ~n2538;
  assign n2540 = n2539 ^ n2502;
  assign n2553 = n2552 ^ n2540;
  assign n2569 = n2568 ^ n2553;
  assign n2372 = n2371 ^ n2360;
  assign n2373 = n2282 ^ n2281;
  assign n2374 = n2373 ^ n2360;
  assign n2375 = n2372 & ~n2374;
  assign n2376 = n2375 ^ n2371;
  assign n2486 = n2485 ^ n2376;
  assign n2487 = n2349 & n2486;
  assign n2489 = n2485 & n2488;
  assign n2490 = ~n2376 & ~n2485;
  assign n2491 = ~n2489 & ~n2490;
  assign n2492 = ~n2487 & n2491;
  assign n2515 = n2514 ^ n2492;
  assign n2535 = n2534 ^ n2514;
  assign n2536 = n2515 & ~n2535;
  assign n2537 = n2536 ^ n2534;
  assign n2570 = n2569 ^ n2537;
  assign n2206 = n2194 ^ n2177;
  assign n2571 = n2570 ^ n2206;
  assign n2574 = n2534 ^ n2515;
  assign n2572 = n2161 ^ n2132;
  assign n2573 = n2572 ^ n2113;
  assign n2575 = n2574 ^ n2573;
  assign n2576 = n2486 ^ n2349;
  assign n2577 = n2576 ^ n2109;
  assign n2578 = n2373 ^ n2372;
  assign n2579 = n1899 ^ n1876;
  assign n2580 = n2578 & n2579;
  assign n2581 = ~n2577 & ~n2580;
  assign n2582 = n1899 & n2578;
  assign n2583 = n2581 & ~n2582;
  assign n2584 = ~n1901 & n2576;
  assign n2585 = ~n2583 & ~n2584;
  assign n2586 = n2108 & ~n2585;
  assign n2587 = n2580 ^ n2576;
  assign n2588 = ~n1902 & ~n2108;
  assign n2589 = n2588 ^ n2580;
  assign n2590 = ~n2587 & n2589;
  assign n2591 = n2590 ^ n2576;
  assign n2592 = ~n2586 & ~n2591;
  assign n2593 = n2592 ^ n2574;
  assign n2594 = ~n2575 & ~n2593;
  assign n2595 = n2594 ^ n2592;
  assign n2596 = n2595 ^ n2206;
  assign n2597 = ~n2571 & n2596;
  assign n2598 = n2597 ^ n2570;
  assign n2599 = n2205 & n2598;
  assign n2600 = n2200 ^ n2197;
  assign n2601 = n2204 & ~n2600;
  assign n2602 = n2601 ^ n2203;
  assign n2603 = ~n2599 & ~n2602;
  assign n2604 = ~n2540 & ~n2551;
  assign n2605 = n2549 & ~n2604;
  assign n2606 = ~n2556 & ~n2566;
  assign n2607 = ~n2565 & ~n2606;
  assign n2608 = ~n2605 & ~n2607;
  assign n2609 = n2607 ^ n2605;
  assign n2610 = n2553 ^ n2537;
  assign n2611 = n2569 & ~n2610;
  assign n2612 = n2611 ^ n2568;
  assign n2613 = ~n2609 & n2612;
  assign n2614 = ~n2608 & ~n2613;
  assign n2615 = ~n2603 & n2614;
  assign n2616 = n2605 & n2607;
  assign n2617 = ~n2612 & ~n2616;
  assign n2618 = n2612 ^ n2609;
  assign n2619 = n2618 ^ n2205;
  assign n2620 = n2619 ^ n2598;
  assign n2621 = n2617 & n2620;
  assign n2622 = n2615 & ~n2621;
  assign n2623 = n2203 & n2605;
  assign n2624 = n2200 & n2551;
  assign n2625 = ~n2623 & ~n2624;
  assign n2626 = n2607 & ~n2625;
  assign n2627 = ~n2197 & n2626;
  assign n2628 = n2200 & n2203;
  assign n2629 = n2607 & n2628;
  assign n2630 = n2197 & ~n2629;
  assign n2631 = ~n2616 & ~n2628;
  assign n2632 = n2630 & ~n2631;
  assign n2633 = ~n2627 & ~n2632;
  assign n2634 = n2612 & ~n2633;
  assign n2635 = ~n2622 & ~n2634;
  assign n2636 = n2608 & ~n2612;
  assign n2638 = ~n2599 & n2636;
  assign n2639 = ~n2608 & ~n2617;
  assign n2640 = ~n2205 & ~n2639;
  assign n2641 = ~n2598 & n2640;
  assign n2642 = ~n2638 & ~n2641;
  assign n2637 = n2598 & ~n2636;
  assign n2643 = n2642 ^ n2637;
  assign n2644 = n2602 & ~n2643;
  assign n2645 = n2644 ^ n2642;
  assign n2646 = n2635 & n2645;
  assign n1630 = x171 & x172;
  assign n1631 = x173 & x174;
  assign n1632 = ~n1630 & ~n1631;
  assign n1633 = ~x171 & ~x172;
  assign n1634 = ~x173 & ~x174;
  assign n1635 = ~n1633 & ~n1634;
  assign n1636 = ~n1632 & n1635;
  assign n1637 = x170 & n1636;
  assign n1638 = n1630 & n1631;
  assign n1639 = ~n1637 & ~n1638;
  assign n1646 = ~x170 & n1636;
  assign n1640 = n1632 & ~n1635;
  assign n1647 = x174 & n1630;
  assign n1648 = x170 & ~n1647;
  assign n1649 = ~n1640 & n1648;
  assign n1650 = ~n1646 & ~n1649;
  assign n1651 = x169 & ~n1650;
  assign n1719 = n1639 & ~n1651;
  assign n1613 = x165 & x166;
  assign n1614 = x167 & x168;
  assign n1618 = n1613 & n1614;
  assign n1610 = ~x165 & ~x166;
  assign n1611 = ~x167 & ~x168;
  assign n1612 = ~n1610 & ~n1611;
  assign n1615 = ~n1613 & ~n1614;
  assign n1616 = ~n1612 & n1615;
  assign n1622 = x163 & x164;
  assign n1624 = ~n1618 & n1622;
  assign n1625 = ~n1616 & n1624;
  assign n1388 = x164 ^ x163;
  assign n1626 = n1388 & n1612;
  assign n1627 = ~n1615 & n1626;
  assign n1628 = ~n1625 & ~n1627;
  assign n1718 = ~n1618 & n1628;
  assign n1720 = n1719 ^ n1718;
  assign n1641 = ~x170 & n1640;
  assign n1642 = n1633 & n1634;
  assign n1643 = ~n1641 & ~n1642;
  assign n1644 = n1639 & n1643;
  assign n1645 = ~x169 & ~n1644;
  assign n1652 = x169 & x170;
  assign n1653 = n1630 & n1652;
  assign n1654 = ~x170 & ~x174;
  assign n1655 = n1633 & n1654;
  assign n1656 = ~n1653 & ~n1655;
  assign n1657 = ~x173 & ~n1656;
  assign n1658 = ~n1651 & ~n1657;
  assign n1659 = ~n1645 & n1658;
  assign n1617 = ~n1388 & n1616;
  assign n1619 = n1610 & n1611;
  assign n1620 = ~n1618 & ~n1619;
  assign n1621 = ~n1617 & n1620;
  assign n1623 = ~n1621 & ~n1622;
  assign n1629 = ~n1623 & n1628;
  assign n1660 = n1659 ^ n1629;
  assign n1383 = x172 ^ x171;
  assign n1382 = x174 ^ x173;
  assign n1384 = n1383 ^ n1382;
  assign n1381 = x170 ^ x169;
  assign n1385 = n1384 ^ n1381;
  assign n1387 = x166 ^ x165;
  assign n1389 = n1388 ^ n1387;
  assign n1386 = x168 ^ x167;
  assign n1390 = n1389 ^ n1386;
  assign n1609 = n1385 & n1390;
  assign n1715 = n1629 ^ n1609;
  assign n1716 = n1660 & ~n1715;
  assign n1717 = n1716 ^ n1659;
  assign n1772 = n1719 ^ n1717;
  assign n1773 = ~n1720 & ~n1772;
  assign n1774 = n1773 ^ n1717;
  assign n1349 = x134 ^ x133;
  assign n1348 = x136 ^ x135;
  assign n1503 = x137 & x138;
  assign n1504 = n1503 ^ x136;
  assign n1505 = n1348 & ~n1504;
  assign n1506 = n1505 ^ x135;
  assign n1507 = n1349 & n1506;
  assign n1508 = ~x135 & ~x136;
  assign n1509 = ~n1503 & n1508;
  assign n1510 = x135 & x136;
  assign n1511 = x133 & x134;
  assign n1512 = ~n1510 & n1511;
  assign n1513 = ~n1509 & n1512;
  assign n1514 = ~n1507 & ~n1513;
  assign n1515 = ~x137 & ~x138;
  assign n1516 = ~n1514 & ~n1515;
  assign n1517 = n1510 & n1511;
  assign n1518 = ~x138 & n1517;
  assign n1519 = ~n1516 & ~n1518;
  assign n1520 = x134 & ~n1515;
  assign n1521 = n1503 & n1510;
  assign n1522 = ~n1520 & ~n1521;
  assign n1523 = n1506 & ~n1522;
  assign n1680 = n1519 & ~n1523;
  assign n1354 = x128 ^ x127;
  assign n1352 = x130 ^ x129;
  assign n1470 = x131 & x132;
  assign n1471 = n1470 ^ x130;
  assign n1472 = n1352 & ~n1471;
  assign n1473 = n1472 ^ x129;
  assign n1474 = n1354 & n1473;
  assign n1475 = ~x129 & ~x130;
  assign n1476 = ~n1470 & n1475;
  assign n1477 = x129 & x130;
  assign n1478 = x127 & x128;
  assign n1479 = ~n1477 & n1478;
  assign n1480 = ~n1476 & n1479;
  assign n1481 = ~n1474 & ~n1480;
  assign n1482 = ~x131 & ~x132;
  assign n1483 = ~n1481 & ~n1482;
  assign n1484 = n1477 & n1478;
  assign n1485 = ~x132 & n1484;
  assign n1486 = ~n1483 & ~n1485;
  assign n1487 = x128 & ~n1482;
  assign n1488 = n1470 & n1477;
  assign n1489 = ~n1487 & ~n1488;
  assign n1490 = n1473 & ~n1489;
  assign n1679 = n1486 & ~n1490;
  assign n1681 = n1680 ^ n1679;
  assign n1524 = n1509 & ~n1520;
  assign n1525 = ~n1523 & ~n1524;
  assign n1526 = ~x133 & ~n1525;
  assign n1527 = n1519 & ~n1526;
  assign n1350 = n1349 ^ n1348;
  assign n1528 = ~x134 & ~x138;
  assign n1529 = ~n1510 & n1528;
  assign n1530 = n1350 & n1529;
  assign n1531 = ~n1517 & ~n1530;
  assign n1532 = ~x137 & ~n1531;
  assign n1533 = n1527 & ~n1532;
  assign n1491 = n1476 & ~n1487;
  assign n1492 = ~x128 & ~n1477;
  assign n1493 = n1482 & n1492;
  assign n1494 = ~n1491 & ~n1493;
  assign n1495 = ~n1490 & n1494;
  assign n1496 = ~x127 & ~n1495;
  assign n1497 = ~x128 & ~x132;
  assign n1498 = n1475 & n1497;
  assign n1499 = ~n1484 & ~n1498;
  assign n1500 = ~x131 & ~n1499;
  assign n1501 = ~n1496 & ~n1500;
  assign n1502 = n1486 & n1501;
  assign n1534 = n1533 ^ n1502;
  assign n1347 = x138 ^ x137;
  assign n1351 = n1350 ^ n1347;
  assign n1353 = x132 ^ x131;
  assign n1355 = n1354 ^ n1353;
  assign n1356 = n1355 ^ n1352;
  assign n1675 = n1351 & n1356;
  assign n1676 = n1675 ^ n1502;
  assign n1677 = n1534 & ~n1676;
  assign n1678 = n1677 ^ n1533;
  assign n1781 = n1680 ^ n1678;
  assign n1782 = ~n1681 & ~n1781;
  assign n1783 = n1782 ^ n1678;
  assign n1682 = n1681 ^ n1678;
  assign n1439 = x147 & x148;
  assign n1440 = x149 & x150;
  assign n1441 = ~n1439 & ~n1440;
  assign n1442 = ~x147 & ~x148;
  assign n1443 = ~x149 & ~x150;
  assign n1444 = ~n1442 & ~n1443;
  assign n1445 = ~n1441 & n1444;
  assign n1446 = x146 & n1445;
  assign n1447 = n1439 & n1440;
  assign n1448 = ~n1446 & ~n1447;
  assign n1449 = n1441 & ~n1444;
  assign n1450 = ~x146 & n1449;
  assign n1451 = n1442 & n1443;
  assign n1452 = ~n1450 & ~n1451;
  assign n1453 = n1448 & n1452;
  assign n1454 = ~x145 & ~n1453;
  assign n1365 = x146 ^ x145;
  assign n1455 = n1365 & n1445;
  assign n1456 = x145 & x146;
  assign n1457 = n1439 & n1456;
  assign n1458 = x150 & n1457;
  assign n1459 = n1458 ^ n1456;
  assign n1460 = ~n1449 & n1459;
  assign n1461 = ~n1455 & ~n1460;
  assign n1462 = ~x146 & ~x150;
  assign n1463 = n1442 & n1462;
  assign n1464 = ~n1457 & ~n1463;
  assign n1465 = ~x149 & ~n1464;
  assign n1466 = n1461 & ~n1465;
  assign n1467 = ~n1454 & n1466;
  assign n1410 = x141 & x142;
  assign n1411 = x143 & x144;
  assign n1412 = ~n1410 & ~n1411;
  assign n1413 = ~x141 & ~x142;
  assign n1414 = ~x143 & ~x144;
  assign n1415 = ~n1413 & ~n1414;
  assign n1416 = ~n1412 & n1415;
  assign n1417 = x140 & n1416;
  assign n1418 = n1410 & n1411;
  assign n1419 = ~n1417 & ~n1418;
  assign n1420 = n1412 & ~n1415;
  assign n1421 = ~x140 & n1420;
  assign n1422 = n1413 & n1414;
  assign n1423 = ~n1421 & ~n1422;
  assign n1424 = n1419 & n1423;
  assign n1425 = ~x139 & ~n1424;
  assign n1360 = x140 ^ x139;
  assign n1426 = n1360 & n1416;
  assign n1427 = x139 & x140;
  assign n1428 = n1410 & n1427;
  assign n1429 = x144 & n1428;
  assign n1430 = n1429 ^ n1427;
  assign n1431 = ~n1420 & n1430;
  assign n1432 = ~n1426 & ~n1431;
  assign n1433 = ~x140 & ~x144;
  assign n1434 = n1413 & n1433;
  assign n1435 = ~n1428 & ~n1434;
  assign n1436 = ~x143 & ~n1435;
  assign n1437 = n1432 & ~n1436;
  assign n1438 = ~n1425 & n1437;
  assign n1468 = n1467 ^ n1438;
  assign n1359 = x142 ^ x141;
  assign n1361 = n1360 ^ n1359;
  assign n1358 = x144 ^ x143;
  assign n1362 = n1361 ^ n1358;
  assign n1364 = x148 ^ x147;
  assign n1366 = n1365 ^ n1364;
  assign n1363 = x150 ^ x149;
  assign n1367 = n1366 ^ n1363;
  assign n1684 = n1362 & n1367;
  assign n1685 = n1684 ^ n1438;
  assign n1686 = n1468 & ~n1685;
  assign n1687 = n1686 ^ n1467;
  assign n1405 = n1362 ^ n1356;
  assign n1407 = n1405 ^ n1351;
  assign n1408 = ~n1367 & n1407;
  assign n1357 = n1356 ^ n1351;
  assign n1406 = ~n1357 & ~n1405;
  assign n1409 = n1408 ^ n1406;
  assign n1469 = n1468 ^ n1409;
  assign n1688 = ~n1469 & ~n1534;
  assign n1368 = n1367 ^ n1362;
  assign n1369 = n1368 ^ n1357;
  assign n1689 = ~n1356 & ~n1684;
  assign n1690 = n1369 & n1689;
  assign n1691 = ~n1362 & ~n1367;
  assign n1692 = ~n1690 & ~n1691;
  assign n1693 = ~n1468 & ~n1692;
  assign n1694 = n1468 & n1684;
  assign n1695 = ~n1693 & ~n1694;
  assign n1696 = ~n1688 & n1695;
  assign n1697 = n1534 & n1675;
  assign n1698 = n1696 & ~n1697;
  assign n1784 = ~n1687 & ~n1698;
  assign n1789 = n1682 & ~n1784;
  assign n1812 = ~n1783 & ~n1789;
  assign n1672 = n1448 & n1461;
  assign n1673 = n1419 & n1432;
  assign n1790 = ~n1672 & ~n1673;
  assign n1785 = ~n1682 & n1784;
  assign n1674 = n1673 ^ n1672;
  assign n1786 = n1687 & n1698;
  assign n1787 = n1674 & ~n1786;
  assign n1788 = ~n1785 & n1787;
  assign n1792 = n1672 & n1673;
  assign n1791 = ~n1786 & ~n1790;
  assign n1793 = n1792 ^ n1791;
  assign n1794 = ~n1789 & ~n1793;
  assign n1795 = n1794 ^ n1792;
  assign n1796 = ~n1788 & ~n1795;
  assign n1797 = n1796 ^ n1783;
  assign n1818 = ~n1790 & ~n1797;
  assign n1819 = ~n1812 & ~n1818;
  assign n1721 = n1720 ^ n1717;
  assign n1539 = x161 & x162;
  assign n1540 = x159 & x160;
  assign n1541 = n1539 & n1540;
  assign n1542 = ~x161 & ~x162;
  assign n1543 = x158 & ~n1542;
  assign n1544 = ~n1541 & ~n1543;
  assign n1372 = x160 ^ x159;
  assign n1545 = n1539 ^ x160;
  assign n1546 = n1372 & ~n1545;
  assign n1547 = n1546 ^ x159;
  assign n1548 = ~n1544 & n1547;
  assign n1549 = ~x159 & ~x160;
  assign n1550 = ~n1539 & n1549;
  assign n1551 = ~n1543 & n1550;
  assign n1552 = ~x158 & ~n1540;
  assign n1553 = n1542 & n1552;
  assign n1554 = ~n1551 & ~n1553;
  assign n1555 = ~n1548 & n1554;
  assign n1556 = ~x157 & ~n1555;
  assign n1557 = x157 & ~n1542;
  assign n1558 = n1547 & n1557;
  assign n1559 = x157 & x158;
  assign n1560 = ~n1558 & ~n1559;
  assign n1561 = ~n1540 & ~n1542;
  assign n1562 = ~n1550 & n1561;
  assign n1563 = ~x162 & n1540;
  assign n1564 = x158 & ~n1563;
  assign n1565 = ~n1562 & n1564;
  assign n1566 = ~n1560 & ~n1565;
  assign n1567 = ~n1556 & ~n1566;
  assign n1568 = n1540 & n1559;
  assign n1569 = ~x158 & ~x162;
  assign n1570 = n1549 & n1569;
  assign n1571 = ~n1568 & ~n1570;
  assign n1572 = ~x161 & ~n1571;
  assign n1573 = n1567 & ~n1572;
  assign n1574 = ~x155 & ~x156;
  assign n1575 = x152 & ~n1574;
  assign n1576 = x155 & x156;
  assign n1577 = x153 & x154;
  assign n1578 = n1576 & n1577;
  assign n1579 = ~n1575 & ~n1578;
  assign n1376 = x154 ^ x153;
  assign n1580 = n1576 ^ x154;
  assign n1581 = n1376 & ~n1580;
  assign n1582 = n1581 ^ x153;
  assign n1583 = ~n1579 & n1582;
  assign n1584 = ~x153 & ~x154;
  assign n1585 = ~n1576 & n1584;
  assign n1586 = ~n1575 & n1585;
  assign n1587 = ~n1583 & ~n1586;
  assign n1588 = ~x151 & ~n1587;
  assign n1589 = x151 & ~n1574;
  assign n1590 = n1582 & n1589;
  assign n1591 = x151 & x152;
  assign n1592 = ~n1590 & ~n1591;
  assign n1593 = ~n1574 & ~n1577;
  assign n1594 = ~n1585 & n1593;
  assign n1595 = ~x156 & n1577;
  assign n1596 = x152 & ~n1595;
  assign n1597 = ~n1594 & n1596;
  assign n1598 = ~n1592 & ~n1597;
  assign n1599 = ~n1588 & ~n1598;
  assign n1600 = x151 & ~n1584;
  assign n1601 = ~x152 & ~x156;
  assign n1602 = ~n1577 & n1601;
  assign n1603 = ~n1600 & n1602;
  assign n1604 = n1577 & n1591;
  assign n1605 = ~n1603 & ~n1604;
  assign n1606 = ~x155 & ~n1605;
  assign n1607 = n1599 & ~n1606;
  assign n1713 = n1573 & n1607;
  assign n1711 = ~n1583 & ~n1598;
  assign n1710 = ~n1548 & ~n1566;
  assign n1712 = n1711 ^ n1710;
  assign n1714 = n1713 ^ n1712;
  assign n1722 = n1721 ^ n1714;
  assign n1661 = n1660 ^ n1609;
  assign n1608 = n1607 ^ n1573;
  assign n1662 = n1661 ^ n1608;
  assign n1377 = x156 ^ x155;
  assign n1378 = n1377 ^ n1376;
  assign n1375 = x152 ^ x151;
  assign n1379 = n1378 ^ n1375;
  assign n1371 = x162 ^ x161;
  assign n1373 = n1372 ^ n1371;
  assign n1370 = x158 ^ x157;
  assign n1374 = n1373 ^ n1370;
  assign n1380 = n1379 ^ n1374;
  assign n1391 = n1390 ^ n1385;
  assign n1536 = n1391 ^ n1379;
  assign n1537 = ~n1380 & n1536;
  assign n1538 = n1537 ^ n1391;
  assign n1707 = n1608 ^ n1538;
  assign n1708 = n1662 & ~n1707;
  assign n1709 = n1708 ^ n1661;
  assign n1723 = n1722 ^ n1709;
  assign n1392 = n1391 ^ n1380;
  assign n1393 = n1369 & n1392;
  assign n1535 = n1534 ^ n1469;
  assign n1701 = n1374 & n1379;
  assign n1702 = n1701 ^ n1662;
  assign n1703 = n1535 & ~n1702;
  assign n1704 = n1393 & ~n1703;
  assign n1663 = n1662 ^ n1538;
  assign n1705 = ~n1535 & n1663;
  assign n1706 = ~n1704 & ~n1705;
  assign n1724 = n1723 ^ n1706;
  assign n1699 = n1698 ^ n1687;
  assign n1683 = n1682 ^ n1674;
  assign n1700 = n1699 ^ n1683;
  assign n1766 = n1706 ^ n1700;
  assign n1767 = ~n1724 & n1766;
  assign n1768 = n1767 ^ n1723;
  assign n1769 = n1721 ^ n1709;
  assign n1770 = ~n1722 & n1769;
  assign n1771 = n1770 ^ n1709;
  assign n1775 = n1713 ^ n1711;
  assign n1776 = ~n1712 & ~n1775;
  assign n1777 = n1776 ^ n1713;
  assign n1813 = ~n1771 & ~n1777;
  assign n1814 = ~n1768 & n1813;
  assign n1836 = ~n1797 & ~n1814;
  assign n1837 = ~n1819 & ~n1836;
  assign n1838 = ~n1774 & ~n1837;
  assign n1839 = ~n1813 & n1819;
  assign n1824 = n1771 & n1777;
  assign n1840 = n1768 & n1824;
  assign n1841 = ~n1839 & ~n1840;
  assign n1842 = n1838 & n1841;
  assign n1820 = n1771 ^ n1768;
  assign n1821 = n1777 ^ n1771;
  assign n1822 = n1820 & ~n1821;
  assign n1823 = n1822 ^ n1768;
  assign n1829 = ~n1819 & ~n1823;
  assign n1778 = n1777 ^ n1774;
  assign n1779 = n1778 ^ n1771;
  assign n1830 = n1779 & ~n1824;
  assign n1831 = ~n1768 & n1830;
  assign n1832 = ~n1812 & ~n1831;
  assign n1833 = n1797 & ~n1832;
  assign n1850 = ~n1829 & ~n1833;
  assign n1851 = ~n1842 & n1850;
  assign n1191 = x107 & x108;
  assign n1192 = x105 & x106;
  assign n1193 = n1191 & n1192;
  assign n1194 = ~x107 & ~x108;
  assign n1195 = x104 & ~n1194;
  assign n1196 = ~n1193 & ~n1195;
  assign n1157 = x106 ^ x105;
  assign n1197 = n1191 ^ x106;
  assign n1198 = n1157 & ~n1197;
  assign n1199 = n1198 ^ x105;
  assign n1200 = ~n1196 & n1199;
  assign n1209 = x103 & ~n1194;
  assign n1210 = n1199 & n1209;
  assign n1211 = x103 & x104;
  assign n1212 = ~n1210 & ~n1211;
  assign n1201 = ~x105 & ~x106;
  assign n1202 = ~n1191 & n1201;
  assign n1213 = ~n1192 & ~n1194;
  assign n1214 = ~n1202 & n1213;
  assign n1215 = ~x108 & n1192;
  assign n1216 = x104 & ~n1215;
  assign n1217 = ~n1214 & n1216;
  assign n1218 = ~n1212 & ~n1217;
  assign n1339 = ~n1200 & ~n1218;
  assign n1203 = ~n1195 & n1202;
  assign n1204 = ~x104 & ~n1192;
  assign n1205 = n1194 & n1204;
  assign n1206 = ~n1203 & ~n1205;
  assign n1207 = ~n1200 & n1206;
  assign n1208 = ~x103 & ~n1207;
  assign n1219 = ~n1208 & ~n1218;
  assign n1220 = n1192 & n1211;
  assign n1221 = ~x104 & ~x108;
  assign n1222 = n1201 & n1221;
  assign n1223 = ~n1220 & ~n1222;
  assign n1224 = ~x107 & ~n1223;
  assign n1225 = n1219 & ~n1224;
  assign n1163 = ~x111 & ~x112;
  assign n1164 = ~x113 & ~x114;
  assign n1165 = ~n1163 & ~n1164;
  assign n1166 = x111 & x112;
  assign n1167 = x113 & x114;
  assign n1168 = ~n1166 & ~n1167;
  assign n1169 = n1165 & ~n1168;
  assign n1170 = x110 & n1169;
  assign n1171 = n1166 & n1167;
  assign n1172 = ~n1170 & ~n1171;
  assign n1173 = ~n1165 & n1168;
  assign n1150 = x112 ^ x111;
  assign n1149 = x114 ^ x113;
  assign n1151 = n1150 ^ n1149;
  assign n1174 = x110 & n1151;
  assign n1175 = n1173 & ~n1174;
  assign n1176 = n1172 & ~n1175;
  assign n1177 = ~x109 & ~n1176;
  assign n1148 = x110 ^ x109;
  assign n1178 = n1148 & n1169;
  assign n1179 = x109 & x110;
  assign n1180 = n1166 & n1179;
  assign n1181 = x114 & n1180;
  assign n1182 = n1181 ^ n1179;
  assign n1183 = ~n1173 & n1182;
  assign n1184 = ~n1178 & ~n1183;
  assign n1185 = ~x110 & ~x114;
  assign n1186 = n1163 & n1185;
  assign n1187 = ~n1180 & ~n1186;
  assign n1188 = ~x113 & ~n1187;
  assign n1189 = n1184 & ~n1188;
  assign n1190 = ~n1177 & n1189;
  assign n1226 = n1225 ^ n1190;
  assign n1152 = n1151 ^ n1148;
  assign n1156 = x108 ^ x107;
  assign n1158 = n1157 ^ n1156;
  assign n1155 = x104 ^ x103;
  assign n1159 = n1158 ^ n1155;
  assign n1314 = n1152 & n1159;
  assign n1336 = n1314 ^ n1190;
  assign n1337 = n1226 & ~n1336;
  assign n1338 = n1337 ^ n1225;
  assign n1340 = n1339 ^ n1338;
  assign n1335 = n1172 & n1184;
  assign n1341 = n1340 ^ n1335;
  assign n1254 = x117 & x118;
  assign n1255 = x119 & x120;
  assign n1256 = ~n1254 & ~n1255;
  assign n1257 = ~x117 & ~x118;
  assign n1258 = ~x119 & ~x120;
  assign n1259 = ~n1257 & ~n1258;
  assign n1260 = ~n1256 & n1259;
  assign n1261 = x116 & n1260;
  assign n1262 = n1254 & n1255;
  assign n1263 = ~n1261 & ~n1262;
  assign n1264 = n1256 & ~n1259;
  assign n1268 = ~n1262 & ~n1264;
  assign n1269 = x116 & ~n1268;
  assign n1270 = ~x116 & ~n1260;
  assign n1271 = x115 & ~n1270;
  assign n1272 = ~n1269 & n1271;
  assign n1332 = n1263 & ~n1272;
  assign n1231 = ~x125 & ~x126;
  assign n1229 = x125 & x126;
  assign n1234 = x123 & x124;
  assign n1246 = ~n1229 & ~n1234;
  assign n1144 = x122 ^ x121;
  assign n1228 = ~x123 & ~x124;
  assign n1247 = n1144 & ~n1228;
  assign n1248 = ~n1246 & n1247;
  assign n1230 = n1228 & ~n1229;
  assign n1241 = x121 & x122;
  assign n1249 = ~n1234 & n1241;
  assign n1250 = ~n1230 & n1249;
  assign n1251 = ~n1248 & ~n1250;
  assign n1252 = ~n1231 & ~n1251;
  assign n1235 = n1229 & n1234;
  assign n1242 = n1234 & n1241;
  assign n1330 = ~n1235 & ~n1242;
  assign n1331 = ~n1252 & n1330;
  assign n1333 = n1332 ^ n1331;
  assign n1265 = ~x116 & n1264;
  assign n1266 = n1263 & ~n1265;
  assign n1267 = ~x115 & ~n1266;
  assign n1139 = x116 ^ x115;
  assign n1273 = n1257 & n1258;
  assign n1274 = n1139 & n1273;
  assign n1275 = ~n1272 & ~n1274;
  assign n1276 = ~n1267 & n1275;
  assign n1232 = x122 & ~n1231;
  assign n1233 = n1230 & ~n1232;
  assign n1236 = ~n1233 & ~n1235;
  assign n1237 = ~x121 & ~n1236;
  assign n1143 = x126 ^ x125;
  assign n1145 = n1144 ^ n1143;
  assign n1142 = x124 ^ x123;
  assign n1146 = n1145 ^ n1142;
  assign n1238 = ~x122 & n1231;
  assign n1239 = ~n1234 & n1238;
  assign n1240 = n1146 & n1239;
  assign n1243 = ~n1229 & n1242;
  assign n1244 = ~n1240 & ~n1243;
  assign n1245 = ~n1237 & n1244;
  assign n1253 = n1245 & ~n1252;
  assign n1277 = n1276 ^ n1253;
  assign n1138 = x118 ^ x117;
  assign n1140 = n1139 ^ n1138;
  assign n1137 = x120 ^ x119;
  assign n1141 = n1140 ^ n1137;
  assign n1317 = n1141 & n1146;
  assign n1327 = n1317 ^ n1253;
  assign n1328 = n1277 & ~n1327;
  assign n1329 = n1328 ^ n1276;
  assign n1334 = n1333 ^ n1329;
  assign n1342 = n1341 ^ n1334;
  assign n1315 = n1226 & n1314;
  assign n1153 = n1152 ^ n1146;
  assign n1160 = n1153 ^ n1141;
  assign n1161 = ~n1159 & n1160;
  assign n1147 = n1146 ^ n1141;
  assign n1154 = ~n1147 & ~n1153;
  assign n1162 = n1161 ^ n1154;
  assign n1227 = n1226 ^ n1162;
  assign n1316 = ~n1227 & ~n1277;
  assign n1318 = n1277 & n1317;
  assign n1280 = n1159 ^ n1152;
  assign n1281 = n1280 ^ n1147;
  assign n1319 = ~n1141 & ~n1314;
  assign n1320 = n1281 & n1319;
  assign n1321 = ~n1152 & ~n1159;
  assign n1322 = ~n1320 & ~n1321;
  assign n1323 = ~n1226 & ~n1322;
  assign n1324 = ~n1318 & ~n1323;
  assign n1325 = ~n1316 & n1324;
  assign n1326 = ~n1315 & n1325;
  assign n1343 = n1342 ^ n1326;
  assign n1732 = n1339 ^ n1326;
  assign n1733 = ~n1340 & n1732;
  assign n1734 = n1733 ^ n1338;
  assign n1735 = n1335 & ~n1734;
  assign n1736 = n1343 & n1735;
  assign n1737 = ~n1338 & n1339;
  assign n1738 = ~n1334 & n1737;
  assign n1739 = ~n1326 & n1738;
  assign n1740 = ~n1736 & ~n1739;
  assign n1729 = n1332 ^ n1329;
  assign n1730 = ~n1333 & ~n1729;
  assign n1731 = n1730 ^ n1329;
  assign n1741 = n1334 & n1734;
  assign n1742 = ~n1343 & n1741;
  assign n1807 = ~n1731 & ~n1742;
  assign n1808 = n1740 & ~n1807;
  assign n1015 = x92 ^ x91;
  assign n1014 = x94 ^ x93;
  assign n1016 = n1015 ^ n1014;
  assign n1013 = x96 ^ x95;
  assign n1017 = n1016 ^ n1013;
  assign n1020 = x98 ^ x97;
  assign n1019 = x100 ^ x99;
  assign n1021 = n1020 ^ n1019;
  assign n1018 = x102 ^ x101;
  assign n1022 = n1021 ^ n1018;
  assign n1025 = n1017 & n1022;
  assign n1057 = x95 & x96;
  assign n1058 = ~x93 & ~x94;
  assign n1059 = ~n1057 & n1058;
  assign n1060 = ~x95 & ~x96;
  assign n1061 = x92 & ~n1060;
  assign n1062 = n1059 & ~n1061;
  assign n1063 = x93 & x94;
  assign n1064 = n1057 & n1063;
  assign n1065 = ~n1062 & ~n1064;
  assign n1066 = ~x91 & ~n1065;
  assign n1067 = ~x92 & n1060;
  assign n1068 = ~n1063 & n1067;
  assign n1069 = n1016 & n1068;
  assign n1070 = x91 & x92;
  assign n1071 = n1063 & n1070;
  assign n1072 = ~n1057 & n1071;
  assign n1073 = ~n1069 & ~n1072;
  assign n1074 = ~n1066 & n1073;
  assign n1075 = ~n1057 & ~n1063;
  assign n1076 = n1015 & ~n1058;
  assign n1077 = ~n1075 & n1076;
  assign n1078 = ~n1063 & n1070;
  assign n1079 = ~n1059 & n1078;
  assign n1080 = ~n1077 & ~n1079;
  assign n1081 = ~n1060 & ~n1080;
  assign n1082 = n1074 & ~n1081;
  assign n1031 = x101 & x102;
  assign n1032 = ~x99 & ~x100;
  assign n1033 = ~n1031 & n1032;
  assign n1034 = ~x101 & ~x102;
  assign n1035 = x98 & ~n1034;
  assign n1036 = n1033 & ~n1035;
  assign n1037 = x99 & x100;
  assign n1038 = n1031 & n1037;
  assign n1039 = ~n1036 & ~n1038;
  assign n1040 = ~x97 & ~n1039;
  assign n1041 = ~x98 & n1034;
  assign n1042 = ~n1037 & n1041;
  assign n1043 = n1021 & n1042;
  assign n1044 = x97 & x98;
  assign n1045 = n1037 & n1044;
  assign n1046 = ~n1031 & n1045;
  assign n1047 = ~n1043 & ~n1046;
  assign n1048 = ~n1040 & n1047;
  assign n1049 = ~n1031 & ~n1037;
  assign n1050 = n1020 & ~n1032;
  assign n1051 = ~n1049 & n1050;
  assign n1052 = ~n1037 & n1044;
  assign n1053 = ~n1033 & n1052;
  assign n1054 = ~n1051 & ~n1053;
  assign n1055 = ~n1034 & ~n1054;
  assign n1056 = n1048 & ~n1055;
  assign n1083 = n1082 ^ n1056;
  assign n1294 = n1025 & n1083;
  assign n1295 = n1056 & n1082;
  assign n1296 = ~n1294 & ~n1295;
  assign n1291 = ~n1064 & ~n1071;
  assign n1292 = ~n1081 & n1291;
  assign n1289 = ~n1038 & ~n1045;
  assign n1290 = ~n1055 & n1289;
  assign n1293 = n1292 ^ n1290;
  assign n1297 = n1296 ^ n1293;
  assign n1106 = x83 & x84;
  assign n1107 = x81 & x82;
  assign n1108 = n1106 & n1107;
  assign n1109 = ~x83 & ~x84;
  assign n1110 = x80 & ~n1109;
  assign n1111 = ~n1108 & ~n1110;
  assign n1003 = x82 ^ x81;
  assign n1112 = n1106 ^ x82;
  assign n1113 = n1003 & ~n1112;
  assign n1114 = n1113 ^ x81;
  assign n1115 = ~n1111 & n1114;
  assign n1118 = ~x81 & ~x82;
  assign n1119 = ~n1106 & n1118;
  assign n1126 = ~n1108 & ~n1119;
  assign n1116 = ~n1107 & n1109;
  assign n1127 = x79 & ~n1116;
  assign n1128 = n1126 & n1127;
  assign n1129 = x79 & ~x80;
  assign n1130 = ~n1128 & ~n1129;
  assign n1131 = ~n1109 & n1114;
  assign n1132 = ~x80 & ~n1131;
  assign n1133 = ~n1130 & ~n1132;
  assign n1309 = ~n1115 & ~n1133;
  assign n1088 = x87 & x88;
  assign n1089 = x89 & x90;
  assign n1093 = n1088 & n1089;
  assign n1085 = ~x87 & ~x88;
  assign n1086 = ~x89 & ~x90;
  assign n1087 = ~n1085 & ~n1086;
  assign n1090 = ~n1088 & ~n1089;
  assign n1091 = ~n1087 & n1090;
  assign n1096 = x85 & x86;
  assign n1097 = ~n1093 & n1096;
  assign n1098 = ~n1091 & n1097;
  assign n1009 = x86 ^ x85;
  assign n1099 = n1087 & ~n1090;
  assign n1100 = n1009 & n1099;
  assign n1101 = ~n1098 & ~n1100;
  assign n1308 = ~n1093 & n1101;
  assign n1310 = n1309 ^ n1308;
  assign n1117 = ~x80 & n1116;
  assign n1120 = ~n1110 & n1119;
  assign n1121 = ~n1117 & ~n1120;
  assign n1122 = ~n1115 & n1121;
  assign n1123 = ~x79 & ~n1122;
  assign n1124 = n1117 & n1118;
  assign n1125 = ~n1123 & ~n1124;
  assign n1134 = n1125 & ~n1133;
  assign n1092 = ~x86 & n1091;
  assign n1094 = ~n1092 & ~n1093;
  assign n1095 = ~x85 & ~n1094;
  assign n1102 = n1085 & ~n1096;
  assign n1103 = n1086 & n1102;
  assign n1104 = n1101 & ~n1103;
  assign n1105 = ~n1095 & n1104;
  assign n1135 = n1134 ^ n1105;
  assign n1004 = x84 ^ x83;
  assign n1005 = n1004 ^ n1003;
  assign n1002 = x80 ^ x79;
  assign n1006 = n1005 ^ n1002;
  assign n1008 = x88 ^ x87;
  assign n1010 = n1009 ^ n1008;
  assign n1007 = x90 ^ x89;
  assign n1011 = n1010 ^ n1007;
  assign n1012 = n1006 & n1011;
  assign n1305 = n1105 ^ n1012;
  assign n1306 = n1135 & ~n1305;
  assign n1307 = n1306 ^ n1134;
  assign n1311 = n1310 ^ n1307;
  assign n1298 = n1012 & n1135;
  assign n1023 = ~n1017 & ~n1022;
  assign n1024 = ~n1012 & n1023;
  assign n1026 = ~n1006 & ~n1011;
  assign n1027 = ~n1025 & n1026;
  assign n1028 = ~n1024 & ~n1027;
  assign n1029 = n1012 & n1025;
  assign n1030 = n1028 & ~n1029;
  assign n1084 = n1083 ^ n1030;
  assign n1299 = n1084 & ~n1135;
  assign n1300 = n1028 ^ n1025;
  assign n1301 = ~n1083 & ~n1300;
  assign n1302 = n1301 ^ n1025;
  assign n1303 = ~n1299 & ~n1302;
  assign n1304 = ~n1298 & n1303;
  assign n1312 = n1311 ^ n1304;
  assign n1756 = n1297 & n1312;
  assign n1751 = ~n1307 & n1309;
  assign n1757 = n1756 ^ n1751;
  assign n1752 = ~n1304 & n1308;
  assign n1758 = n1752 ^ n1751;
  assign n1759 = n1757 & ~n1758;
  assign n1760 = n1759 ^ n1756;
  assign n1748 = n1296 ^ n1292;
  assign n1749 = ~n1293 & n1748;
  assign n1750 = n1749 ^ n1296;
  assign n1753 = ~n1751 & ~n1752;
  assign n1754 = ~n1297 & n1312;
  assign n1755 = n1753 & n1754;
  assign n1805 = n1750 & ~n1755;
  assign n1806 = ~n1760 & ~n1805;
  assign n1809 = n1808 ^ n1806;
  assign n1761 = ~n1755 & ~n1760;
  assign n1762 = n1761 ^ n1750;
  assign n1313 = n1312 ^ n1297;
  assign n1344 = n1343 ^ n1313;
  assign n1278 = n1277 ^ n1227;
  assign n1136 = n1135 ^ n1084;
  assign n1279 = n1278 ^ n1136;
  assign n1283 = n1011 ^ n1006;
  assign n1282 = n1022 ^ n1017;
  assign n1284 = n1283 ^ n1282;
  assign n1285 = n1281 & n1284;
  assign n1286 = n1285 ^ n1136;
  assign n1287 = ~n1279 & ~n1286;
  assign n1288 = n1287 ^ n1278;
  assign n1745 = n1313 ^ n1288;
  assign n1746 = ~n1344 & ~n1745;
  assign n1747 = n1746 ^ n1343;
  assign n1763 = n1762 ^ n1747;
  assign n1743 = n1740 & ~n1742;
  assign n1744 = n1743 ^ n1731;
  assign n1802 = n1747 ^ n1744;
  assign n1803 = ~n1763 & ~n1802;
  assign n1804 = n1803 ^ n1762;
  assign n1847 = n1808 ^ n1804;
  assign n1848 = ~n1809 & ~n1847;
  assign n1849 = n1848 ^ n1804;
  assign n1852 = n1851 ^ n1849;
  assign n1810 = n1809 ^ n1804;
  assign n1764 = n1763 ^ n1744;
  assign n1346 = ~n1279 & n1285;
  assign n1394 = n1285 & n1393;
  assign n1395 = n1284 ^ n1281;
  assign n1396 = n1392 ^ n1369;
  assign n1397 = n1396 ^ n1284;
  assign n1398 = n1395 & ~n1397;
  assign n1399 = n1398 ^ n1281;
  assign n1400 = n1399 ^ n1285;
  assign n1401 = ~n1393 & ~n1400;
  assign n1402 = n1401 ^ n1285;
  assign n1403 = ~n1279 & ~n1402;
  assign n1404 = ~n1394 & ~n1403;
  assign n1664 = n1663 ^ n1535;
  assign n1665 = n1404 & n1664;
  assign n1666 = ~n1346 & ~n1665;
  assign n1667 = n1279 & ~n1399;
  assign n1668 = ~n1393 & ~n1667;
  assign n1669 = ~n1664 & ~n1668;
  assign n1670 = n1666 & ~n1669;
  assign n1345 = n1344 ^ n1288;
  assign n1671 = n1670 ^ n1345;
  assign n1725 = n1724 ^ n1700;
  assign n1726 = n1725 ^ n1345;
  assign n1727 = n1671 & n1726;
  assign n1728 = n1727 ^ n1670;
  assign n1765 = n1764 ^ n1728;
  assign n1780 = n1779 ^ n1768;
  assign n1798 = n1797 ^ n1780;
  assign n1799 = n1798 ^ n1728;
  assign n1800 = ~n1765 & n1799;
  assign n1801 = n1800 ^ n1764;
  assign n1811 = n1810 ^ n1801;
  assign n1815 = n1812 & ~n1814;
  assign n1816 = n1797 & ~n1815;
  assign n1817 = n1774 & ~n1816;
  assign n1825 = n1824 ^ n1823;
  assign n1826 = ~n1819 & ~n1825;
  assign n1827 = n1826 ^ n1824;
  assign n1828 = n1817 & n1827;
  assign n1834 = ~n1829 & n1833;
  assign n1835 = ~n1828 & ~n1834;
  assign n1843 = n1835 & ~n1842;
  assign n1844 = n1843 ^ n1801;
  assign n1845 = ~n1811 & n1844;
  assign n1846 = n1845 ^ n1843;
  assign n1853 = n1852 ^ n1846;
  assign n2647 = n2646 ^ n1853;
  assign n2648 = n1843 ^ n1811;
  assign n2649 = n2648 ^ n2620;
  assign n2667 = n2595 ^ n2571;
  assign n2661 = n1725 ^ n1671;
  assign n2650 = n1396 ^ n1395;
  assign n2651 = ~n2578 & ~n2579;
  assign n2652 = n2650 & ~n2651;
  assign n2653 = ~n2577 & n2652;
  assign n2654 = n1402 ^ n1279;
  assign n2655 = n2654 ^ n1664;
  assign n2656 = ~n2653 & n2655;
  assign n2657 = ~n2580 & ~n2652;
  assign n2658 = n2657 ^ n2577;
  assign n2659 = ~n2581 & ~n2658;
  assign n2660 = ~n2656 & ~n2659;
  assign n2662 = n2661 ^ n2660;
  assign n2663 = n2592 ^ n2575;
  assign n2664 = n2663 ^ n2661;
  assign n2665 = n2662 & ~n2664;
  assign n2666 = n2665 ^ n2663;
  assign n2668 = n2667 ^ n2666;
  assign n2669 = n1798 ^ n1765;
  assign n2670 = n2669 ^ n2666;
  assign n2671 = ~n2668 & ~n2670;
  assign n2672 = n2671 ^ n2667;
  assign n2673 = n2672 ^ n2648;
  assign n2674 = ~n2649 & ~n2673;
  assign n2675 = n2674 ^ n2620;
  assign n2676 = n2675 ^ n1853;
  assign n2677 = n2647 & ~n2676;
  assign n2678 = n2677 ^ n2646;
  assign n2679 = n1851 ^ n1846;
  assign n2680 = n1852 & ~n2679;
  assign n2681 = n2680 ^ n1846;
  assign n2682 = ~n2678 & n2681;
  assign n3547 = x314 ^ x313;
  assign n3548 = x316 ^ x315;
  assign n3549 = x317 & x318;
  assign n3550 = n3549 ^ x316;
  assign n3551 = n3548 & ~n3550;
  assign n3552 = n3551 ^ x315;
  assign n3553 = n3547 & n3552;
  assign n3554 = ~x315 & ~x316;
  assign n3555 = ~n3549 & n3554;
  assign n3556 = x315 & x316;
  assign n3557 = x313 & x314;
  assign n3558 = ~n3556 & n3557;
  assign n3559 = ~n3555 & n3558;
  assign n3560 = ~n3553 & ~n3559;
  assign n3561 = ~x317 & ~x318;
  assign n3562 = ~n3560 & ~n3561;
  assign n3563 = n3556 & n3557;
  assign n3564 = ~x318 & n3563;
  assign n3565 = ~n3562 & ~n3564;
  assign n3566 = x314 & ~n3561;
  assign n3567 = n3549 & n3556;
  assign n3568 = ~n3566 & ~n3567;
  assign n3569 = n3552 & ~n3568;
  assign n3570 = n3555 & ~n3566;
  assign n3571 = ~n3569 & ~n3570;
  assign n3572 = ~x313 & ~n3571;
  assign n3573 = n3565 & ~n3572;
  assign n3574 = n3548 ^ n3547;
  assign n3575 = ~x314 & ~x318;
  assign n3576 = ~n3556 & n3575;
  assign n3577 = n3574 & n3576;
  assign n3578 = ~n3563 & ~n3577;
  assign n3579 = ~x317 & ~n3578;
  assign n3580 = n3573 & ~n3579;
  assign n3512 = ~x311 & ~x312;
  assign n3513 = x308 & ~n3512;
  assign n3514 = x311 & x312;
  assign n3515 = x309 & x310;
  assign n3516 = n3514 & n3515;
  assign n3517 = ~n3513 & ~n3516;
  assign n3518 = x310 ^ x309;
  assign n3519 = n3514 ^ x310;
  assign n3520 = n3518 & ~n3519;
  assign n3521 = n3520 ^ x309;
  assign n3522 = ~n3517 & n3521;
  assign n3523 = ~x309 & ~x310;
  assign n3524 = ~n3514 & n3523;
  assign n3525 = ~n3513 & n3524;
  assign n3526 = ~n3522 & ~n3525;
  assign n3527 = ~x307 & ~n3526;
  assign n3528 = x307 & ~n3512;
  assign n3529 = n3521 & n3528;
  assign n3530 = x307 & x308;
  assign n3531 = ~n3529 & ~n3530;
  assign n3532 = ~n3512 & ~n3515;
  assign n3533 = ~n3524 & n3532;
  assign n3534 = ~x312 & n3515;
  assign n3535 = x308 & ~n3534;
  assign n3536 = ~n3533 & n3535;
  assign n3537 = ~n3531 & ~n3536;
  assign n3538 = ~n3527 & ~n3537;
  assign n3539 = x307 & ~n3523;
  assign n3540 = ~x308 & ~x312;
  assign n3541 = ~n3515 & n3540;
  assign n3542 = ~n3539 & n3541;
  assign n3543 = n3515 & n3530;
  assign n3544 = ~n3542 & ~n3543;
  assign n3545 = ~x311 & ~n3544;
  assign n3546 = n3538 & ~n3545;
  assign n3581 = n3580 ^ n3546;
  assign n3583 = x312 ^ x311;
  assign n3584 = n3583 ^ n3518;
  assign n3582 = x308 ^ x307;
  assign n3585 = n3584 ^ n3582;
  assign n3586 = x318 ^ x317;
  assign n3587 = n3586 ^ n3574;
  assign n3588 = n3585 & n3587;
  assign n3589 = n3581 & n3588;
  assign n3620 = ~x305 & ~x306;
  assign n3621 = ~x303 & ~x304;
  assign n3622 = ~n3620 & ~n3621;
  assign n3623 = x305 & x306;
  assign n3624 = x303 & x304;
  assign n3625 = ~n3623 & ~n3624;
  assign n3626 = n3622 & ~n3625;
  assign n3627 = x302 & n3626;
  assign n3628 = n3623 & n3624;
  assign n3629 = ~n3627 & ~n3628;
  assign n3630 = ~n3622 & n3625;
  assign n3631 = ~x302 & n3630;
  assign n3632 = n3620 & n3621;
  assign n3633 = ~n3631 & ~n3632;
  assign n3634 = n3629 & n3633;
  assign n3635 = ~x301 & ~n3634;
  assign n3636 = x302 ^ x301;
  assign n3637 = n3626 & n3636;
  assign n3638 = x301 & x302;
  assign n3639 = n3624 & n3638;
  assign n3640 = x306 & n3639;
  assign n3641 = n3640 ^ n3638;
  assign n3642 = ~n3630 & n3641;
  assign n3643 = ~n3637 & ~n3642;
  assign n3644 = ~x302 & ~x306;
  assign n3645 = n3621 & n3644;
  assign n3646 = ~n3639 & ~n3645;
  assign n3647 = ~x305 & ~n3646;
  assign n3648 = n3643 & ~n3647;
  assign n3649 = ~n3635 & n3648;
  assign n3590 = ~x297 & ~x298;
  assign n3591 = ~x299 & ~x300;
  assign n3592 = ~n3590 & ~n3591;
  assign n3593 = x297 & x298;
  assign n3594 = x299 & x300;
  assign n3595 = ~n3593 & ~n3594;
  assign n3596 = n3592 & ~n3595;
  assign n3597 = x296 & n3596;
  assign n3598 = n3593 & n3594;
  assign n3599 = ~n3597 & ~n3598;
  assign n3600 = ~n3592 & n3595;
  assign n3601 = ~x296 & n3600;
  assign n3602 = n3590 & n3591;
  assign n3603 = ~n3601 & ~n3602;
  assign n3604 = n3599 & n3603;
  assign n3605 = ~x295 & ~n3604;
  assign n3606 = ~x296 & n3596;
  assign n3607 = x300 & n3593;
  assign n3608 = x296 & ~n3607;
  assign n3609 = ~n3600 & n3608;
  assign n3610 = ~n3606 & ~n3609;
  assign n3611 = x295 & ~n3610;
  assign n3612 = x295 & x296;
  assign n3613 = n3593 & n3612;
  assign n3614 = ~x296 & ~x300;
  assign n3615 = n3590 & n3614;
  assign n3616 = ~n3613 & ~n3615;
  assign n3617 = ~x299 & ~n3616;
  assign n3618 = ~n3611 & ~n3617;
  assign n3619 = ~n3605 & n3618;
  assign n3650 = n3649 ^ n3619;
  assign n3657 = x304 ^ x303;
  assign n3658 = n3657 ^ n3636;
  assign n3656 = x306 ^ x305;
  assign n3659 = n3658 ^ n3656;
  assign n3653 = x298 ^ x297;
  assign n3652 = x300 ^ x299;
  assign n3654 = n3653 ^ n3652;
  assign n3651 = x296 ^ x295;
  assign n3655 = n3654 ^ n3651;
  assign n3660 = n3659 ^ n3655;
  assign n3661 = n3587 ^ n3585;
  assign n3662 = n3661 ^ n3659;
  assign n3663 = ~n3660 & n3662;
  assign n3664 = n3663 ^ n3661;
  assign n3665 = ~n3650 & ~n3664;
  assign n3666 = ~n3589 & ~n3665;
  assign n3667 = n3655 & n3659;
  assign n3668 = n3667 ^ n3664;
  assign n3669 = ~n3588 & ~n3668;
  assign n3670 = n3669 ^ n3667;
  assign n3671 = n3670 ^ n3650;
  assign n3672 = ~n3581 & ~n3671;
  assign n3673 = n3650 & n3667;
  assign n3674 = ~n3672 & ~n3673;
  assign n3675 = n3666 & n3674;
  assign n3680 = n3599 & ~n3611;
  assign n3679 = n3629 & n3643;
  assign n3681 = n3680 ^ n3679;
  assign n3676 = n3667 ^ n3619;
  assign n3677 = n3650 & ~n3676;
  assign n3678 = n3677 ^ n3649;
  assign n3682 = n3681 ^ n3678;
  assign n3683 = n3565 & ~n3569;
  assign n3684 = ~n3682 & n3683;
  assign n3685 = ~n3675 & n3684;
  assign n3686 = ~n3522 & ~n3537;
  assign n3687 = n3588 ^ n3546;
  assign n3688 = n3581 & ~n3687;
  assign n3689 = n3688 ^ n3580;
  assign n3690 = ~n3686 & n3689;
  assign n3691 = n3685 & ~n3690;
  assign n3692 = n3680 ^ n3678;
  assign n3693 = ~n3681 & ~n3692;
  assign n3694 = n3693 ^ n3678;
  assign n3695 = ~n3691 & n3694;
  assign n3696 = n3682 & ~n3683;
  assign n3697 = n3675 & n3696;
  assign n3698 = ~n3695 & ~n3697;
  assign n3699 = n3683 ^ n3682;
  assign n3700 = n3682 ^ n3675;
  assign n3701 = n3699 & n3700;
  assign n3702 = n3701 ^ n3675;
  assign n3703 = n3690 & n3702;
  assign n3704 = n3698 & ~n3703;
  assign n3705 = n3699 ^ n3675;
  assign n3706 = n3686 & ~n3689;
  assign n3707 = ~n3705 & n3706;
  assign n3708 = ~n3704 & ~n3707;
  assign n4052 = x339 & x340;
  assign n4053 = x341 & x342;
  assign n4054 = ~n4052 & ~n4053;
  assign n4055 = ~x339 & ~x340;
  assign n4056 = ~x341 & ~x342;
  assign n4057 = ~n4055 & ~n4056;
  assign n4058 = ~n4054 & n4057;
  assign n4059 = x338 & n4058;
  assign n4060 = n4052 & n4053;
  assign n4061 = ~n4059 & ~n4060;
  assign n4062 = n4054 & ~n4057;
  assign n4066 = ~n4060 & ~n4062;
  assign n4067 = x338 & ~n4066;
  assign n4068 = ~x338 & ~n4058;
  assign n4069 = x337 & ~n4068;
  assign n4070 = ~n4067 & n4069;
  assign n4162 = n4061 & ~n4070;
  assign n4028 = x335 & x336;
  assign n4029 = x333 & x334;
  assign n4030 = ~n4028 & ~n4029;
  assign n4031 = ~x335 & ~x336;
  assign n4032 = ~x333 & ~x334;
  assign n4033 = ~n4031 & ~n4032;
  assign n4034 = ~n4030 & n4033;
  assign n4035 = x332 & n4034;
  assign n4036 = n4028 & n4029;
  assign n4037 = ~n4035 & ~n4036;
  assign n4038 = n4030 & ~n4033;
  assign n4042 = ~n4036 & ~n4038;
  assign n4043 = x332 & ~n4042;
  assign n4044 = ~x332 & ~n4034;
  assign n4045 = x331 & ~n4044;
  assign n4046 = ~n4043 & n4045;
  assign n4161 = n4037 & ~n4046;
  assign n4163 = n4162 ^ n4161;
  assign n4063 = ~x338 & n4062;
  assign n4064 = n4061 & ~n4063;
  assign n4065 = ~x337 & ~n4064;
  assign n3882 = x338 ^ x337;
  assign n4071 = n4055 & n4056;
  assign n4072 = n3882 & n4071;
  assign n4073 = ~n4070 & ~n4072;
  assign n4074 = ~n4065 & n4073;
  assign n3881 = x342 ^ x341;
  assign n3883 = n3882 ^ n3881;
  assign n3880 = x340 ^ x339;
  assign n3884 = n3883 ^ n3880;
  assign n3887 = x332 ^ x331;
  assign n3886 = x334 ^ x333;
  assign n3888 = n3887 ^ n3886;
  assign n3885 = x336 ^ x335;
  assign n3889 = n3888 ^ n3885;
  assign n4051 = n3884 & n3889;
  assign n4075 = n4074 ^ n4051;
  assign n4039 = ~x332 & n4038;
  assign n4040 = n4037 & ~n4039;
  assign n4041 = ~x331 & ~n4040;
  assign n4047 = n4031 & n4032;
  assign n4048 = n3887 & n4047;
  assign n4049 = ~n4046 & ~n4048;
  assign n4050 = ~n4041 & n4049;
  assign n4158 = n4051 ^ n4050;
  assign n4159 = n4075 & ~n4158;
  assign n4160 = n4159 ^ n4074;
  assign n4249 = n4162 ^ n4160;
  assign n4250 = ~n4163 & ~n4249;
  assign n4251 = n4250 ^ n4160;
  assign n4077 = x323 & x324;
  assign n4078 = x321 & x322;
  assign n4079 = ~n4077 & ~n4078;
  assign n4080 = ~x323 & ~x324;
  assign n4081 = ~x321 & ~x322;
  assign n4082 = ~n4080 & ~n4081;
  assign n4083 = ~n4079 & n4082;
  assign n4084 = x320 & n4083;
  assign n4085 = n4077 & n4078;
  assign n4086 = ~n4084 & ~n4085;
  assign n3876 = x320 ^ x319;
  assign n4093 = n3876 & n4083;
  assign n4087 = n4079 & ~n4082;
  assign n4094 = x319 & x320;
  assign n4095 = n4078 & n4094;
  assign n4096 = x324 & n4095;
  assign n4097 = n4096 ^ n4094;
  assign n4098 = ~n4087 & n4097;
  assign n4099 = ~n4093 & ~n4098;
  assign n4155 = n4086 & n4099;
  assign n4107 = x329 & x330;
  assign n4108 = x327 & x328;
  assign n4109 = ~n4107 & ~n4108;
  assign n4110 = ~x329 & ~x330;
  assign n4111 = ~x327 & ~x328;
  assign n4112 = ~n4110 & ~n4111;
  assign n4113 = ~n4109 & n4112;
  assign n4114 = x326 & n4113;
  assign n4115 = n4107 & n4108;
  assign n4116 = ~n4114 & ~n4115;
  assign n3871 = x326 ^ x325;
  assign n4123 = n3871 & n4113;
  assign n4117 = n4109 & ~n4112;
  assign n4124 = x325 & x326;
  assign n4125 = n4108 & n4124;
  assign n4126 = x330 & n4125;
  assign n4127 = n4126 ^ n4124;
  assign n4128 = ~n4117 & n4127;
  assign n4129 = ~n4123 & ~n4128;
  assign n4154 = n4116 & n4129;
  assign n4156 = n4155 ^ n4154;
  assign n4118 = ~x326 & n4117;
  assign n4119 = n4110 & n4111;
  assign n4120 = ~n4118 & ~n4119;
  assign n4121 = n4116 & n4120;
  assign n4122 = ~x325 & ~n4121;
  assign n4130 = ~x326 & ~x330;
  assign n4131 = n4111 & n4130;
  assign n4132 = ~n4125 & ~n4131;
  assign n4133 = ~x329 & ~n4132;
  assign n4134 = n4129 & ~n4133;
  assign n4135 = ~n4122 & n4134;
  assign n3870 = x328 ^ x327;
  assign n3872 = n3871 ^ n3870;
  assign n3869 = x330 ^ x329;
  assign n3873 = n3872 ^ n3869;
  assign n3875 = x322 ^ x321;
  assign n3877 = n3876 ^ n3875;
  assign n3874 = x324 ^ x323;
  assign n3878 = n3877 ^ n3874;
  assign n4106 = n3873 & n3878;
  assign n4136 = n4135 ^ n4106;
  assign n4088 = ~x320 & n4087;
  assign n4089 = n4080 & n4081;
  assign n4090 = ~n4088 & ~n4089;
  assign n4091 = n4086 & n4090;
  assign n4092 = ~x319 & ~n4091;
  assign n4100 = ~x320 & ~x324;
  assign n4101 = n4081 & n4100;
  assign n4102 = ~n4095 & ~n4101;
  assign n4103 = ~x323 & ~n4102;
  assign n4104 = n4099 & ~n4103;
  assign n4105 = ~n4092 & n4104;
  assign n4151 = n4106 ^ n4105;
  assign n4152 = n4136 & ~n4151;
  assign n4153 = n4152 ^ n4135;
  assign n4246 = n4155 ^ n4153;
  assign n4247 = ~n4156 & ~n4246;
  assign n4248 = n4247 ^ n4153;
  assign n4252 = n4251 ^ n4248;
  assign n4164 = n4163 ^ n4160;
  assign n4157 = n4156 ^ n4153;
  assign n4165 = n4164 ^ n4157;
  assign n4137 = n4136 ^ n4105;
  assign n4076 = n4075 ^ n4050;
  assign n4138 = n4137 ^ n4076;
  assign n3879 = n3878 ^ n3873;
  assign n3890 = n3889 ^ n3884;
  assign n3898 = n3879 & n3890;
  assign n4148 = n4076 ^ n3898;
  assign n4149 = n4138 & ~n4148;
  assign n4150 = n4149 ^ n4137;
  assign n4243 = n4157 ^ n4150;
  assign n4244 = n4165 & ~n4243;
  assign n4245 = n4244 ^ n4164;
  assign n4253 = n4252 ^ n4245;
  assign n3859 = x344 ^ x343;
  assign n3858 = x346 ^ x345;
  assign n3994 = x347 & x348;
  assign n3995 = n3994 ^ x346;
  assign n3996 = n3858 & ~n3995;
  assign n3997 = n3996 ^ x345;
  assign n3998 = n3859 & n3997;
  assign n3999 = ~x345 & ~x346;
  assign n4000 = ~n3994 & n3999;
  assign n4001 = x345 & x346;
  assign n4002 = x343 & x344;
  assign n4003 = ~n4001 & n4002;
  assign n4004 = ~n4000 & n4003;
  assign n4005 = ~n3998 & ~n4004;
  assign n4006 = ~x347 & ~x348;
  assign n4007 = ~n4005 & ~n4006;
  assign n4008 = n4001 & n4002;
  assign n4009 = ~x348 & n4008;
  assign n4010 = ~n4007 & ~n4009;
  assign n4011 = x344 & ~n4006;
  assign n4012 = n3994 & n4001;
  assign n4013 = ~n4011 & ~n4012;
  assign n4014 = n3997 & ~n4013;
  assign n4172 = n4010 & ~n4014;
  assign n3965 = x351 & x352;
  assign n3973 = x353 & x354;
  assign n3974 = ~n3965 & ~n3973;
  assign n3975 = ~x353 & ~x354;
  assign n3976 = ~x351 & ~x352;
  assign n3977 = ~n3975 & ~n3976;
  assign n3978 = n3974 & ~n3977;
  assign n3969 = x349 & x350;
  assign n3970 = n3965 & n3969;
  assign n3979 = x354 & n3970;
  assign n3980 = n3979 ^ n3969;
  assign n3981 = ~n3978 & n3980;
  assign n3864 = x350 ^ x349;
  assign n3982 = n3864 & ~n3974;
  assign n3983 = n3977 & n3982;
  assign n3984 = ~n3981 & ~n3983;
  assign n3862 = x354 ^ x353;
  assign n3986 = x353 ^ x350;
  assign n3987 = ~n3862 & n3986;
  assign n3988 = n3987 ^ x350;
  assign n4170 = n3965 & n3988;
  assign n4171 = n3984 & ~n4170;
  assign n4173 = n4172 ^ n4171;
  assign n3863 = x352 ^ x351;
  assign n3865 = n3864 ^ n3863;
  assign n3966 = ~x350 & ~x354;
  assign n3967 = ~n3965 & n3966;
  assign n3968 = n3865 & n3967;
  assign n3971 = ~n3968 & ~n3970;
  assign n3972 = ~x353 & ~n3971;
  assign n3985 = ~n3972 & n3984;
  assign n3989 = n3988 ^ x352;
  assign n3990 = ~n3863 & ~n3989;
  assign n3991 = ~x349 & n3990;
  assign n3992 = n3985 & ~n3991;
  assign n3860 = n3859 ^ n3858;
  assign n3857 = x348 ^ x347;
  assign n3861 = n3860 ^ n3857;
  assign n3866 = n3865 ^ n3862;
  assign n3964 = n3861 & n3866;
  assign n3993 = n3992 ^ n3964;
  assign n4015 = n4000 & ~n4011;
  assign n4016 = ~n4014 & ~n4015;
  assign n4017 = ~x343 & ~n4016;
  assign n4018 = n4010 & ~n4017;
  assign n4019 = ~x344 & ~x348;
  assign n4020 = ~n4001 & n4019;
  assign n4021 = n3860 & n4020;
  assign n4022 = ~n4008 & ~n4021;
  assign n4023 = ~x347 & ~n4022;
  assign n4024 = n4018 & ~n4023;
  assign n4167 = n4024 ^ n3992;
  assign n4168 = ~n3993 & n4167;
  assign n4169 = n4168 ^ n4024;
  assign n4238 = n4172 ^ n4169;
  assign n4239 = ~n4173 & ~n4238;
  assign n4240 = n4239 ^ n4169;
  assign n3904 = x365 & x366;
  assign n3905 = x363 & x364;
  assign n3906 = ~n3904 & ~n3905;
  assign n3907 = ~x365 & ~x366;
  assign n3908 = ~x363 & ~x364;
  assign n3909 = ~n3907 & ~n3908;
  assign n3910 = ~n3906 & n3909;
  assign n3911 = x362 & n3910;
  assign n3912 = n3904 & n3905;
  assign n3913 = ~n3911 & ~n3912;
  assign n3848 = x362 ^ x361;
  assign n3920 = n3848 & n3910;
  assign n3914 = n3906 & ~n3909;
  assign n3921 = x361 & x362;
  assign n3922 = n3905 & n3921;
  assign n3923 = x366 & n3922;
  assign n3924 = n3923 ^ n3921;
  assign n3925 = ~n3914 & n3924;
  assign n3926 = ~n3920 & ~n3925;
  assign n4182 = n3913 & n3926;
  assign n3933 = x359 & x360;
  assign n3934 = x357 & x358;
  assign n3935 = ~n3933 & ~n3934;
  assign n3936 = ~x359 & ~x360;
  assign n3937 = ~x357 & ~x358;
  assign n3938 = ~n3936 & ~n3937;
  assign n3939 = ~n3935 & n3938;
  assign n3940 = x356 & n3939;
  assign n3941 = n3933 & n3934;
  assign n3942 = ~n3940 & ~n3941;
  assign n3853 = x356 ^ x355;
  assign n3949 = n3853 & n3939;
  assign n3943 = n3935 & ~n3938;
  assign n3950 = x355 & x356;
  assign n3951 = n3934 & n3950;
  assign n3952 = x360 & n3951;
  assign n3953 = n3952 ^ n3950;
  assign n3954 = ~n3943 & n3953;
  assign n3955 = ~n3949 & ~n3954;
  assign n4181 = n3942 & n3955;
  assign n4183 = n4182 ^ n4181;
  assign n3944 = ~x356 & n3943;
  assign n3945 = n3936 & n3937;
  assign n3946 = ~n3944 & ~n3945;
  assign n3947 = n3942 & n3946;
  assign n3948 = ~x355 & ~n3947;
  assign n3956 = ~x356 & ~x360;
  assign n3957 = n3937 & n3956;
  assign n3958 = ~n3951 & ~n3957;
  assign n3959 = ~x359 & ~n3958;
  assign n3960 = n3955 & ~n3959;
  assign n3961 = ~n3948 & n3960;
  assign n3915 = ~x362 & n3914;
  assign n3916 = n3907 & n3908;
  assign n3917 = ~n3915 & ~n3916;
  assign n3918 = n3913 & n3917;
  assign n3919 = ~x361 & ~n3918;
  assign n3927 = ~x362 & ~x366;
  assign n3928 = n3908 & n3927;
  assign n3929 = ~n3922 & ~n3928;
  assign n3930 = ~x365 & ~n3929;
  assign n3931 = n3926 & ~n3930;
  assign n3932 = ~n3919 & n3931;
  assign n3962 = n3961 ^ n3932;
  assign n3847 = x364 ^ x363;
  assign n3849 = n3848 ^ n3847;
  assign n3846 = x366 ^ x365;
  assign n3850 = n3849 ^ n3846;
  assign n3852 = x358 ^ x357;
  assign n3854 = n3853 ^ n3852;
  assign n3851 = x360 ^ x359;
  assign n3855 = n3854 ^ n3851;
  assign n3901 = n3850 & n3855;
  assign n4178 = n3932 ^ n3901;
  assign n4179 = n3962 & ~n4178;
  assign n4180 = n4179 ^ n3961;
  assign n4235 = n4182 ^ n4180;
  assign n4236 = ~n4183 & ~n4235;
  assign n4237 = n4236 ^ n4180;
  assign n4241 = n4240 ^ n4237;
  assign n4184 = n4183 ^ n4180;
  assign n3856 = n3855 ^ n3850;
  assign n3867 = n3866 ^ n3861;
  assign n3902 = n3856 & n3867;
  assign n3903 = ~n3901 & ~n3902;
  assign n3963 = n3962 ^ n3903;
  assign n4025 = n4024 ^ n3993;
  assign n4175 = n4025 ^ n3902;
  assign n4176 = n3963 & n4175;
  assign n4177 = n4176 ^ n4025;
  assign n4185 = n4184 ^ n4177;
  assign n4174 = n4173 ^ n4169;
  assign n4232 = n4177 ^ n4174;
  assign n4233 = n4185 & ~n4232;
  assign n4234 = n4233 ^ n4184;
  assign n4242 = n4241 ^ n4234;
  assign n4254 = n4253 ^ n4242;
  assign n4186 = n4185 ^ n4174;
  assign n4166 = n4165 ^ n4150;
  assign n4187 = n4186 ^ n4166;
  assign n4143 = n4138 ^ n3898;
  assign n3868 = n3867 ^ n3856;
  assign n3891 = n3890 ^ n3879;
  assign n3899 = n3868 & n3891;
  assign n4144 = n4143 ^ n3899;
  assign n4026 = n4025 ^ n3963;
  assign n4145 = n4026 ^ n3899;
  assign n4146 = n4144 & n4145;
  assign n4147 = n4146 ^ n4143;
  assign n4229 = n4166 ^ n4147;
  assign n4230 = n4187 & ~n4229;
  assign n4231 = n4230 ^ n4186;
  assign n4255 = n4254 ^ n4231;
  assign n4188 = n4187 ^ n4147;
  assign n3840 = n3671 ^ n3581;
  assign n3804 = ~x275 & ~x276;
  assign n3805 = x272 & ~n3804;
  assign n3806 = x275 & x276;
  assign n3807 = x273 & x274;
  assign n3808 = n3806 & n3807;
  assign n3809 = ~n3805 & ~n3808;
  assign n3710 = x274 ^ x273;
  assign n3810 = n3806 ^ x274;
  assign n3811 = n3710 & ~n3810;
  assign n3812 = n3811 ^ x273;
  assign n3813 = ~n3809 & n3812;
  assign n3814 = ~x273 & ~x274;
  assign n3815 = ~n3806 & n3814;
  assign n3816 = ~n3805 & n3815;
  assign n3817 = ~n3813 & ~n3816;
  assign n3818 = ~x271 & ~n3817;
  assign n3819 = x271 & ~n3804;
  assign n3820 = n3812 & n3819;
  assign n3821 = x271 & x272;
  assign n3822 = ~n3820 & ~n3821;
  assign n3823 = ~n3804 & ~n3807;
  assign n3824 = ~n3815 & n3823;
  assign n3825 = ~x276 & n3807;
  assign n3826 = x272 & ~n3825;
  assign n3827 = ~n3824 & n3826;
  assign n3828 = ~n3822 & ~n3827;
  assign n3829 = ~n3818 & ~n3828;
  assign n3830 = x271 & ~n3814;
  assign n3831 = ~x272 & ~x276;
  assign n3832 = ~n3830 & n3831;
  assign n3833 = ~n3807 & ~n3832;
  assign n3834 = n3807 & ~n3821;
  assign n3835 = ~x275 & ~n3834;
  assign n3836 = ~n3833 & n3835;
  assign n3837 = n3829 & ~n3836;
  assign n3778 = x279 & x280;
  assign n3779 = x281 & x282;
  assign n3780 = ~n3778 & ~n3779;
  assign n3727 = x278 ^ x277;
  assign n3781 = ~x279 & ~x280;
  assign n3782 = n3727 & ~n3781;
  assign n3783 = ~n3780 & n3782;
  assign n3784 = ~n3779 & n3781;
  assign n3785 = x277 & x278;
  assign n3786 = ~n3778 & n3785;
  assign n3787 = ~n3784 & n3786;
  assign n3788 = ~n3783 & ~n3787;
  assign n3789 = ~x281 & ~x282;
  assign n3790 = ~n3788 & ~n3789;
  assign n3726 = x282 ^ x281;
  assign n3728 = n3727 ^ n3726;
  assign n3725 = x280 ^ x279;
  assign n3729 = n3728 ^ n3725;
  assign n3791 = ~x278 & ~n3778;
  assign n3792 = n3789 & n3791;
  assign n3793 = n3729 & n3792;
  assign n3794 = n3778 & n3785;
  assign n3795 = ~n3779 & n3794;
  assign n3796 = ~n3793 & ~n3795;
  assign n3797 = ~n3790 & n3796;
  assign n3798 = x278 & ~n3789;
  assign n3799 = n3784 & ~n3798;
  assign n3800 = n3778 & n3779;
  assign n3801 = ~n3799 & ~n3800;
  assign n3802 = ~x277 & ~n3801;
  assign n3803 = n3797 & ~n3802;
  assign n3838 = n3837 ^ n3803;
  assign n3722 = x290 ^ x289;
  assign n3756 = x291 & x292;
  assign n3757 = x293 & x294;
  assign n3758 = ~n3756 & ~n3757;
  assign n3759 = ~x291 & ~x292;
  assign n3760 = ~x293 & ~x294;
  assign n3761 = ~n3759 & ~n3760;
  assign n3762 = n3758 & ~n3761;
  assign n3763 = ~n3722 & n3762;
  assign n3764 = n3756 & n3757;
  assign n3765 = n3759 & n3760;
  assign n3766 = ~n3764 & ~n3765;
  assign n3767 = ~n3763 & n3766;
  assign n3768 = x289 & x290;
  assign n3769 = ~n3767 & ~n3768;
  assign n3770 = n3722 & n3761;
  assign n3771 = ~n3758 & n3770;
  assign n3772 = ~n3764 & n3768;
  assign n3773 = ~n3762 & n3772;
  assign n3774 = ~n3771 & ~n3773;
  assign n3775 = ~n3769 & n3774;
  assign n3716 = x284 ^ x283;
  assign n3736 = ~x285 & ~x286;
  assign n3737 = ~x287 & ~x288;
  assign n3738 = ~n3736 & ~n3737;
  assign n3739 = x285 & x286;
  assign n3740 = x287 & x288;
  assign n3741 = ~n3739 & ~n3740;
  assign n3742 = ~n3738 & n3741;
  assign n3743 = ~n3716 & n3742;
  assign n3744 = n3739 & n3740;
  assign n3745 = n3736 & n3737;
  assign n3746 = ~n3744 & ~n3745;
  assign n3747 = ~n3743 & n3746;
  assign n3748 = x283 & x284;
  assign n3749 = ~n3747 & ~n3748;
  assign n3750 = ~n3744 & n3748;
  assign n3751 = ~n3742 & n3750;
  assign n3752 = n3716 & n3738;
  assign n3753 = ~n3741 & n3752;
  assign n3754 = ~n3751 & ~n3753;
  assign n3755 = ~n3749 & n3754;
  assign n3776 = n3775 ^ n3755;
  assign n3715 = x286 ^ x285;
  assign n3717 = n3716 ^ n3715;
  assign n3714 = x288 ^ x287;
  assign n3718 = n3717 ^ n3714;
  assign n3711 = x276 ^ x275;
  assign n3712 = n3711 ^ n3710;
  assign n3709 = x272 ^ x271;
  assign n3713 = n3712 ^ n3709;
  assign n3719 = n3718 ^ n3713;
  assign n3721 = x292 ^ x291;
  assign n3723 = n3722 ^ n3721;
  assign n3720 = x294 ^ x293;
  assign n3724 = n3723 ^ n3720;
  assign n3730 = n3729 ^ n3724;
  assign n3731 = n3719 & n3730;
  assign n3733 = n3713 & n3718;
  assign n3732 = n3724 & n3729;
  assign n3734 = n3733 ^ n3732;
  assign n3735 = ~n3731 & ~n3734;
  assign n3777 = n3776 ^ n3735;
  assign n3839 = n3838 ^ n3777;
  assign n3841 = n3840 ^ n3839;
  assign n3842 = n3661 ^ n3660;
  assign n3843 = n3730 ^ n3719;
  assign n3844 = n3842 & n3843;
  assign n3845 = n3841 & n3844;
  assign n3892 = n3891 ^ n3868;
  assign n3893 = n3843 ^ n3842;
  assign n3894 = n3892 & n3893;
  assign n3895 = ~n3844 & ~n3894;
  assign n3896 = ~n3841 & n3895;
  assign n3897 = ~n3845 & ~n3896;
  assign n3900 = ~n3898 & ~n3899;
  assign n4027 = n4026 ^ n3900;
  assign n4139 = n4138 ^ n4027;
  assign n4140 = n3841 & n3894;
  assign n4141 = ~n4139 & ~n4140;
  assign n4142 = n3897 & ~n4141;
  assign n4189 = n4188 ^ n4142;
  assign n4212 = ~n3735 & n3776;
  assign n4213 = n3732 & n3733;
  assign n4214 = ~n4212 & ~n4213;
  assign n4215 = ~n3838 & ~n4214;
  assign n4205 = n3713 & n3729;
  assign n4216 = n3735 & ~n3776;
  assign n4217 = n3838 & ~n4216;
  assign n4218 = ~n4205 & n4217;
  assign n4219 = ~n4215 & ~n4218;
  assign n4197 = n3718 & n3724;
  assign n4220 = n3776 & n4197;
  assign n4221 = ~n4219 & ~n4220;
  assign n4209 = ~n3813 & ~n3828;
  assign n4206 = n4205 ^ n3803;
  assign n4207 = n3838 & ~n4206;
  assign n4208 = n4207 ^ n3837;
  assign n4210 = n4209 ^ n4208;
  assign n4202 = ~n3744 & n3754;
  assign n4201 = ~n3764 & n3774;
  assign n4203 = n4202 ^ n4201;
  assign n4198 = n4197 ^ n3755;
  assign n4199 = n3776 & ~n4198;
  assign n4200 = n4199 ^ n3775;
  assign n4204 = n4203 ^ n4200;
  assign n4211 = n4210 ^ n4204;
  assign n4222 = n4221 ^ n4211;
  assign n4195 = ~n3794 & ~n3800;
  assign n4196 = ~n3790 & n4195;
  assign n4223 = n4222 ^ n4196;
  assign n4192 = n3844 ^ n3839;
  assign n4193 = n3841 & n4192;
  assign n4194 = n4193 ^ n3840;
  assign n4224 = n4223 ^ n4194;
  assign n4190 = n3689 ^ n3686;
  assign n4191 = n4190 ^ n3705;
  assign n4225 = n4224 ^ n4191;
  assign n4226 = n4225 ^ n4188;
  assign n4227 = ~n4189 & ~n4226;
  assign n4228 = n4227 ^ n4225;
  assign n4256 = n4255 ^ n4228;
  assign n4277 = n3675 & n3682;
  assign n4278 = n3708 & n4277;
  assign n4279 = n3702 ^ n3689;
  assign n4280 = n4190 & ~n4279;
  assign n4281 = ~n3691 & n4280;
  assign n4282 = n4281 ^ n3691;
  assign n4283 = ~n4278 & ~n4282;
  assign n4284 = n4283 ^ n3694;
  assign n4263 = n4196 & ~n4222;
  assign n4264 = n4221 ^ n4208;
  assign n4265 = n4210 & n4264;
  assign n4266 = n4265 ^ n4221;
  assign n4267 = n4263 & ~n4266;
  assign n4268 = ~n4208 & n4209;
  assign n4269 = ~n4204 & n4268;
  assign n4270 = ~n4221 & n4269;
  assign n4271 = ~n4267 & ~n4270;
  assign n4272 = n4204 & n4266;
  assign n4273 = ~n4223 & n4272;
  assign n4274 = n4271 & ~n4273;
  assign n4260 = n4202 ^ n4200;
  assign n4261 = ~n4203 & ~n4260;
  assign n4262 = n4261 ^ n4200;
  assign n4275 = n4274 ^ n4262;
  assign n4257 = n4194 ^ n4191;
  assign n4258 = ~n4224 & n4257;
  assign n4259 = n4258 ^ n4223;
  assign n4276 = n4275 ^ n4259;
  assign n4285 = n4284 ^ n4276;
  assign n4286 = n4285 ^ n4228;
  assign n4287 = n4256 & ~n4286;
  assign n4288 = n4287 ^ n4285;
  assign n4289 = ~n4234 & ~n4253;
  assign n4290 = n4240 ^ n4231;
  assign n4291 = ~n4241 & n4290;
  assign n4292 = n4291 ^ n4231;
  assign n4293 = n4289 & ~n4292;
  assign n4294 = ~n4237 & ~n4240;
  assign n4295 = ~n4231 & n4294;
  assign n4296 = n4234 & n4253;
  assign n4297 = n4295 & ~n4296;
  assign n4298 = ~n4293 & ~n4297;
  assign n4299 = n4292 & n4296;
  assign n4300 = n4237 & n4240;
  assign n4301 = n4231 & n4300;
  assign n4302 = n4251 ^ n4245;
  assign n4303 = ~n4252 & n4302;
  assign n4304 = n4303 ^ n4245;
  assign n4305 = ~n4301 & ~n4304;
  assign n4306 = ~n4248 & ~n4251;
  assign n4307 = ~n4245 & n4306;
  assign n4308 = ~n4305 & ~n4307;
  assign n4309 = ~n4299 & ~n4308;
  assign n4310 = n4298 & ~n4309;
  assign n4314 = n4248 & n4251;
  assign n4315 = n4245 & n4314;
  assign n4316 = n4234 & n4315;
  assign n4317 = n4292 & n4316;
  assign n4318 = n4310 & ~n4317;
  assign n4311 = ~n4262 & ~n4273;
  assign n4312 = n4271 & ~n4311;
  assign n4313 = ~n4310 & n4312;
  assign n4319 = n4318 ^ n4313;
  assign n4320 = n4288 & n4319;
  assign n4321 = n4320 ^ n4318;
  assign n4322 = n4284 ^ n4275;
  assign n4323 = ~n4276 & n4322;
  assign n4324 = n4323 ^ n4284;
  assign n4325 = n4321 & ~n4324;
  assign n4326 = ~n4288 & n4313;
  assign n4327 = ~n4298 & ~n4304;
  assign n4328 = ~n4324 & n4327;
  assign n4329 = n4326 & ~n4328;
  assign n4330 = ~n4325 & ~n4329;
  assign n4331 = ~n3708 & ~n4330;
  assign n4333 = n4312 ^ n4288;
  assign n4332 = n4324 ^ n3708;
  assign n4334 = n4333 ^ n4332;
  assign n4335 = ~n4327 & n4334;
  assign n4336 = ~n4310 & ~n4335;
  assign n4337 = ~n4331 & ~n4336;
  assign n4338 = ~n3708 & ~n4324;
  assign n4339 = ~n4316 & n4338;
  assign n4340 = ~n4288 & n4339;
  assign n4341 = ~n4312 & ~n4340;
  assign n4342 = n3708 & n4324;
  assign n4343 = n4327 & ~n4342;
  assign n4344 = n4288 & ~n4338;
  assign n4345 = n4343 & ~n4344;
  assign n4346 = n4341 & ~n4345;
  assign n4347 = n4288 & n4342;
  assign n4348 = ~n4310 & ~n4347;
  assign n4349 = ~n4338 & ~n4348;
  assign n4350 = ~n4288 & n4318;
  assign n4351 = ~n4342 & n4350;
  assign n4352 = n4349 & ~n4351;
  assign n4353 = n4346 & ~n4352;
  assign n4354 = n4337 & ~n4353;
  assign n2892 = ~x395 & ~x396;
  assign n2893 = ~x393 & ~x394;
  assign n2894 = ~n2892 & ~n2893;
  assign n2895 = x395 & x396;
  assign n2896 = x393 & x394;
  assign n2897 = ~n2895 & ~n2896;
  assign n2898 = n2894 & ~n2897;
  assign n2899 = x392 & n2898;
  assign n2900 = n2895 & n2896;
  assign n2901 = ~n2899 & ~n2900;
  assign n2908 = x392 ^ x391;
  assign n2909 = n2898 & n2908;
  assign n2902 = ~n2894 & n2897;
  assign n2910 = x391 & x392;
  assign n2911 = n2896 & n2910;
  assign n2912 = x396 & n2911;
  assign n2913 = n2912 ^ n2910;
  assign n2914 = ~n2902 & n2913;
  assign n2915 = ~n2909 & ~n2914;
  assign n2933 = n2901 & n2915;
  assign n2864 = ~x401 & ~x402;
  assign n2861 = x401 & x402;
  assign n2867 = x399 & x400;
  assign n2884 = ~n2861 & ~n2867;
  assign n2862 = ~x399 & ~x400;
  assign n2872 = x398 ^ x397;
  assign n2885 = ~n2862 & n2872;
  assign n2886 = ~n2884 & n2885;
  assign n2863 = ~n2861 & n2862;
  assign n2879 = x397 & x398;
  assign n2887 = ~n2867 & n2879;
  assign n2888 = ~n2863 & n2887;
  assign n2889 = ~n2886 & ~n2888;
  assign n2890 = ~n2864 & ~n2889;
  assign n2868 = n2861 & n2867;
  assign n2880 = n2867 & n2879;
  assign n2931 = ~n2868 & ~n2880;
  assign n2932 = ~n2890 & n2931;
  assign n2934 = n2933 ^ n2932;
  assign n2903 = ~x392 & n2902;
  assign n2904 = n2892 & n2893;
  assign n2905 = ~n2903 & ~n2904;
  assign n2906 = n2901 & n2905;
  assign n2907 = ~x391 & ~n2906;
  assign n2916 = ~x392 & ~x396;
  assign n2917 = n2893 & n2916;
  assign n2918 = ~n2911 & ~n2917;
  assign n2919 = ~x395 & ~n2918;
  assign n2920 = n2915 & ~n2919;
  assign n2921 = ~n2907 & n2920;
  assign n2865 = x398 & ~n2864;
  assign n2866 = n2863 & ~n2865;
  assign n2869 = ~n2866 & ~n2868;
  assign n2870 = ~x397 & ~n2869;
  assign n2873 = x402 ^ x401;
  assign n2874 = n2873 ^ n2872;
  assign n2871 = x400 ^ x399;
  assign n2875 = n2874 ^ n2871;
  assign n2876 = ~x398 & n2864;
  assign n2877 = ~n2867 & n2876;
  assign n2878 = n2875 & n2877;
  assign n2881 = ~n2861 & n2880;
  assign n2882 = ~n2878 & ~n2881;
  assign n2883 = ~n2870 & n2882;
  assign n2891 = n2883 & ~n2890;
  assign n2922 = n2921 ^ n2891;
  assign n2924 = x394 ^ x393;
  assign n2925 = n2924 ^ n2908;
  assign n2923 = x396 ^ x395;
  assign n2926 = n2925 ^ n2923;
  assign n2927 = n2875 & n2926;
  assign n2928 = n2927 ^ n2891;
  assign n2929 = n2922 & ~n2928;
  assign n2930 = n2929 ^ n2921;
  assign n2935 = n2934 ^ n2930;
  assign n2936 = ~x413 & ~x414;
  assign n2937 = ~x411 & ~x412;
  assign n2938 = ~n2936 & ~n2937;
  assign n2939 = x413 & x414;
  assign n2940 = x411 & x412;
  assign n2941 = ~n2939 & ~n2940;
  assign n2942 = ~n2938 & n2941;
  assign n2945 = x414 ^ x413;
  assign n2944 = x412 ^ x411;
  assign n2946 = n2945 ^ n2944;
  assign n2943 = x410 ^ x409;
  assign n2947 = n2946 ^ n2943;
  assign n2948 = x409 & ~n2947;
  assign n2949 = ~n2942 & n2948;
  assign n2950 = x410 & n2938;
  assign n2951 = n2950 ^ n2939;
  assign n2952 = n2940 ^ n2939;
  assign n2953 = n2951 & ~n2952;
  assign n2954 = n2953 ^ n2950;
  assign n2955 = ~n2949 & ~n2954;
  assign n2956 = ~x407 & ~x408;
  assign n2957 = ~x405 & ~x406;
  assign n2958 = ~n2956 & ~n2957;
  assign n2959 = x407 & x408;
  assign n2960 = x405 & x406;
  assign n2961 = ~n2959 & ~n2960;
  assign n2962 = n2958 & ~n2961;
  assign n2963 = x404 & n2962;
  assign n2964 = n2959 & n2960;
  assign n2965 = ~n2963 & ~n2964;
  assign n2966 = x404 ^ x403;
  assign n2967 = n2962 & n2966;
  assign n2968 = ~n2958 & n2961;
  assign n2969 = x403 & x404;
  assign n2970 = n2960 & n2969;
  assign n2971 = x408 & n2970;
  assign n2972 = n2971 ^ n2969;
  assign n2973 = ~n2968 & n2972;
  assign n2974 = ~n2967 & ~n2973;
  assign n2975 = n2965 & n2974;
  assign n2976 = ~n2955 & ~n2975;
  assign n2977 = ~n2935 & ~n2976;
  assign n3003 = ~x410 & n2942;
  assign n3004 = n2936 & n2937;
  assign n3005 = ~n3003 & ~n3004;
  assign n3006 = ~n2954 & n3005;
  assign n3007 = ~n2948 & ~n3006;
  assign n3008 = n2939 & n2940;
  assign n3009 = n2949 & ~n3008;
  assign n3010 = ~n3007 & ~n3009;
  assign n2992 = ~x404 & n2968;
  assign n2993 = n2956 & n2957;
  assign n2994 = ~n2992 & ~n2993;
  assign n2995 = n2965 & n2994;
  assign n2996 = ~x403 & ~n2995;
  assign n2997 = ~x404 & ~x408;
  assign n2998 = n2957 & n2997;
  assign n2999 = ~n2970 & ~n2998;
  assign n3000 = ~x407 & ~n2999;
  assign n3001 = n2974 & ~n3000;
  assign n3002 = ~n2996 & n3001;
  assign n3011 = n3010 ^ n3002;
  assign n2988 = n2875 & n2947;
  assign n3012 = n3011 ^ n2988;
  assign n2983 = x406 ^ x405;
  assign n2984 = n2983 ^ n2966;
  assign n2982 = x408 ^ x407;
  assign n2985 = n2984 ^ n2982;
  assign n2989 = n2926 & n2985;
  assign n3013 = n3012 ^ n2989;
  assign n2981 = n2947 ^ n2875;
  assign n2986 = n2985 ^ n2926;
  assign n2987 = n2981 & n2986;
  assign n2990 = ~n2988 & ~n2989;
  assign n2991 = n2987 & n2990;
  assign n3014 = n3013 ^ n2991;
  assign n3015 = ~n2922 & n3014;
  assign n3016 = n2947 & n2985;
  assign n3017 = n3011 & n3016;
  assign n3018 = n2922 & n2927;
  assign n3019 = ~n3017 & ~n3018;
  assign n3020 = ~n3015 & n3019;
  assign n3021 = ~n2987 & n2990;
  assign n3022 = ~n3011 & n3021;
  assign n3023 = n3020 & ~n3022;
  assign n3024 = n3016 ^ n3002;
  assign n3025 = n3011 & ~n3024;
  assign n3026 = n3025 ^ n3010;
  assign n3027 = ~n3023 & ~n3026;
  assign n3028 = n2935 & ~n3027;
  assign n3029 = n2975 ^ n2955;
  assign n3030 = n3029 ^ n3026;
  assign n3031 = n3030 ^ n2935;
  assign n3032 = n3031 ^ n3023;
  assign n3033 = n2955 & n2975;
  assign n3034 = n3032 & n3033;
  assign n3035 = ~n3028 & n3034;
  assign n3036 = n3023 & n3026;
  assign n3037 = n2935 & ~n3033;
  assign n3038 = n3036 & n3037;
  assign n3039 = n3027 ^ n2976;
  assign n3040 = n2976 ^ n2935;
  assign n3041 = n3039 & ~n3040;
  assign n3042 = ~n3038 & n3041;
  assign n3043 = n3042 ^ n3038;
  assign n3044 = ~n3035 & ~n3043;
  assign n2978 = n2933 ^ n2930;
  assign n2979 = ~n2934 & ~n2978;
  assign n2980 = n2979 ^ n2930;
  assign n3045 = n3044 ^ n2980;
  assign n3046 = n2977 & n3045;
  assign n3047 = n2976 & n3028;
  assign n3048 = ~n2980 & ~n3036;
  assign n3049 = ~n3047 & n3048;
  assign n3050 = ~n3034 & ~n3049;
  assign n3051 = ~n3046 & n3050;
  assign n2705 = x389 & x390;
  assign n2706 = x387 & x388;
  assign n2707 = ~n2705 & ~n2706;
  assign n2708 = ~x389 & ~x390;
  assign n2709 = ~x387 & ~x388;
  assign n2710 = ~n2708 & ~n2709;
  assign n2711 = ~n2707 & n2710;
  assign n2712 = x386 & n2711;
  assign n2713 = n2705 & n2706;
  assign n2714 = ~n2712 & ~n2713;
  assign n2721 = x386 ^ x385;
  assign n2722 = n2711 & n2721;
  assign n2715 = n2707 & ~n2710;
  assign n2723 = x385 & x386;
  assign n2724 = n2706 & n2723;
  assign n2725 = x390 & n2724;
  assign n2726 = n2725 ^ n2723;
  assign n2727 = ~n2715 & n2726;
  assign n2728 = ~n2722 & ~n2727;
  assign n2749 = n2714 & n2728;
  assign n2686 = x381 & x382;
  assign n2687 = x383 & x384;
  assign n2691 = n2686 & n2687;
  assign n2683 = ~x381 & ~x382;
  assign n2684 = ~x383 & ~x384;
  assign n2685 = ~n2683 & ~n2684;
  assign n2688 = ~n2686 & ~n2687;
  assign n2694 = x380 ^ x379;
  assign n2695 = ~n2688 & n2694;
  assign n2696 = n2685 & n2695;
  assign n2689 = ~n2685 & n2688;
  assign n2697 = x379 & x380;
  assign n2698 = ~n2691 & n2697;
  assign n2699 = ~n2689 & n2698;
  assign n2700 = ~n2696 & ~n2699;
  assign n2748 = ~n2691 & n2700;
  assign n2750 = n2749 ^ n2748;
  assign n2716 = ~x386 & n2715;
  assign n2717 = n2708 & n2709;
  assign n2718 = ~n2716 & ~n2717;
  assign n2719 = n2714 & n2718;
  assign n2720 = ~x385 & ~n2719;
  assign n2729 = ~x386 & ~x390;
  assign n2730 = n2709 & n2729;
  assign n2731 = ~n2724 & ~n2730;
  assign n2732 = ~x389 & ~n2731;
  assign n2733 = n2728 & ~n2732;
  assign n2734 = ~n2720 & n2733;
  assign n2690 = ~x380 & n2689;
  assign n2692 = ~n2690 & ~n2691;
  assign n2693 = ~x379 & ~n2692;
  assign n2701 = n2683 & ~n2697;
  assign n2702 = n2684 & n2701;
  assign n2703 = n2700 & ~n2702;
  assign n2704 = ~n2693 & n2703;
  assign n2735 = n2734 ^ n2704;
  assign n2737 = x388 ^ x387;
  assign n2738 = n2737 ^ n2721;
  assign n2736 = x390 ^ x389;
  assign n2739 = n2738 ^ n2736;
  assign n2741 = x384 ^ x383;
  assign n2742 = n2741 ^ n2694;
  assign n2740 = x382 ^ x381;
  assign n2743 = n2742 ^ n2740;
  assign n2744 = n2739 & n2743;
  assign n2745 = n2744 ^ n2704;
  assign n2746 = n2735 & ~n2745;
  assign n2747 = n2746 ^ n2734;
  assign n2751 = n2750 ^ n2747;
  assign n2752 = ~x371 & ~x372;
  assign n2753 = ~x369 & ~x370;
  assign n2754 = ~n2752 & ~n2753;
  assign n2755 = x371 & x372;
  assign n2756 = x369 & x370;
  assign n2757 = ~n2755 & ~n2756;
  assign n2758 = n2754 & ~n2757;
  assign n2759 = x368 & n2758;
  assign n2760 = n2755 & n2756;
  assign n2761 = ~n2759 & ~n2760;
  assign n2762 = x368 ^ x367;
  assign n2763 = n2758 & n2762;
  assign n2764 = ~n2754 & n2757;
  assign n2765 = x367 & x368;
  assign n2766 = n2756 & n2765;
  assign n2767 = x372 & n2766;
  assign n2768 = n2767 ^ n2765;
  assign n2769 = ~n2764 & n2768;
  assign n2770 = ~n2763 & ~n2769;
  assign n2771 = n2761 & n2770;
  assign n2772 = n2751 & ~n2771;
  assign n2816 = n2743 ^ n2739;
  assign n2822 = x372 ^ x371;
  assign n2823 = n2822 ^ n2762;
  assign n2821 = x370 ^ x369;
  assign n2824 = n2823 ^ n2821;
  assign n2818 = x378 ^ x377;
  assign n2783 = x374 ^ x373;
  assign n2819 = n2818 ^ n2783;
  assign n2817 = x376 ^ x375;
  assign n2820 = n2819 ^ n2817;
  assign n2825 = n2824 ^ n2820;
  assign n2826 = n2816 & n2825;
  assign n2827 = n2820 & n2824;
  assign n2828 = n2827 ^ n2744;
  assign n2829 = ~n2826 & ~n2828;
  assign n2830 = n2829 ^ n2735;
  assign n2804 = ~x368 & n2764;
  assign n2805 = n2752 & n2753;
  assign n2806 = ~n2804 & ~n2805;
  assign n2807 = n2761 & n2806;
  assign n2808 = ~x367 & ~n2807;
  assign n2809 = ~x368 & ~x372;
  assign n2810 = n2753 & n2809;
  assign n2811 = ~n2766 & ~n2810;
  assign n2812 = ~x371 & ~n2811;
  assign n2813 = n2770 & ~n2812;
  assign n2814 = ~n2808 & n2813;
  assign n2773 = ~x377 & ~x378;
  assign n2774 = ~x375 & ~x376;
  assign n2775 = ~n2773 & ~n2774;
  assign n2776 = x377 & x378;
  assign n2777 = x375 & x376;
  assign n2778 = ~n2776 & ~n2777;
  assign n2779 = n2775 & ~n2778;
  assign n2780 = x374 & n2779;
  assign n2781 = n2776 & n2777;
  assign n2782 = ~n2780 & ~n2781;
  assign n2785 = ~n2775 & n2778;
  assign n2793 = ~x374 & n2785;
  assign n2794 = n2773 & n2774;
  assign n2795 = ~n2793 & ~n2794;
  assign n2796 = n2782 & n2795;
  assign n2797 = ~x373 & ~n2796;
  assign n2784 = n2779 & n2783;
  assign n2786 = x373 & x374;
  assign n2787 = n2777 & n2786;
  assign n2788 = x378 & n2787;
  assign n2789 = n2788 ^ n2786;
  assign n2790 = ~n2785 & n2789;
  assign n2791 = ~n2784 & ~n2790;
  assign n2798 = ~x374 & ~x378;
  assign n2799 = n2774 & n2798;
  assign n2800 = ~n2787 & ~n2799;
  assign n2801 = ~x377 & ~n2800;
  assign n2802 = n2791 & ~n2801;
  assign n2803 = ~n2797 & n2802;
  assign n2815 = n2814 ^ n2803;
  assign n2831 = n2830 ^ n2815;
  assign n2832 = ~n2815 & ~n2827;
  assign n2833 = n2831 & ~n2832;
  assign n2834 = ~n2735 & ~n2833;
  assign n2835 = ~n2815 & ~n2830;
  assign n2836 = n2735 & n2744;
  assign n2837 = n2815 & n2827;
  assign n2838 = ~n2836 & ~n2837;
  assign n2839 = ~n2835 & n2838;
  assign n2840 = ~n2834 & n2839;
  assign n2792 = n2782 & n2791;
  assign n2841 = n2840 ^ n2792;
  assign n2842 = n2827 ^ n2814;
  assign n2843 = ~n2815 & n2842;
  assign n2844 = n2843 ^ n2827;
  assign n2845 = n2844 ^ n2792;
  assign n2846 = ~n2841 & n2845;
  assign n2847 = n2846 ^ n2840;
  assign n2848 = ~n2772 & ~n2847;
  assign n2849 = n2844 ^ n2771;
  assign n2850 = n2849 ^ n2751;
  assign n2851 = n2850 ^ n2841;
  assign n2852 = ~n2751 & n2771;
  assign n2853 = ~n2851 & ~n2852;
  assign n2854 = n2848 & ~n2853;
  assign n2855 = n2847 & n2853;
  assign n2856 = n2749 ^ n2747;
  assign n2857 = ~n2750 & ~n2856;
  assign n2858 = n2857 ^ n2747;
  assign n2859 = ~n2855 & ~n2858;
  assign n2860 = ~n2854 & ~n2859;
  assign n3052 = n3051 ^ n2860;
  assign n3056 = n3014 ^ n2922;
  assign n3053 = n2986 ^ n2981;
  assign n3054 = n2825 ^ n2816;
  assign n3055 = n3053 & n3054;
  assign n3057 = n3056 ^ n3055;
  assign n3058 = n3056 ^ n2831;
  assign n3059 = ~n3057 & ~n3058;
  assign n3060 = n3059 ^ n2831;
  assign n3061 = n3060 ^ n2851;
  assign n3062 = n3060 ^ n3032;
  assign n3063 = ~n3061 & n3062;
  assign n3064 = n3063 ^ n2851;
  assign n3065 = n3064 ^ n3045;
  assign n3066 = ~n2854 & ~n2855;
  assign n3067 = n3066 ^ n2858;
  assign n3068 = n3067 ^ n3064;
  assign n3069 = ~n3065 & n3068;
  assign n3070 = n3069 ^ n3067;
  assign n3071 = n3070 ^ n3051;
  assign n3072 = ~n3052 & n3071;
  assign n3073 = n3072 ^ n3070;
  assign n3291 = x452 ^ x451;
  assign n3292 = x454 ^ x453;
  assign n3293 = x455 & x456;
  assign n3294 = n3293 ^ x454;
  assign n3295 = n3292 & ~n3294;
  assign n3296 = n3295 ^ x453;
  assign n3297 = n3291 & n3296;
  assign n3298 = ~x453 & ~x454;
  assign n3299 = ~n3293 & n3298;
  assign n3300 = x453 & x454;
  assign n3301 = x451 & x452;
  assign n3302 = ~n3300 & n3301;
  assign n3303 = ~n3299 & n3302;
  assign n3304 = ~n3297 & ~n3303;
  assign n3305 = ~x455 & ~x456;
  assign n3306 = ~n3304 & ~n3305;
  assign n3307 = n3300 & n3301;
  assign n3308 = ~x456 & n3307;
  assign n3309 = ~n3306 & ~n3308;
  assign n3310 = x452 & ~n3305;
  assign n3311 = n3293 & n3300;
  assign n3312 = ~n3310 & ~n3311;
  assign n3313 = n3296 & ~n3312;
  assign n3314 = n3299 & ~n3310;
  assign n3315 = ~x452 & ~n3300;
  assign n3316 = n3305 & n3315;
  assign n3317 = ~n3314 & ~n3316;
  assign n3318 = ~n3313 & n3317;
  assign n3319 = ~x451 & ~n3318;
  assign n3320 = ~x452 & ~x456;
  assign n3321 = n3298 & n3320;
  assign n3322 = ~n3307 & ~n3321;
  assign n3323 = ~x455 & ~n3322;
  assign n3324 = ~n3319 & ~n3323;
  assign n3325 = n3309 & n3324;
  assign n3256 = x458 ^ x457;
  assign n3257 = x460 ^ x459;
  assign n3258 = x461 & x462;
  assign n3259 = n3258 ^ x460;
  assign n3260 = n3257 & ~n3259;
  assign n3261 = n3260 ^ x459;
  assign n3262 = n3256 & n3261;
  assign n3263 = ~x459 & ~x460;
  assign n3264 = ~n3258 & n3263;
  assign n3265 = x459 & x460;
  assign n3266 = x457 & x458;
  assign n3267 = ~n3265 & n3266;
  assign n3268 = ~n3264 & n3267;
  assign n3269 = ~n3262 & ~n3268;
  assign n3270 = ~x461 & ~x462;
  assign n3271 = ~n3269 & ~n3270;
  assign n3272 = n3265 & n3266;
  assign n3273 = ~x462 & n3272;
  assign n3274 = ~n3271 & ~n3273;
  assign n3275 = x458 & ~n3270;
  assign n3276 = n3258 & n3265;
  assign n3277 = ~n3275 & ~n3276;
  assign n3278 = n3261 & ~n3277;
  assign n3279 = n3264 & ~n3275;
  assign n3280 = ~x458 & ~n3265;
  assign n3281 = n3270 & n3280;
  assign n3282 = ~n3279 & ~n3281;
  assign n3283 = ~n3278 & n3282;
  assign n3284 = ~x457 & ~n3283;
  assign n3285 = ~x458 & ~x462;
  assign n3286 = n3263 & n3285;
  assign n3287 = ~n3272 & ~n3286;
  assign n3288 = ~x461 & ~n3287;
  assign n3289 = ~n3284 & ~n3288;
  assign n3290 = n3274 & n3289;
  assign n3326 = n3325 ^ n3290;
  assign n3327 = x456 ^ x455;
  assign n3328 = n3327 ^ n3291;
  assign n3329 = n3328 ^ n3292;
  assign n3330 = x462 ^ x461;
  assign n3331 = n3330 ^ n3256;
  assign n3332 = n3331 ^ n3257;
  assign n3333 = n3329 & n3332;
  assign n3334 = n3333 ^ n3325;
  assign n3335 = ~n3326 & n3334;
  assign n3336 = n3335 ^ n3333;
  assign n3430 = n3332 ^ n3329;
  assign n3417 = x444 ^ x443;
  assign n3345 = x442 ^ x441;
  assign n3418 = n3417 ^ n3345;
  assign n3416 = x440 ^ x439;
  assign n3419 = n3418 ^ n3416;
  assign n3413 = x450 ^ x449;
  assign n3381 = x448 ^ x447;
  assign n3414 = n3413 ^ n3381;
  assign n3412 = x446 ^ x445;
  assign n3415 = n3414 ^ n3412;
  assign n3431 = n3419 ^ n3415;
  assign n3432 = n3430 & n3431;
  assign n3420 = n3415 & n3419;
  assign n3433 = n3420 ^ n3333;
  assign n3434 = ~n3432 & ~n3433;
  assign n3375 = x449 & x450;
  assign n3376 = x447 & x448;
  assign n3377 = n3375 & n3376;
  assign n3378 = ~x449 & ~x450;
  assign n3379 = x446 & ~n3378;
  assign n3380 = ~n3377 & ~n3379;
  assign n3382 = n3375 ^ x448;
  assign n3383 = n3381 & ~n3382;
  assign n3384 = n3383 ^ x447;
  assign n3385 = ~n3380 & n3384;
  assign n3386 = ~x447 & ~x448;
  assign n3387 = ~n3375 & n3386;
  assign n3388 = ~n3379 & n3387;
  assign n3389 = ~x446 & ~n3376;
  assign n3390 = n3378 & n3389;
  assign n3391 = ~n3388 & ~n3390;
  assign n3392 = ~n3385 & n3391;
  assign n3393 = ~x445 & ~n3392;
  assign n3394 = x445 & ~n3378;
  assign n3395 = n3384 & n3394;
  assign n3396 = x445 & x446;
  assign n3397 = ~n3395 & ~n3396;
  assign n3398 = ~n3376 & ~n3378;
  assign n3399 = ~n3387 & n3398;
  assign n3400 = ~x450 & n3376;
  assign n3401 = x446 & ~n3400;
  assign n3402 = ~n3399 & n3401;
  assign n3403 = ~n3397 & ~n3402;
  assign n3404 = ~n3393 & ~n3403;
  assign n3405 = n3376 & n3396;
  assign n3406 = ~x446 & ~x450;
  assign n3407 = n3386 & n3406;
  assign n3408 = ~n3405 & ~n3407;
  assign n3409 = ~x449 & ~n3408;
  assign n3410 = n3404 & ~n3409;
  assign n3339 = x443 & x444;
  assign n3340 = x441 & x442;
  assign n3341 = n3339 & n3340;
  assign n3342 = ~x443 & ~x444;
  assign n3343 = x440 & ~n3342;
  assign n3344 = ~n3341 & ~n3343;
  assign n3346 = n3339 ^ x442;
  assign n3347 = n3345 & ~n3346;
  assign n3348 = n3347 ^ x441;
  assign n3349 = ~n3344 & n3348;
  assign n3350 = ~x441 & ~x442;
  assign n3351 = ~n3339 & n3350;
  assign n3352 = ~n3343 & n3351;
  assign n3353 = ~x440 & ~n3340;
  assign n3354 = n3342 & n3353;
  assign n3355 = ~n3352 & ~n3354;
  assign n3356 = ~n3349 & n3355;
  assign n3357 = ~x439 & ~n3356;
  assign n3358 = x439 & ~n3342;
  assign n3359 = n3348 & n3358;
  assign n3360 = x439 & x440;
  assign n3361 = ~n3359 & ~n3360;
  assign n3362 = ~n3340 & ~n3342;
  assign n3363 = ~n3351 & n3362;
  assign n3364 = ~x444 & n3340;
  assign n3365 = x440 & ~n3364;
  assign n3366 = ~n3363 & n3365;
  assign n3367 = ~n3361 & ~n3366;
  assign n3368 = ~n3357 & ~n3367;
  assign n3369 = n3340 & n3360;
  assign n3370 = ~x440 & ~x444;
  assign n3371 = n3350 & n3370;
  assign n3372 = ~n3369 & ~n3371;
  assign n3373 = ~x443 & ~n3372;
  assign n3374 = n3368 & ~n3373;
  assign n3411 = n3410 ^ n3374;
  assign n3435 = n3434 ^ n3411;
  assign n3436 = n3435 ^ n3326;
  assign n3437 = n3326 & ~n3333;
  assign n3438 = ~n3436 & ~n3437;
  assign n3439 = n3420 ^ n3411;
  assign n3440 = ~n3432 & ~n3439;
  assign n3441 = ~n3438 & ~n3440;
  assign n3429 = n3274 & ~n3278;
  assign n3442 = n3441 ^ n3429;
  assign n3425 = ~n3349 & ~n3367;
  assign n3424 = ~n3385 & ~n3403;
  assign n3426 = n3425 ^ n3424;
  assign n3421 = n3420 ^ n3374;
  assign n3422 = n3411 & ~n3421;
  assign n3423 = n3422 ^ n3410;
  assign n3427 = n3426 ^ n3423;
  assign n3337 = n3309 & ~n3313;
  assign n3338 = n3337 ^ n3336;
  assign n3428 = n3427 ^ n3338;
  assign n3443 = n3442 ^ n3428;
  assign n3444 = ~n3336 & n3443;
  assign n3445 = n3429 ^ n3337;
  assign n3446 = ~n3442 & ~n3445;
  assign n3447 = n3446 ^ n3441;
  assign n3448 = n3444 & ~n3447;
  assign n3449 = n3429 & ~n3441;
  assign n3450 = n3337 & ~n3427;
  assign n3451 = n3449 & n3450;
  assign n3452 = ~n3448 & ~n3451;
  assign n3453 = n3427 & n3447;
  assign n3454 = ~n3443 & n3453;
  assign n3455 = n3425 ^ n3423;
  assign n3456 = ~n3426 & ~n3455;
  assign n3457 = n3456 ^ n3423;
  assign n3458 = ~n3454 & ~n3457;
  assign n3459 = n3452 & ~n3458;
  assign n3074 = x423 & x424;
  assign n3079 = x425 & x426;
  assign n3084 = n3074 & n3079;
  assign n3087 = x422 ^ x421;
  assign n3078 = ~x423 & ~x424;
  assign n3088 = ~n3078 & n3079;
  assign n3075 = ~x425 & ~x426;
  assign n3089 = n3074 & ~n3075;
  assign n3090 = ~n3088 & ~n3089;
  assign n3091 = n3087 & ~n3090;
  assign n3080 = n3078 & ~n3079;
  assign n3092 = x421 & x422;
  assign n3093 = ~n3080 & n3092;
  assign n3076 = ~n3074 & n3075;
  assign n3094 = ~n3076 & ~n3084;
  assign n3095 = n3093 & n3094;
  assign n3096 = ~n3091 & ~n3095;
  assign n3142 = ~n3084 & n3096;
  assign n3103 = ~x419 & ~x420;
  assign n3100 = x419 & x420;
  assign n3106 = x417 & x418;
  assign n3121 = ~n3100 & ~n3106;
  assign n3101 = ~x417 & ~x418;
  assign n3111 = x416 ^ x415;
  assign n3122 = ~n3101 & n3111;
  assign n3123 = ~n3121 & n3122;
  assign n3102 = ~n3100 & n3101;
  assign n3116 = x415 & x416;
  assign n3124 = ~n3106 & n3116;
  assign n3125 = ~n3102 & n3124;
  assign n3126 = ~n3123 & ~n3125;
  assign n3127 = ~n3103 & ~n3126;
  assign n3107 = n3100 & n3106;
  assign n3117 = n3106 & n3116;
  assign n3140 = ~n3107 & ~n3117;
  assign n3141 = ~n3127 & n3140;
  assign n3143 = n3142 ^ n3141;
  assign n3104 = x416 & ~n3103;
  assign n3105 = n3102 & ~n3104;
  assign n3108 = ~n3105 & ~n3107;
  assign n3109 = ~x415 & ~n3108;
  assign n3110 = x418 ^ x417;
  assign n3112 = n3111 ^ n3110;
  assign n3113 = ~x416 & n3103;
  assign n3114 = ~n3106 & n3113;
  assign n3115 = n3112 & n3114;
  assign n3118 = ~n3100 & n3117;
  assign n3119 = ~n3115 & ~n3118;
  assign n3120 = ~n3109 & n3119;
  assign n3128 = n3120 & ~n3127;
  assign n3077 = ~x422 & n3076;
  assign n3081 = x422 & ~n3075;
  assign n3082 = n3080 & ~n3081;
  assign n3083 = ~n3077 & ~n3082;
  assign n3085 = n3083 & ~n3084;
  assign n3086 = ~x421 & ~n3085;
  assign n3097 = n3077 & n3078;
  assign n3098 = n3096 & ~n3097;
  assign n3099 = ~n3086 & n3098;
  assign n3129 = n3128 ^ n3099;
  assign n3131 = x426 ^ x425;
  assign n3132 = n3131 ^ n3087;
  assign n3130 = x424 ^ x423;
  assign n3133 = n3132 ^ n3130;
  assign n3134 = x420 ^ x419;
  assign n3135 = n3134 ^ n3112;
  assign n3136 = n3133 & n3135;
  assign n3137 = n3136 ^ n3128;
  assign n3138 = ~n3129 & n3137;
  assign n3139 = n3138 ^ n3136;
  assign n3144 = n3143 ^ n3139;
  assign n3220 = x438 ^ x437;
  assign n3192 = x434 ^ x433;
  assign n3191 = x436 ^ x435;
  assign n3193 = n3192 ^ n3191;
  assign n3221 = n3220 ^ n3193;
  assign n3218 = x432 ^ x431;
  assign n3209 = x428 ^ x427;
  assign n3208 = x430 ^ x429;
  assign n3210 = n3209 ^ n3208;
  assign n3219 = n3218 ^ n3210;
  assign n3226 = n3221 ^ n3219;
  assign n3227 = n3135 ^ n3133;
  assign n3228 = n3227 ^ n3219;
  assign n3229 = ~n3226 & n3228;
  assign n3230 = n3229 ^ n3227;
  assign n3222 = n3219 & n3221;
  assign n3231 = n3230 ^ n3222;
  assign n3232 = ~n3136 & ~n3231;
  assign n3233 = n3232 ^ n3222;
  assign n3234 = n3233 ^ n3129;
  assign n3164 = x431 & x432;
  assign n3165 = x429 & x430;
  assign n3166 = ~n3164 & ~n3165;
  assign n3167 = ~x431 & ~x432;
  assign n3168 = ~x429 & ~x430;
  assign n3169 = ~n3167 & ~n3168;
  assign n3170 = n3166 & ~n3169;
  assign n3171 = x427 & x428;
  assign n3172 = n3165 & n3171;
  assign n3173 = x432 & n3172;
  assign n3174 = n3173 ^ n3171;
  assign n3175 = ~n3170 & n3174;
  assign n3176 = n3164 & n3165;
  assign n3177 = ~n3175 & ~n3176;
  assign n3178 = ~n3166 & n3169;
  assign n3179 = ~x428 & n3178;
  assign n3180 = ~x427 & n3179;
  assign n3181 = n3180 ^ n3178;
  assign n3182 = n3177 & ~n3181;
  assign n3201 = x428 & ~n3167;
  assign n3202 = ~n3164 & n3168;
  assign n3203 = ~n3201 & n3202;
  assign n3204 = n3182 & ~n3203;
  assign n3205 = x427 & ~n3175;
  assign n3206 = ~n3179 & n3205;
  assign n3207 = ~n3204 & ~n3206;
  assign n3211 = ~x428 & ~x432;
  assign n3212 = ~n3165 & n3211;
  assign n3213 = n3210 & n3212;
  assign n3214 = ~n3172 & ~n3213;
  assign n3215 = ~x431 & ~n3214;
  assign n3216 = ~n3207 & ~n3215;
  assign n3145 = x437 & x438;
  assign n3146 = x435 & x436;
  assign n3147 = n3145 & n3146;
  assign n3148 = ~n3145 & ~n3146;
  assign n3149 = ~x437 & ~x438;
  assign n3150 = ~x435 & ~x436;
  assign n3151 = ~n3149 & ~n3150;
  assign n3152 = ~n3148 & n3151;
  assign n3153 = ~x434 & n3152;
  assign n3154 = ~x433 & n3153;
  assign n3155 = n3154 ^ n3152;
  assign n3156 = ~n3147 & ~n3155;
  assign n3185 = x434 & ~n3149;
  assign n3186 = ~n3145 & n3150;
  assign n3187 = ~n3185 & n3186;
  assign n3188 = n3156 & ~n3187;
  assign n3189 = x433 & ~n3153;
  assign n3190 = ~n3188 & ~n3189;
  assign n3157 = n3148 & ~n3151;
  assign n3158 = x433 & x434;
  assign n3159 = n3146 & n3158;
  assign n3160 = x438 & n3159;
  assign n3161 = n3160 ^ n3158;
  assign n3162 = ~n3157 & n3161;
  assign n3194 = ~x434 & ~x438;
  assign n3195 = ~n3146 & n3194;
  assign n3196 = n3193 & n3195;
  assign n3197 = ~n3159 & ~n3196;
  assign n3198 = ~x437 & ~n3197;
  assign n3199 = ~n3162 & ~n3198;
  assign n3200 = ~n3190 & n3199;
  assign n3217 = n3216 ^ n3200;
  assign n3235 = n3234 ^ n3217;
  assign n3236 = n3129 & ~n3136;
  assign n3237 = ~n3235 & ~n3236;
  assign n3238 = ~n3217 & ~n3231;
  assign n3239 = n3238 ^ n3222;
  assign n3240 = ~n3237 & ~n3239;
  assign n3223 = n3217 & ~n3222;
  assign n3224 = ~n3200 & ~n3216;
  assign n3225 = ~n3223 & ~n3224;
  assign n3241 = n3240 ^ n3225;
  assign n3163 = n3156 & ~n3162;
  assign n3183 = n3182 ^ n3163;
  assign n3184 = n3183 ^ n3144;
  assign n3242 = n3241 ^ n3184;
  assign n3243 = n3144 & ~n3242;
  assign n3244 = n3225 & n3240;
  assign n3245 = ~n3163 & ~n3182;
  assign n3246 = ~n3244 & ~n3245;
  assign n3247 = n3183 & n3241;
  assign n3248 = n3246 & ~n3247;
  assign n3249 = ~n3243 & n3248;
  assign n3250 = n3243 & ~n3246;
  assign n3251 = n3142 ^ n3139;
  assign n3252 = ~n3143 & ~n3251;
  assign n3253 = n3252 ^ n3139;
  assign n3254 = ~n3250 & ~n3253;
  assign n3255 = ~n3249 & ~n3254;
  assign n3460 = n3459 ^ n3255;
  assign n3472 = ~n3249 & ~n3250;
  assign n3473 = n3472 ^ n3253;
  assign n3461 = n3431 ^ n3430;
  assign n3462 = n3227 ^ n3226;
  assign n3463 = n3461 & n3462;
  assign n3464 = n3463 ^ n3235;
  assign n3465 = n3463 ^ n3436;
  assign n3466 = ~n3464 & n3465;
  assign n3467 = n3466 ^ n3235;
  assign n3468 = n3467 ^ n3242;
  assign n3469 = n3467 ^ n3443;
  assign n3470 = ~n3468 & n3469;
  assign n3471 = n3470 ^ n3242;
  assign n3474 = n3473 ^ n3471;
  assign n3475 = n3452 & ~n3454;
  assign n3476 = n3475 ^ n3457;
  assign n3477 = n3476 ^ n3471;
  assign n3478 = n3474 & ~n3477;
  assign n3479 = n3478 ^ n3473;
  assign n3480 = n3479 ^ n3459;
  assign n3481 = ~n3460 & n3480;
  assign n3482 = n3481 ^ n3479;
  assign n3483 = n3073 & n3482;
  assign n3485 = n3070 ^ n3052;
  assign n3484 = n3479 ^ n3460;
  assign n3486 = n3485 ^ n3484;
  assign n3502 = n3476 ^ n3474;
  assign n3496 = n3468 ^ n3443;
  assign n3490 = n3057 ^ n2831;
  assign n3487 = n3054 ^ n3053;
  assign n3488 = n3462 ^ n3461;
  assign n3489 = n3487 & n3488;
  assign n3491 = n3490 ^ n3489;
  assign n3492 = n3464 ^ n3436;
  assign n3493 = n3492 ^ n3489;
  assign n3494 = ~n3491 & ~n3493;
  assign n3495 = n3494 ^ n3490;
  assign n3497 = n3496 ^ n3495;
  assign n3498 = n3061 ^ n3032;
  assign n3499 = n3498 ^ n3496;
  assign n3500 = ~n3497 & n3499;
  assign n3501 = n3500 ^ n3498;
  assign n3503 = n3502 ^ n3501;
  assign n3504 = n3067 ^ n3065;
  assign n3505 = n3504 ^ n3501;
  assign n3506 = ~n3503 & n3505;
  assign n3507 = n3506 ^ n3502;
  assign n3508 = n3507 ^ n3484;
  assign n3509 = n3486 & ~n3508;
  assign n3510 = n3509 ^ n3485;
  assign n3511 = n3483 & n3510;
  assign n4355 = n4354 ^ n3511;
  assign n4356 = n3708 & n4288;
  assign n4357 = n4313 & n4324;
  assign n4358 = ~n4356 & ~n4357;
  assign n4359 = n4327 & ~n4358;
  assign n4360 = n3708 & ~n4324;
  assign n4361 = n4326 & n4360;
  assign n4362 = n4312 & n4317;
  assign n4363 = n4342 & n4362;
  assign n4364 = ~n4361 & ~n4363;
  assign n4365 = ~n4359 & n4364;
  assign n4366 = ~n4331 & n4365;
  assign n4367 = ~n4353 & n4366;
  assign n4368 = ~n4355 & ~n4367;
  assign n4393 = n3507 ^ n3486;
  assign n4387 = n3504 ^ n3503;
  assign n4381 = n3498 ^ n3497;
  assign n4373 = n3492 ^ n3490;
  assign n4369 = n3893 ^ n3892;
  assign n4370 = n3488 ^ n3487;
  assign n4371 = n4369 & n4370;
  assign n4372 = ~n3489 & ~n4371;
  assign n4374 = n4373 ^ n4372;
  assign n4375 = n3895 ^ n3841;
  assign n4376 = n4375 ^ n4139;
  assign n4377 = n4374 & ~n4376;
  assign n4378 = n4373 & n4376;
  assign n4379 = n4371 & ~n4378;
  assign n4380 = ~n4377 & ~n4379;
  assign n4382 = n4381 ^ n4380;
  assign n4383 = n4225 ^ n4189;
  assign n4384 = n4383 ^ n4380;
  assign n4385 = n4382 & ~n4384;
  assign n4386 = n4385 ^ n4381;
  assign n4388 = n4387 ^ n4386;
  assign n4389 = n4285 ^ n4256;
  assign n4390 = n4389 ^ n4386;
  assign n4391 = n4388 & ~n4390;
  assign n4392 = n4391 ^ n4387;
  assign n4394 = n4393 ^ n4392;
  assign n4395 = ~n4318 & ~n4327;
  assign n4396 = n4395 ^ n4334;
  assign n4397 = n4396 ^ n4393;
  assign n4398 = n4394 & n4397;
  assign n4399 = n4398 ^ n4396;
  assign n4404 = ~n3073 & ~n3482;
  assign n4405 = ~n3510 & n4404;
  assign n4400 = n3482 ^ n3073;
  assign n4401 = n3510 ^ n3073;
  assign n4402 = ~n4400 & n4401;
  assign n4403 = n4402 ^ n3510;
  assign n4406 = n4405 ^ n4403;
  assign n4407 = n4399 & n4406;
  assign n4408 = n4407 ^ n4405;
  assign n4409 = n4368 & ~n4408;
  assign n4410 = ~n4366 & ~n4405;
  assign n4411 = ~n4353 & ~n4410;
  assign n4412 = ~n4399 & ~n4403;
  assign n4413 = ~n4405 & ~n4412;
  assign n4414 = n4413 ^ n4337;
  assign n4415 = n4411 & n4414;
  assign n4416 = ~n4409 & ~n4415;
  assign n4446 = n2675 ^ n2647;
  assign n4419 = n4396 ^ n4394;
  assign n4417 = n2672 ^ n2620;
  assign n4418 = n4417 ^ n2648;
  assign n4420 = n4419 ^ n4418;
  assign n4437 = n2669 ^ n2668;
  assign n4431 = n4383 ^ n4382;
  assign n4425 = n2658 ^ n2655;
  assign n4421 = n4370 ^ n4369;
  assign n4422 = n2579 ^ n2578;
  assign n4423 = n4422 ^ n2650;
  assign n4424 = n4421 & n4423;
  assign n4426 = n4425 ^ n4424;
  assign n4427 = n4376 ^ n4374;
  assign n4428 = n4427 ^ n4424;
  assign n4429 = ~n4426 & n4428;
  assign n4430 = n4429 ^ n4425;
  assign n4432 = n4431 ^ n4430;
  assign n4433 = n2663 ^ n2662;
  assign n4434 = n4433 ^ n4430;
  assign n4435 = n4432 & ~n4434;
  assign n4436 = n4435 ^ n4431;
  assign n4438 = n4437 ^ n4436;
  assign n4439 = n4389 ^ n4388;
  assign n4440 = n4439 ^ n4436;
  assign n4441 = n4438 & ~n4440;
  assign n4442 = n4441 ^ n4437;
  assign n4443 = n4442 ^ n4418;
  assign n4444 = ~n4420 & n4443;
  assign n4445 = n4444 ^ n4419;
  assign n4447 = n4446 ^ n4445;
  assign n4449 = n4399 ^ n4367;
  assign n4448 = n4400 ^ n3510;
  assign n4450 = n4449 ^ n4448;
  assign n4451 = n4450 ^ n4446;
  assign n4452 = n4447 & ~n4451;
  assign n4453 = n4452 ^ n4450;
  assign n4454 = ~n4416 & ~n4453;
  assign n4455 = n2682 & ~n4454;
  assign n4456 = ~n4354 & n4409;
  assign n4457 = n4337 & ~n4412;
  assign n4458 = n4367 & ~n4457;
  assign n4459 = ~n4405 & ~n4458;
  assign n4460 = ~n4456 & n4459;
  assign n4461 = ~n4454 & ~n4460;
  assign n4462 = ~n4455 & ~n4461;
  assign n4463 = n4416 & n4453;
  assign n4464 = ~n2602 & n2635;
  assign n4465 = n2642 & ~n4464;
  assign n4466 = ~n4463 & n4465;
  assign n4467 = ~n4462 & ~n4466;
  assign n4468 = n2682 & ~n4460;
  assign n4469 = ~n4467 & ~n4468;
  assign n4470 = ~n4461 & n4465;
  assign n4471 = n2678 & ~n2681;
  assign n4472 = n4460 & ~n4463;
  assign n4473 = ~n4471 & ~n4472;
  assign n4474 = ~n4470 & n4473;
  assign n4475 = n4469 & ~n4474;
  assign n5039 = x53 & x54;
  assign n5040 = x51 & x52;
  assign n5041 = ~n5039 & ~n5040;
  assign n5042 = ~x53 & ~x54;
  assign n5043 = ~x51 & ~x52;
  assign n5044 = ~n5042 & ~n5043;
  assign n5045 = ~n5041 & n5044;
  assign n5046 = x50 & n5045;
  assign n5047 = n5039 & n5040;
  assign n5048 = ~n5046 & ~n5047;
  assign n5049 = n5041 & ~n5044;
  assign n5050 = ~x50 & n5049;
  assign n5051 = n5048 & ~n5050;
  assign n5052 = ~x49 & ~n5051;
  assign n5053 = ~n5047 & ~n5049;
  assign n5054 = x50 & ~n5053;
  assign n5055 = ~x50 & ~n5045;
  assign n5056 = x49 & ~n5055;
  assign n5057 = ~n5054 & n5056;
  assign n4478 = x50 ^ x49;
  assign n5058 = n5042 & n5043;
  assign n5059 = n4478 & n5058;
  assign n5060 = ~n5057 & ~n5059;
  assign n5061 = ~n5052 & n5060;
  assign n5010 = x47 & x48;
  assign n5011 = x45 & x46;
  assign n5012 = ~n5010 & ~n5011;
  assign n5013 = ~x47 & ~x48;
  assign n5014 = ~x45 & ~x46;
  assign n5015 = ~n5013 & ~n5014;
  assign n5016 = ~n5012 & n5015;
  assign n5017 = x44 & n5016;
  assign n5018 = n5010 & n5011;
  assign n5019 = ~n5017 & ~n5018;
  assign n5020 = n5012 & ~n5015;
  assign n5021 = ~x44 & n5020;
  assign n5022 = n5013 & n5014;
  assign n5023 = ~n5021 & ~n5022;
  assign n5024 = n5019 & n5023;
  assign n5025 = ~x43 & ~n5024;
  assign n4483 = x44 ^ x43;
  assign n5026 = n4483 & n5016;
  assign n5027 = x43 & x44;
  assign n5028 = n5011 & n5027;
  assign n5029 = x48 & n5028;
  assign n5030 = n5029 ^ n5027;
  assign n5031 = ~n5020 & n5030;
  assign n5032 = ~n5026 & ~n5031;
  assign n5033 = ~x44 & ~x48;
  assign n5034 = n5014 & n5033;
  assign n5035 = ~n5028 & ~n5034;
  assign n5036 = ~x47 & ~n5035;
  assign n5037 = n5032 & ~n5036;
  assign n5038 = ~n5025 & n5037;
  assign n5062 = n5061 ^ n5038;
  assign n5102 = x39 & x40;
  assign n5103 = x41 & x42;
  assign n5104 = ~n5102 & ~n5103;
  assign n5105 = ~x39 & ~x40;
  assign n5106 = ~x41 & ~x42;
  assign n5107 = ~n5105 & ~n5106;
  assign n5108 = ~n5104 & n5107;
  assign n5109 = x38 & n5108;
  assign n5110 = n5102 & n5103;
  assign n5111 = ~n5109 & ~n5110;
  assign n5112 = x38 & ~n5106;
  assign n5113 = ~n5103 & n5105;
  assign n5114 = ~n5112 & n5113;
  assign n5115 = n5111 & ~n5114;
  assign n5116 = ~x37 & ~n5115;
  assign n4494 = x38 ^ x37;
  assign n4493 = x40 ^ x39;
  assign n4495 = n4494 ^ n4493;
  assign n5117 = ~x38 & ~x42;
  assign n5118 = ~n5102 & n5117;
  assign n5119 = n4495 & n5118;
  assign n5120 = x37 & x38;
  assign n5121 = n5102 & n5120;
  assign n5122 = ~n5119 & ~n5121;
  assign n5123 = ~x41 & ~n5122;
  assign n5124 = n5104 & ~n5107;
  assign n5125 = x42 & n5121;
  assign n5126 = n5125 ^ n5120;
  assign n5127 = ~n5124 & n5126;
  assign n5128 = n4494 & n5108;
  assign n5129 = ~n5127 & ~n5128;
  assign n5130 = ~n5123 & n5129;
  assign n5131 = ~n5116 & n5130;
  assign n5072 = x33 & x34;
  assign n5073 = x35 & x36;
  assign n5074 = ~n5072 & ~n5073;
  assign n5075 = ~x33 & ~x34;
  assign n5076 = ~x35 & ~x36;
  assign n5077 = ~n5075 & ~n5076;
  assign n5078 = ~n5074 & n5077;
  assign n5079 = x32 & n5078;
  assign n5080 = n5072 & n5073;
  assign n5081 = ~n5079 & ~n5080;
  assign n5082 = n5074 & ~n5077;
  assign n5083 = ~x32 & n5082;
  assign n5084 = n5075 & n5076;
  assign n5085 = ~n5083 & ~n5084;
  assign n5086 = n5081 & n5085;
  assign n5087 = ~x31 & ~n5086;
  assign n5088 = ~x32 & n5078;
  assign n5089 = x36 & n5072;
  assign n5090 = x32 & ~n5089;
  assign n5091 = ~n5082 & n5090;
  assign n5092 = ~n5088 & ~n5091;
  assign n5093 = x31 & ~n5092;
  assign n5094 = x31 & x32;
  assign n5095 = n5072 & n5094;
  assign n5096 = ~x32 & ~x36;
  assign n5097 = n5075 & n5096;
  assign n5098 = ~n5095 & ~n5097;
  assign n5099 = ~x35 & ~n5098;
  assign n5100 = ~n5093 & ~n5099;
  assign n5101 = ~n5087 & n5100;
  assign n5132 = n5131 ^ n5101;
  assign n4489 = x34 ^ x33;
  assign n4488 = x36 ^ x35;
  assign n4490 = n4489 ^ n4488;
  assign n4487 = x32 ^ x31;
  assign n4491 = n4490 ^ n4487;
  assign n4492 = x42 ^ x41;
  assign n4496 = n4495 ^ n4492;
  assign n5063 = n4491 & n4496;
  assign n4477 = x52 ^ x51;
  assign n4479 = n4478 ^ n4477;
  assign n4476 = x54 ^ x53;
  assign n4480 = n4479 ^ n4476;
  assign n4482 = x46 ^ x45;
  assign n4484 = n4483 ^ n4482;
  assign n4481 = x48 ^ x47;
  assign n4485 = n4484 ^ n4481;
  assign n5064 = ~n4480 & ~n4485;
  assign n5065 = ~n5063 & n5064;
  assign n5066 = n4480 & n4485;
  assign n5067 = ~n4491 & ~n4496;
  assign n5068 = ~n5066 & n5067;
  assign n5069 = ~n5065 & ~n5068;
  assign n5070 = n5063 & n5066;
  assign n5071 = n5069 & ~n5070;
  assign n5133 = n5132 ^ n5071;
  assign n6115 = n5133 ^ n5066;
  assign n6116 = ~n5062 & n6115;
  assign n6117 = n6116 ^ n5066;
  assign n6118 = n5069 ^ n5063;
  assign n6119 = ~n5132 & ~n6118;
  assign n6120 = n6119 ^ n5063;
  assign n6121 = ~n6117 & ~n6120;
  assign n6111 = n5062 & ~n5066;
  assign n6112 = ~n5038 & ~n5061;
  assign n6113 = ~n6111 & ~n6112;
  assign n6109 = n5048 & ~n5057;
  assign n6108 = n5019 & n5032;
  assign n6110 = n6109 ^ n6108;
  assign n6114 = n6113 ^ n6110;
  assign n6122 = n6121 ^ n6114;
  assign n6103 = ~n5063 & n5132;
  assign n6104 = ~n5101 & ~n5131;
  assign n6105 = ~n6103 & ~n6104;
  assign n6102 = n5081 & ~n5093;
  assign n6106 = n6105 ^ n6102;
  assign n6101 = n5111 & n5129;
  assign n6107 = n6106 ^ n6101;
  assign n6255 = n6114 ^ n6107;
  assign n6256 = n6122 & ~n6255;
  assign n6257 = n6256 ^ n6121;
  assign n6258 = n6113 ^ n6109;
  assign n6259 = ~n6110 & ~n6258;
  assign n6260 = n6259 ^ n6113;
  assign n6261 = n6102 ^ n6101;
  assign n6262 = ~n6106 & ~n6261;
  assign n6263 = n6262 ^ n6105;
  assign n6536 = n6260 & n6263;
  assign n6537 = n6257 & n6536;
  assign n4506 = x62 ^ x61;
  assign n4924 = x65 & x66;
  assign n4933 = ~x63 & ~x64;
  assign n4938 = n4924 & ~n4933;
  assign n4928 = x63 & x64;
  assign n4929 = ~x65 & ~x66;
  assign n4939 = n4928 & ~n4929;
  assign n4940 = ~n4938 & ~n4939;
  assign n4941 = n4506 & ~n4940;
  assign n4505 = x64 ^ x63;
  assign n4925 = n4924 ^ x64;
  assign n4926 = ~n4505 & ~n4925;
  assign n4930 = ~n4928 & n4929;
  assign n4942 = x61 & x62;
  assign n4943 = ~n4930 & n4942;
  assign n4944 = ~n4926 & n4943;
  assign n4945 = ~n4941 & ~n4944;
  assign n6127 = n4924 & n4928;
  assign n6128 = n4945 & ~n6127;
  assign n4927 = ~x61 & n4926;
  assign n4931 = ~x62 & n4930;
  assign n4932 = ~n4927 & ~n4931;
  assign n4934 = x61 & ~n4933;
  assign n4935 = x62 & ~n4929;
  assign n4936 = ~n4934 & ~n4935;
  assign n4937 = ~n4932 & n4936;
  assign n4946 = ~n4937 & n4945;
  assign n4899 = x57 & x58;
  assign n4900 = ~x59 & ~x60;
  assign n4901 = ~n4899 & n4900;
  assign n4902 = ~x56 & n4901;
  assign n4903 = x59 & x60;
  assign n4904 = ~x57 & ~x58;
  assign n4905 = ~n4903 & n4904;
  assign n4906 = x56 & ~n4900;
  assign n4907 = n4905 & ~n4906;
  assign n4908 = ~n4902 & ~n4907;
  assign n4909 = n4899 & n4903;
  assign n4910 = n4908 & ~n4909;
  assign n4911 = ~x55 & ~n4910;
  assign n4912 = ~n4901 & ~n4909;
  assign n4913 = x55 & x56;
  assign n4914 = ~n4905 & n4913;
  assign n4915 = n4912 & n4914;
  assign n4501 = x56 ^ x55;
  assign n4916 = n4903 & ~n4904;
  assign n4917 = n4899 & ~n4900;
  assign n4918 = ~n4916 & ~n4917;
  assign n4919 = n4501 & ~n4918;
  assign n4920 = ~n4915 & ~n4919;
  assign n4921 = n4902 & n4904;
  assign n4922 = n4920 & ~n4921;
  assign n4923 = ~n4911 & n4922;
  assign n4947 = n4946 ^ n4923;
  assign n4500 = x58 ^ x57;
  assign n4502 = n4501 ^ n4500;
  assign n4499 = x60 ^ x59;
  assign n4503 = n4502 ^ n4499;
  assign n4507 = n4506 ^ n4505;
  assign n4504 = x66 ^ x65;
  assign n4508 = n4507 ^ n4504;
  assign n4895 = n4503 & n4508;
  assign n6124 = n4923 ^ n4895;
  assign n6125 = n4947 & ~n6124;
  assign n6126 = n6125 ^ n4946;
  assign n6129 = ~n4909 & n4920;
  assign n4978 = x75 & x76;
  assign n4979 = x77 & x78;
  assign n4980 = ~n4978 & ~n4979;
  assign n4981 = ~x75 & ~x76;
  assign n4982 = ~x77 & ~x78;
  assign n4983 = ~n4981 & ~n4982;
  assign n4984 = ~n4980 & n4983;
  assign n4985 = x74 & n4984;
  assign n4986 = n4978 & n4979;
  assign n4987 = ~n4985 & ~n4986;
  assign n4988 = n4980 & ~n4983;
  assign n4989 = ~x74 & n4988;
  assign n4990 = n4981 & n4982;
  assign n4991 = ~n4989 & ~n4990;
  assign n4992 = n4987 & n4991;
  assign n4993 = ~x73 & ~n4992;
  assign n4517 = x74 ^ x73;
  assign n4994 = n4517 & n4984;
  assign n4995 = x73 & x74;
  assign n4996 = n4978 & n4995;
  assign n4997 = x78 & n4996;
  assign n4998 = n4997 ^ n4995;
  assign n4999 = ~n4988 & n4998;
  assign n5000 = ~n4994 & ~n4999;
  assign n5001 = ~x74 & ~x78;
  assign n5002 = n4981 & n5001;
  assign n5003 = ~n4996 & ~n5002;
  assign n5004 = ~x77 & ~n5003;
  assign n5005 = n5000 & ~n5004;
  assign n5006 = ~n4993 & n5005;
  assign n4949 = x69 & x70;
  assign n4950 = x71 & x72;
  assign n4951 = ~n4949 & ~n4950;
  assign n4952 = ~x69 & ~x70;
  assign n4953 = ~x71 & ~x72;
  assign n4954 = ~n4952 & ~n4953;
  assign n4955 = ~n4951 & n4954;
  assign n4956 = x68 & n4955;
  assign n4957 = n4949 & n4950;
  assign n4958 = ~n4956 & ~n4957;
  assign n4959 = n4951 & ~n4954;
  assign n4960 = ~x68 & n4959;
  assign n4961 = n4952 & n4953;
  assign n4962 = ~n4960 & ~n4961;
  assign n4963 = n4958 & n4962;
  assign n4964 = ~x67 & ~n4963;
  assign n4512 = x68 ^ x67;
  assign n4965 = n4512 & n4955;
  assign n4966 = x67 & x68;
  assign n4967 = n4949 & n4966;
  assign n4968 = x72 & n4967;
  assign n4969 = n4968 ^ n4966;
  assign n4970 = ~n4959 & n4969;
  assign n4971 = ~n4965 & ~n4970;
  assign n4972 = ~x68 & ~x72;
  assign n4973 = n4952 & n4972;
  assign n4974 = ~n4967 & ~n4973;
  assign n4975 = ~x71 & ~n4974;
  assign n4976 = n4971 & ~n4975;
  assign n4977 = ~n4964 & n4976;
  assign n5007 = n5006 ^ n4977;
  assign n4509 = n4508 ^ n4503;
  assign n4516 = x76 ^ x75;
  assign n4518 = n4517 ^ n4516;
  assign n4515 = x78 ^ x77;
  assign n4519 = n4518 ^ n4515;
  assign n4511 = x70 ^ x69;
  assign n4513 = n4512 ^ n4511;
  assign n4510 = x72 ^ x71;
  assign n4514 = n4513 ^ n4510;
  assign n4520 = n4519 ^ n4514;
  assign n4894 = n4509 & n4520;
  assign n4896 = n4514 & n4519;
  assign n4897 = n4896 ^ n4895;
  assign n4898 = ~n4894 & ~n4897;
  assign n4948 = n4947 ^ n4898;
  assign n5008 = n5007 ^ n4948;
  assign n6140 = ~n4896 & ~n5007;
  assign n6141 = n5008 & ~n6140;
  assign n6142 = ~n4947 & ~n6141;
  assign n6143 = n4895 & n4947;
  assign n6144 = n4948 ^ n4896;
  assign n6145 = ~n5007 & ~n6144;
  assign n6146 = n6145 ^ n4896;
  assign n6147 = ~n6143 & ~n6146;
  assign n6148 = ~n6142 & n6147;
  assign n6270 = n6129 & ~n6148;
  assign n6271 = ~n6126 & n6270;
  assign n6272 = ~n6128 & ~n6271;
  assign n6135 = n4896 & n5007;
  assign n6136 = n4977 & n5006;
  assign n6137 = ~n6135 & ~n6136;
  assign n6133 = n4987 & n5000;
  assign n6132 = n4958 & n4971;
  assign n6134 = n6133 ^ n6132;
  assign n6138 = n6137 ^ n6134;
  assign n6130 = n6129 ^ n6128;
  assign n6131 = n6130 ^ n6126;
  assign n6139 = n6138 ^ n6131;
  assign n6149 = n6148 ^ n6139;
  assign n6273 = ~n6138 & n6149;
  assign n6274 = ~n6272 & ~n6273;
  assign n6275 = n6129 ^ n6126;
  assign n6276 = n6148 ^ n6129;
  assign n6277 = n6275 & ~n6276;
  assign n6278 = n6277 ^ n6148;
  assign n6279 = n6274 & ~n6278;
  assign n6280 = n6273 & n6278;
  assign n6281 = ~n6279 & ~n6280;
  assign n6267 = n6137 ^ n6133;
  assign n6268 = ~n6134 & n6267;
  assign n6269 = n6268 ^ n6137;
  assign n6282 = n6281 ^ n6269;
  assign n6532 = n6269 & ~n6280;
  assign n6533 = ~n6279 & ~n6532;
  assign n6534 = ~n6260 & ~n6263;
  assign n6535 = ~n6257 & n6534;
  assign n6538 = ~n6535 & ~n6537;
  assign n6539 = n6533 & n6538;
  assign n6540 = ~n6282 & ~n6539;
  assign n6123 = n6122 ^ n6107;
  assign n6150 = n6149 ^ n6123;
  assign n5134 = n5133 ^ n5062;
  assign n6097 = n5134 ^ n5008;
  assign n4497 = n4496 ^ n4491;
  assign n4486 = n4485 ^ n4480;
  assign n4498 = n4497 ^ n4486;
  assign n4521 = n4520 ^ n4509;
  assign n4893 = n4498 & n4521;
  assign n6098 = n5134 ^ n4893;
  assign n6099 = ~n6097 & ~n6098;
  assign n6100 = n6099 ^ n5008;
  assign n6252 = n6123 ^ n6100;
  assign n6253 = ~n6150 & n6252;
  assign n6254 = n6253 ^ n6149;
  assign n6264 = n6263 ^ n6260;
  assign n6541 = n6263 ^ n6257;
  assign n6542 = ~n6264 & n6541;
  assign n6543 = n6542 ^ n6257;
  assign n6544 = ~n6254 & n6543;
  assign n6545 = n6540 & ~n6544;
  assign n6571 = ~n6537 & n6545;
  assign n6548 = ~n6254 & ~n6535;
  assign n6549 = ~n6543 & ~n6548;
  assign n6572 = ~n6279 & ~n6549;
  assign n6573 = n6282 & ~n6572;
  assign n6574 = ~n6571 & ~n6573;
  assign n4528 = x5 ^ x4;
  assign n4529 = n4528 ^ x3;
  assign n4530 = x2 ^ x1;
  assign n4531 = n4530 ^ x0;
  assign n5170 = n4529 & n4531;
  assign n5180 = x1 ^ x0;
  assign n5181 = ~n4530 & n5180;
  assign n5182 = n5181 ^ x0;
  assign n5177 = x4 ^ x3;
  assign n5178 = ~n4528 & n5177;
  assign n5179 = n5178 ^ x3;
  assign n5183 = n5182 ^ n5179;
  assign n6157 = n5170 & n5183;
  assign n6158 = n5179 & n5182;
  assign n6159 = ~n6157 & ~n6158;
  assign n5136 = x995 & x996;
  assign n5137 = x993 & x994;
  assign n5138 = ~n5136 & ~n5137;
  assign n5139 = ~x995 & ~x996;
  assign n5140 = ~x993 & ~x994;
  assign n5141 = ~n5139 & ~n5140;
  assign n5142 = ~n5138 & n5141;
  assign n5143 = x992 & n5142;
  assign n5144 = n5136 & n5137;
  assign n5145 = ~n5143 & ~n5144;
  assign n4525 = x992 ^ x991;
  assign n5152 = n4525 & n5142;
  assign n5146 = n5138 & ~n5141;
  assign n5153 = x991 & x992;
  assign n5154 = n5137 & n5153;
  assign n5155 = x996 & n5154;
  assign n5156 = n5155 ^ n5153;
  assign n5157 = ~n5146 & n5156;
  assign n5158 = ~n5152 & ~n5157;
  assign n6156 = n5145 & n5158;
  assign n6160 = n6159 ^ n6156;
  assign n4533 = x999 ^ x998;
  assign n5174 = x998 ^ x997;
  assign n5175 = ~n4533 & n5174;
  assign n5176 = n5175 ^ x997;
  assign n5184 = n5183 ^ n5176;
  assign n4534 = n4533 ^ x997;
  assign n5166 = x6 & n4534;
  assign n4532 = n4531 ^ n4529;
  assign n4535 = n4534 ^ x6;
  assign n5167 = n4535 ^ n4531;
  assign n5168 = ~n4532 & n5167;
  assign n5169 = n5168 ^ n4535;
  assign n5171 = n5170 ^ n5169;
  assign n5172 = ~n5166 & ~n5171;
  assign n5173 = n5172 ^ n5170;
  assign n5185 = n5184 ^ n5173;
  assign n6164 = ~n5176 & ~n5185;
  assign n6165 = ~n5171 & ~n5183;
  assign n6166 = n6165 ^ n5170;
  assign n6167 = ~n5166 & n6166;
  assign n6168 = ~n6164 & ~n6167;
  assign n4524 = x994 ^ x993;
  assign n4526 = n4525 ^ n4524;
  assign n4523 = x996 ^ x995;
  assign n4527 = n4526 ^ n4523;
  assign n4536 = n4535 ^ n4532;
  assign n5165 = n4527 & n4536;
  assign n5186 = n5185 ^ n5165;
  assign n5147 = ~x992 & n5146;
  assign n5148 = n5139 & n5140;
  assign n5149 = ~n5147 & ~n5148;
  assign n5150 = n5145 & n5149;
  assign n5151 = ~x991 & ~n5150;
  assign n5159 = ~x992 & ~x996;
  assign n5160 = n5140 & n5159;
  assign n5161 = ~n5154 & ~n5160;
  assign n5162 = ~x995 & ~n5161;
  assign n5163 = n5158 & ~n5162;
  assign n5164 = ~n5151 & n5163;
  assign n6161 = n5165 ^ n5164;
  assign n6162 = ~n5186 & ~n6161;
  assign n6163 = n6162 ^ n5185;
  assign n6169 = n6168 ^ n6163;
  assign n6244 = n6160 & ~n6169;
  assign n6241 = ~n6163 & n6168;
  assign n6242 = ~n6156 & ~n6159;
  assign n6245 = ~n6241 & ~n6242;
  assign n6246 = ~n6244 & n6245;
  assign n4545 = x10 ^ x9;
  assign n4544 = x8 ^ x7;
  assign n4546 = n4545 ^ n4544;
  assign n4543 = x12 ^ x11;
  assign n4547 = n4546 ^ n4543;
  assign n4540 = x16 ^ x15;
  assign n4539 = x18 ^ x17;
  assign n4541 = n4540 ^ n4539;
  assign n4538 = x14 ^ x13;
  assign n4542 = n4541 ^ n4538;
  assign n4548 = n4547 ^ n4542;
  assign n4556 = x28 ^ x27;
  assign n4555 = x30 ^ x29;
  assign n4557 = n4556 ^ n4555;
  assign n4554 = x26 ^ x25;
  assign n4558 = n4557 ^ n4554;
  assign n4551 = x22 ^ x21;
  assign n4550 = x20 ^ x19;
  assign n4552 = n4551 ^ n4550;
  assign n4549 = x24 ^ x23;
  assign n4553 = n4552 ^ n4549;
  assign n4559 = n4558 ^ n4553;
  assign n5188 = n4559 ^ n4547;
  assign n5189 = ~n4548 & n5188;
  assign n5190 = n5189 ^ n4559;
  assign n5299 = x23 & x24;
  assign n5300 = x21 & x22;
  assign n5301 = ~n5299 & ~n5300;
  assign n5302 = ~x23 & ~x24;
  assign n5303 = ~x21 & ~x22;
  assign n5304 = ~n5302 & ~n5303;
  assign n5305 = ~n5301 & n5304;
  assign n5306 = x20 & n5305;
  assign n5307 = n5299 & n5300;
  assign n5308 = ~n5306 & ~n5307;
  assign n5309 = n5301 & ~n5304;
  assign n5310 = ~x20 & n5309;
  assign n5311 = n5302 & n5303;
  assign n5312 = ~n5310 & ~n5311;
  assign n5313 = n5308 & n5312;
  assign n5314 = ~x19 & ~n5313;
  assign n5315 = ~x20 & ~n5305;
  assign n5316 = x19 & ~n5309;
  assign n5317 = ~n5315 & n5316;
  assign n5318 = x20 & x24;
  assign n5319 = n5300 & n5318;
  assign n5320 = n5317 & ~n5319;
  assign n5321 = x21 ^ x20;
  assign n5322 = x24 ^ x22;
  assign n5323 = ~n4551 & ~n5322;
  assign n5324 = ~n5321 & n5323;
  assign n5325 = ~x23 & n5324;
  assign n5326 = ~n5320 & ~n5325;
  assign n5327 = ~n5314 & n5326;
  assign n5264 = ~x29 & ~x30;
  assign n5265 = x25 & ~n5264;
  assign n5266 = x29 & x30;
  assign n5267 = n5266 ^ x28;
  assign n5268 = n4556 & ~n5267;
  assign n5269 = n5268 ^ x27;
  assign n5270 = n5265 & n5269;
  assign n5271 = x25 & x26;
  assign n5272 = ~n5270 & ~n5271;
  assign n5273 = ~x27 & ~x28;
  assign n5274 = ~n5266 & n5273;
  assign n5275 = x27 & x28;
  assign n5276 = ~n5264 & ~n5275;
  assign n5277 = ~n5274 & n5276;
  assign n5278 = ~x30 & n5275;
  assign n5279 = x26 & ~n5278;
  assign n5280 = ~n5277 & n5279;
  assign n5281 = ~n5272 & ~n5280;
  assign n5282 = n5266 & n5275;
  assign n5283 = x26 & ~n5264;
  assign n5284 = ~n5282 & ~n5283;
  assign n5285 = n5269 & ~n5284;
  assign n5286 = ~x26 & ~n5275;
  assign n5287 = n5264 & n5286;
  assign n5288 = n5274 & ~n5283;
  assign n5289 = ~n5287 & ~n5288;
  assign n5290 = ~n5285 & n5289;
  assign n5291 = ~x25 & ~n5290;
  assign n5292 = ~n5281 & ~n5291;
  assign n5293 = n5271 & n5275;
  assign n5294 = ~x26 & ~x30;
  assign n5295 = n5273 & n5294;
  assign n5296 = ~n5293 & ~n5295;
  assign n5297 = ~x29 & ~n5296;
  assign n5298 = n5292 & ~n5297;
  assign n5328 = n5327 ^ n5298;
  assign n5263 = n4553 & n4558;
  assign n5329 = n5328 ^ n5263;
  assign n6187 = ~n5190 & ~n5329;
  assign n5227 = ~x17 & ~x18;
  assign n5228 = x13 & ~n5227;
  assign n5229 = x17 & x18;
  assign n5230 = n5229 ^ x16;
  assign n5231 = n4540 & ~n5230;
  assign n5232 = n5231 ^ x15;
  assign n5233 = n5228 & n5232;
  assign n5234 = x13 & x14;
  assign n5235 = ~n5233 & ~n5234;
  assign n5236 = ~x15 & ~x16;
  assign n5237 = ~n5229 & n5236;
  assign n5238 = x15 & x16;
  assign n5239 = ~n5227 & ~n5238;
  assign n5240 = ~n5237 & n5239;
  assign n5241 = ~x18 & n5238;
  assign n5242 = x14 & ~n5241;
  assign n5243 = ~n5240 & n5242;
  assign n5244 = ~n5235 & ~n5243;
  assign n5245 = n5229 & n5238;
  assign n5246 = x14 & ~n5227;
  assign n5247 = ~n5245 & ~n5246;
  assign n5248 = n5232 & ~n5247;
  assign n5249 = ~x14 & ~n5238;
  assign n5250 = n5227 & n5249;
  assign n5251 = n5237 & ~n5246;
  assign n5252 = ~n5250 & ~n5251;
  assign n5253 = ~n5248 & n5252;
  assign n5254 = ~x13 & ~n5253;
  assign n5255 = ~n5244 & ~n5254;
  assign n5256 = n5234 & n5238;
  assign n5257 = ~x14 & ~x18;
  assign n5258 = n5236 & n5257;
  assign n5259 = ~n5256 & ~n5258;
  assign n5260 = ~x17 & ~n5259;
  assign n5261 = n5255 & ~n5260;
  assign n5193 = ~x11 & ~x12;
  assign n5194 = x8 & ~n5193;
  assign n5195 = ~x9 & ~x10;
  assign n5196 = x11 & x12;
  assign n5197 = n5195 & ~n5196;
  assign n5198 = ~n5194 & n5197;
  assign n5200 = n5194 & ~n5195;
  assign n5199 = x9 & x10;
  assign n5201 = n5200 ^ n5199;
  assign n5202 = n5199 ^ n5196;
  assign n5203 = n5201 & ~n5202;
  assign n5204 = n5203 ^ n5200;
  assign n5205 = ~n5198 & ~n5204;
  assign n5206 = ~x7 & ~n5205;
  assign n5207 = ~n5196 & ~n5199;
  assign n5208 = ~n5193 & ~n5195;
  assign n5209 = ~x8 & ~n5208;
  assign n5210 = x8 & x9;
  assign n5211 = x12 & n5210;
  assign n5212 = x7 & ~n5211;
  assign n5213 = ~n5209 & n5212;
  assign n5214 = ~n5207 & n5213;
  assign n5215 = x7 & n4545;
  assign n5216 = n5194 & n5215;
  assign n5217 = ~n5214 & ~n5216;
  assign n5218 = ~x11 & ~n5215;
  assign n5220 = x7 & x8;
  assign n5219 = ~x8 & ~x12;
  assign n5221 = n5220 ^ n5219;
  assign n5222 = ~n5199 & n5221;
  assign n5223 = n5222 ^ n5220;
  assign n5224 = n5218 & n5223;
  assign n5225 = n5217 & ~n5224;
  assign n5226 = ~n5206 & n5225;
  assign n5262 = n5261 ^ n5226;
  assign n6178 = n4542 & n4547;
  assign n6188 = n5262 & ~n6178;
  assign n6189 = ~n6187 & n6188;
  assign n6190 = n5190 & ~n5262;
  assign n6191 = n5329 & n6190;
  assign n6192 = ~n6189 & ~n6191;
  assign n6183 = ~n5204 & n5217;
  assign n6182 = ~n5244 & ~n5248;
  assign n6184 = n6183 ^ n6182;
  assign n6179 = n6178 ^ n5261;
  assign n6180 = ~n5262 & n6179;
  assign n6181 = n6180 ^ n6178;
  assign n6185 = n6184 ^ n6181;
  assign n6175 = ~n5281 & ~n5285;
  assign n6174 = n5308 & ~n5317;
  assign n6176 = n6175 ^ n6174;
  assign n6171 = n5298 ^ n5263;
  assign n6172 = n5328 & ~n6171;
  assign n6173 = n6172 ^ n5327;
  assign n6177 = n6176 ^ n6173;
  assign n6186 = n6185 ^ n6177;
  assign n6193 = n6192 ^ n6186;
  assign n6170 = n6169 ^ n6160;
  assign n6194 = n6193 ^ n6170;
  assign n5330 = n5329 ^ n5262;
  assign n4537 = n4536 ^ n4527;
  assign n4560 = n4559 ^ n4548;
  assign n5191 = n4537 & n4560;
  assign n5192 = n5191 ^ n5190;
  assign n5331 = n5330 ^ n5192;
  assign n5187 = n5186 ^ n5164;
  assign n6153 = n5191 ^ n5187;
  assign n6154 = n5331 & ~n6153;
  assign n6155 = n6154 ^ n5191;
  assign n6228 = n6170 ^ n6155;
  assign n6229 = n6194 & n6228;
  assign n6230 = n6229 ^ n6193;
  assign n6243 = n6241 & n6242;
  assign n6512 = n6230 & ~n6243;
  assign n6237 = n6175 ^ n6173;
  assign n6238 = ~n6176 & ~n6237;
  assign n6239 = n6238 ^ n6173;
  assign n6234 = n6183 ^ n6181;
  assign n6235 = ~n6184 & ~n6234;
  assign n6236 = n6235 ^ n6181;
  assign n6240 = n6239 ^ n6236;
  assign n6231 = n6192 ^ n6185;
  assign n6232 = ~n6186 & ~n6231;
  assign n6233 = n6232 ^ n6192;
  assign n6520 = n6236 ^ n6233;
  assign n6521 = n6240 & n6520;
  assign n6522 = n6521 ^ n6239;
  assign n6523 = ~n6512 & n6522;
  assign n6524 = n6236 & n6239;
  assign n6525 = ~n6233 & n6524;
  assign n6526 = ~n6523 & ~n6525;
  assign n6527 = ~n6246 & ~n6526;
  assign n6575 = n6574 ^ n6527;
  assign n6513 = ~n6239 & n6246;
  assign n6514 = ~n6512 & ~n6513;
  assign n6247 = ~n6243 & ~n6246;
  assign n6248 = n6247 ^ n6240;
  assign n6249 = n6248 ^ n6233;
  assign n6250 = n6249 ^ n6230;
  assign n6515 = ~n6236 & n6250;
  assign n6516 = ~n6514 & n6515;
  assign n6517 = n6230 & n6513;
  assign n6518 = ~n6516 & ~n6517;
  assign n6519 = n6233 & ~n6518;
  assign n6528 = ~n6236 & n6517;
  assign n6529 = ~n6527 & ~n6528;
  assign n6530 = ~n6519 & n6529;
  assign n6265 = n6264 ^ n6257;
  assign n6266 = n6265 ^ n6254;
  assign n6283 = n6282 ^ n6266;
  assign n6508 = n6283 ^ n6250;
  assign n6151 = n6150 ^ n6100;
  assign n4522 = n4521 ^ n4498;
  assign n4561 = n4560 ^ n4537;
  assign n6035 = n4522 & n4561;
  assign n5332 = n5331 ^ n5187;
  assign n6093 = n6035 ^ n5332;
  assign n5009 = n5008 ^ n4893;
  assign n5135 = n5134 ^ n5009;
  assign n6094 = n6035 ^ n5135;
  assign n6095 = ~n6093 & n6094;
  assign n6096 = n6095 ^ n5332;
  assign n6152 = n6151 ^ n6096;
  assign n6195 = n6194 ^ n6155;
  assign n6225 = n6195 ^ n6096;
  assign n6226 = ~n6152 & n6225;
  assign n6227 = n6226 ^ n6151;
  assign n6509 = n6283 ^ n6227;
  assign n6510 = n6508 & ~n6509;
  assign n6511 = n6510 ^ n6250;
  assign n6531 = n6530 ^ n6511;
  assign n6546 = ~n6533 & n6537;
  assign n6547 = n6545 & ~n6546;
  assign n6550 = n6549 ^ n6279;
  assign n6551 = n6282 & n6550;
  assign n6552 = ~n6547 & ~n6551;
  assign n6553 = n6254 & n6535;
  assign n6554 = ~n6533 & n6553;
  assign n6555 = ~n6552 & ~n6554;
  assign n6568 = n6555 ^ n6530;
  assign n6569 = ~n6531 & n6568;
  assign n6570 = n6569 ^ n6555;
  assign n6576 = n6575 ^ n6570;
  assign n6614 = ~n6527 & ~n6574;
  assign n6615 = ~n6576 & ~n6614;
  assign n4783 = ~x989 & ~x990;
  assign n4784 = x985 & ~n4783;
  assign n4598 = x988 ^ x987;
  assign n4785 = x989 & x990;
  assign n4786 = n4785 ^ x988;
  assign n4787 = n4598 & ~n4786;
  assign n4788 = n4787 ^ x987;
  assign n4789 = n4784 & n4788;
  assign n4790 = x985 & x986;
  assign n4791 = ~n4789 & ~n4790;
  assign n4792 = ~x987 & ~x988;
  assign n4793 = ~n4785 & n4792;
  assign n4794 = x987 & x988;
  assign n4795 = ~n4783 & ~n4794;
  assign n4796 = ~n4793 & n4795;
  assign n4797 = ~x990 & n4794;
  assign n4798 = x986 & ~n4797;
  assign n4799 = ~n4796 & n4798;
  assign n4800 = ~n4791 & ~n4799;
  assign n4801 = n4785 & n4794;
  assign n4802 = x986 & ~n4783;
  assign n4803 = ~n4801 & ~n4802;
  assign n4804 = n4788 & ~n4803;
  assign n6086 = ~n4800 & ~n4804;
  assign n4755 = ~x983 & ~x984;
  assign n4603 = x982 ^ x981;
  assign n4756 = x983 & x984;
  assign n4757 = n4756 ^ x982;
  assign n4758 = n4603 & ~n4757;
  assign n4759 = n4758 ^ x981;
  assign n4760 = ~n4755 & n4759;
  assign n4761 = ~x980 & ~n4760;
  assign n4762 = ~x981 & ~x982;
  assign n4763 = ~n4756 & n4762;
  assign n4764 = x979 & ~n4763;
  assign n4765 = x981 & x982;
  assign n4766 = n4755 & ~n4765;
  assign n4767 = n4756 & n4765;
  assign n4768 = ~n4766 & ~n4767;
  assign n4769 = n4764 & n4768;
  assign n4770 = x979 & ~x980;
  assign n4771 = ~n4769 & ~n4770;
  assign n4772 = ~n4761 & ~n4771;
  assign n4773 = x980 & ~n4755;
  assign n4774 = ~n4767 & ~n4773;
  assign n4775 = n4759 & ~n4774;
  assign n6085 = ~n4772 & ~n4775;
  assign n6087 = n6086 ^ n6085;
  assign n4805 = n4793 & ~n4802;
  assign n4806 = ~n4804 & ~n4805;
  assign n4807 = ~x985 & ~n4806;
  assign n4808 = ~n4800 & ~n4807;
  assign n4599 = x986 ^ x985;
  assign n4600 = n4599 ^ n4598;
  assign n4809 = ~x986 & ~x990;
  assign n4810 = ~n4794 & n4809;
  assign n4811 = n4600 & n4810;
  assign n4812 = n4790 & n4794;
  assign n4813 = ~n4811 & ~n4812;
  assign n4814 = ~x989 & ~n4813;
  assign n4815 = n4808 & ~n4814;
  assign n4776 = n4763 & ~n4773;
  assign n4777 = ~n4775 & ~n4776;
  assign n4778 = ~x979 & ~n4777;
  assign n4779 = ~n4772 & ~n4778;
  assign n4604 = x984 ^ x983;
  assign n4605 = n4604 ^ n4603;
  assign n4602 = x980 ^ x979;
  assign n4606 = n4605 ^ n4602;
  assign n4780 = ~x980 & n4766;
  assign n4781 = n4606 & n4780;
  assign n4782 = n4779 & ~n4781;
  assign n4816 = n4815 ^ n4782;
  assign n4597 = x990 ^ x989;
  assign n4601 = n4600 ^ n4597;
  assign n4817 = n4601 & n4606;
  assign n6082 = n4817 ^ n4815;
  assign n6083 = ~n4816 & n6082;
  assign n6084 = n6083 ^ n4817;
  assign n6088 = n6087 ^ n6084;
  assign n4593 = x974 ^ x973;
  assign n4591 = x976 ^ x975;
  assign n4854 = x977 & x978;
  assign n4855 = n4854 ^ x976;
  assign n4856 = n4591 & ~n4855;
  assign n4857 = n4856 ^ x975;
  assign n4858 = n4593 & n4857;
  assign n4859 = ~x975 & ~x976;
  assign n4860 = ~n4854 & n4859;
  assign n4861 = x975 & x976;
  assign n4862 = x973 & x974;
  assign n4863 = ~n4861 & n4862;
  assign n4864 = ~n4860 & n4863;
  assign n4865 = ~n4858 & ~n4864;
  assign n4866 = ~x977 & ~x978;
  assign n4867 = ~n4865 & ~n4866;
  assign n4868 = n4861 & n4862;
  assign n4869 = ~x978 & n4868;
  assign n4870 = ~n4867 & ~n4869;
  assign n4871 = n4854 & n4861;
  assign n4872 = x974 & ~n4866;
  assign n4873 = ~n4871 & ~n4872;
  assign n4874 = n4857 & ~n4873;
  assign n6079 = n4870 & ~n4874;
  assign n4826 = ~x969 & ~x970;
  assign n4827 = ~x971 & ~x972;
  assign n4828 = ~n4826 & ~n4827;
  assign n4829 = x969 & x970;
  assign n4830 = x971 & x972;
  assign n4831 = ~n4829 & ~n4830;
  assign n4832 = n4828 & ~n4831;
  assign n4833 = x968 & n4832;
  assign n4834 = n4829 & n4830;
  assign n4835 = ~n4833 & ~n4834;
  assign n4586 = x968 ^ x967;
  assign n4841 = n4586 & n4832;
  assign n4836 = ~n4828 & n4831;
  assign n4842 = x967 & x968;
  assign n4843 = n4829 & n4842;
  assign n4844 = x972 & n4843;
  assign n4845 = n4844 ^ n4842;
  assign n4846 = ~n4836 & n4845;
  assign n4847 = ~n4841 & ~n4846;
  assign n6078 = n4835 & n4847;
  assign n6080 = n6079 ^ n6078;
  assign n4875 = n4860 & ~n4872;
  assign n4876 = ~x974 & ~n4861;
  assign n4877 = n4866 & n4876;
  assign n4878 = ~n4875 & ~n4877;
  assign n4879 = ~n4874 & n4878;
  assign n4880 = ~x973 & ~n4879;
  assign n4881 = ~x974 & ~x978;
  assign n4882 = n4859 & n4881;
  assign n4883 = ~n4868 & ~n4882;
  assign n4884 = ~x977 & ~n4883;
  assign n4885 = ~n4880 & ~n4884;
  assign n4886 = n4870 & n4885;
  assign n4588 = x970 ^ x969;
  assign n4587 = x972 ^ x971;
  assign n4589 = n4588 ^ n4587;
  assign n4837 = x968 & n4589;
  assign n4838 = n4836 & ~n4837;
  assign n4839 = n4835 & ~n4838;
  assign n4840 = ~x967 & ~n4839;
  assign n4848 = ~x968 & ~x972;
  assign n4849 = n4826 & n4848;
  assign n4850 = ~n4843 & ~n4849;
  assign n4851 = ~x971 & ~n4850;
  assign n4852 = n4847 & ~n4851;
  assign n4853 = ~n4840 & n4852;
  assign n4887 = n4886 ^ n4853;
  assign n4590 = n4589 ^ n4586;
  assign n4592 = x978 ^ x977;
  assign n4594 = n4593 ^ n4592;
  assign n4595 = n4594 ^ n4591;
  assign n4820 = n4590 & n4595;
  assign n6075 = n4853 ^ n4820;
  assign n6076 = n4887 & ~n6075;
  assign n6077 = n6076 ^ n4886;
  assign n6081 = n6080 ^ n6077;
  assign n6089 = n6088 ^ n6081;
  assign n6068 = n4820 & n4887;
  assign n4818 = ~n4590 & ~n4595;
  assign n4819 = ~n4817 & n4818;
  assign n4821 = ~n4601 & ~n4606;
  assign n4822 = ~n4820 & n4821;
  assign n4823 = ~n4819 & ~n4822;
  assign n4824 = n4817 & n4820;
  assign n4825 = n4823 & ~n4824;
  assign n4888 = n4887 ^ n4825;
  assign n6069 = ~n4816 & n4888;
  assign n6070 = n4816 & n4817;
  assign n6071 = ~n4823 & ~n4887;
  assign n6072 = ~n6070 & ~n6071;
  assign n6073 = ~n6069 & n6072;
  assign n6074 = ~n6068 & n6073;
  assign n6090 = n6089 ^ n6074;
  assign n6311 = n6079 ^ n6077;
  assign n6312 = ~n6080 & ~n6311;
  assign n6313 = n6312 ^ n6077;
  assign n6314 = n6088 & n6313;
  assign n6315 = ~n6090 & n6314;
  assign n6316 = ~n6074 & ~n6088;
  assign n6317 = ~n6313 & n6316;
  assign n6318 = ~n6315 & ~n6317;
  assign n6319 = n6078 & n6079;
  assign n6320 = ~n6077 & n6319;
  assign n6321 = n6090 & n6320;
  assign n6322 = n6318 & ~n6321;
  assign n6308 = n6086 ^ n6084;
  assign n6309 = ~n6087 & ~n6308;
  assign n6310 = n6309 ^ n6084;
  assign n6323 = n6322 ^ n6310;
  assign n6501 = ~n6078 & ~n6079;
  assign n6502 = n6323 & ~n6501;
  assign n6503 = ~n6310 & ~n6315;
  assign n6504 = ~n6502 & ~n6503;
  assign n4643 = x951 & x952;
  assign n4644 = x953 & x954;
  assign n4645 = ~n4643 & ~n4644;
  assign n4646 = ~x951 & ~x952;
  assign n4647 = ~x953 & ~x954;
  assign n4648 = ~n4646 & ~n4647;
  assign n4649 = ~n4645 & n4648;
  assign n4650 = x950 & n4649;
  assign n4651 = n4643 & n4644;
  assign n4652 = ~n4650 & ~n4651;
  assign n4658 = n4645 & ~n4648;
  assign n4659 = x949 & x950;
  assign n4660 = n4643 & n4659;
  assign n4661 = x954 & n4660;
  assign n4662 = n4661 ^ n4659;
  assign n4663 = ~n4658 & n4662;
  assign n4576 = x950 ^ x949;
  assign n4664 = n4576 & n4649;
  assign n4665 = ~n4663 & ~n4664;
  assign n6047 = n4652 & n4665;
  assign n4613 = x945 & x946;
  assign n4614 = x947 & x948;
  assign n4615 = ~n4613 & ~n4614;
  assign n4616 = ~x945 & ~x946;
  assign n4617 = ~x947 & ~x948;
  assign n4618 = ~n4616 & ~n4617;
  assign n4619 = ~n4615 & n4618;
  assign n4620 = x944 & n4619;
  assign n4621 = n4613 & n4614;
  assign n4622 = ~n4620 & ~n4621;
  assign n4628 = n4615 & ~n4618;
  assign n4629 = x943 & x944;
  assign n4630 = n4613 & n4629;
  assign n4631 = x948 & n4630;
  assign n4632 = n4631 ^ n4629;
  assign n4633 = ~n4628 & n4632;
  assign n4581 = x944 ^ x943;
  assign n4634 = n4581 & n4619;
  assign n4635 = ~n4633 & ~n4634;
  assign n6048 = n4622 & n4635;
  assign n6299 = ~n6047 & ~n6048;
  assign n6289 = n6047 & n6048;
  assign n4717 = ~x959 & ~x960;
  assign n4718 = x956 & ~n4717;
  assign n4719 = x959 & x960;
  assign n4720 = x957 & x958;
  assign n4721 = n4719 & n4720;
  assign n4722 = ~n4718 & ~n4721;
  assign n4564 = x958 ^ x957;
  assign n4723 = n4719 ^ x958;
  assign n4724 = n4564 & ~n4723;
  assign n4725 = n4724 ^ x957;
  assign n4726 = ~n4722 & n4725;
  assign n4732 = x955 & ~n4717;
  assign n4733 = n4725 & n4732;
  assign n4734 = x955 & x956;
  assign n4735 = ~n4733 & ~n4734;
  assign n4727 = ~x957 & ~x958;
  assign n4728 = ~n4719 & n4727;
  assign n4736 = ~n4717 & ~n4720;
  assign n4737 = ~n4728 & n4736;
  assign n4738 = ~x960 & n4720;
  assign n4739 = x956 & ~n4738;
  assign n4740 = ~n4737 & n4739;
  assign n4741 = ~n4735 & ~n4740;
  assign n6055 = ~n4726 & ~n4741;
  assign n4683 = ~x965 & ~x966;
  assign n4684 = x962 & ~n4683;
  assign n4685 = x965 & x966;
  assign n4686 = x963 & x964;
  assign n4687 = n4685 & n4686;
  assign n4688 = ~n4684 & ~n4687;
  assign n4569 = x964 ^ x963;
  assign n4689 = n4685 ^ x964;
  assign n4690 = n4569 & ~n4689;
  assign n4691 = n4690 ^ x963;
  assign n4692 = ~n4688 & n4691;
  assign n4698 = x961 & ~n4683;
  assign n4699 = n4691 & n4698;
  assign n4700 = x961 & x962;
  assign n4701 = ~n4699 & ~n4700;
  assign n4693 = ~x963 & ~x964;
  assign n4694 = ~n4685 & n4693;
  assign n4702 = ~n4683 & ~n4686;
  assign n4703 = ~n4694 & n4702;
  assign n4704 = ~x966 & n4686;
  assign n4705 = x962 & ~n4704;
  assign n4706 = ~n4703 & n4705;
  assign n4707 = ~n4701 & ~n4706;
  assign n6054 = ~n4692 & ~n4707;
  assign n6056 = n6055 ^ n6054;
  assign n4729 = ~n4718 & n4728;
  assign n4730 = ~n4726 & ~n4729;
  assign n4731 = ~x955 & ~n4730;
  assign n4742 = ~n4731 & ~n4741;
  assign n4743 = x955 & ~n4727;
  assign n4744 = ~x956 & ~x960;
  assign n4745 = ~n4720 & n4744;
  assign n4746 = ~n4743 & n4745;
  assign n4747 = n4720 & n4734;
  assign n4748 = ~n4746 & ~n4747;
  assign n4749 = ~x959 & ~n4748;
  assign n4750 = n4742 & ~n4749;
  assign n4695 = ~n4684 & n4694;
  assign n4696 = ~n4692 & ~n4695;
  assign n4697 = ~x961 & ~n4696;
  assign n4708 = ~n4697 & ~n4707;
  assign n4709 = x961 & ~n4693;
  assign n4710 = ~x962 & ~x966;
  assign n4711 = ~n4686 & n4710;
  assign n4712 = ~n4709 & n4711;
  assign n4713 = n4686 & n4700;
  assign n4714 = ~n4712 & ~n4713;
  assign n4715 = ~x965 & ~n4714;
  assign n4716 = n4708 & ~n4715;
  assign n4751 = n4750 ^ n4716;
  assign n4565 = x960 ^ x959;
  assign n4566 = n4565 ^ n4564;
  assign n4563 = x956 ^ x955;
  assign n4567 = n4566 ^ n4563;
  assign n4570 = x966 ^ x965;
  assign n4571 = n4570 ^ n4569;
  assign n4568 = x962 ^ x961;
  assign n4572 = n4571 ^ n4568;
  assign n4674 = n4567 & n4572;
  assign n6051 = n4716 ^ n4674;
  assign n6052 = n4751 & ~n6051;
  assign n6053 = n6052 ^ n4750;
  assign n6057 = n6056 ^ n6053;
  assign n4653 = x950 & ~n4647;
  assign n4654 = ~n4644 & n4646;
  assign n4655 = ~n4653 & n4654;
  assign n4656 = n4652 & ~n4655;
  assign n4657 = ~x949 & ~n4656;
  assign n4575 = x952 ^ x951;
  assign n4577 = n4576 ^ n4575;
  assign n4666 = ~x950 & ~x954;
  assign n4667 = ~n4643 & n4666;
  assign n4668 = n4577 & n4667;
  assign n4669 = ~n4660 & ~n4668;
  assign n4670 = ~x953 & ~n4669;
  assign n4671 = n4665 & ~n4670;
  assign n4672 = ~n4657 & n4671;
  assign n4623 = x944 & ~n4617;
  assign n4624 = ~n4614 & n4616;
  assign n4625 = ~n4623 & n4624;
  assign n4626 = n4622 & ~n4625;
  assign n4627 = ~x943 & ~n4626;
  assign n4580 = x946 ^ x945;
  assign n4582 = n4581 ^ n4580;
  assign n4636 = ~x944 & ~x948;
  assign n4637 = ~n4613 & n4636;
  assign n4638 = n4582 & n4637;
  assign n4639 = ~n4630 & ~n4638;
  assign n4640 = ~x947 & ~n4639;
  assign n4641 = n4635 & ~n4640;
  assign n4642 = ~n4627 & n4641;
  assign n4673 = n4672 ^ n4642;
  assign n4574 = x954 ^ x953;
  assign n4578 = n4577 ^ n4574;
  assign n4579 = x948 ^ x947;
  assign n4583 = n4582 ^ n4579;
  assign n4677 = n4578 & n4583;
  assign n6044 = n4677 ^ n4672;
  assign n6045 = ~n4673 & n6044;
  assign n6046 = n6045 ^ n4677;
  assign n6290 = n6057 ^ n6046;
  assign n4675 = ~n4578 & ~n4583;
  assign n4676 = ~n4674 & n4675;
  assign n4678 = ~n4567 & ~n4572;
  assign n4679 = ~n4677 & n4678;
  assign n4680 = ~n4676 & ~n4679;
  assign n4681 = n4674 & n4677;
  assign n4682 = n4680 & ~n4681;
  assign n4752 = n4751 ^ n4682;
  assign n6059 = ~n4673 & n4752;
  assign n6060 = n4673 & n4677;
  assign n6061 = ~n4680 & ~n4751;
  assign n6062 = ~n6060 & ~n6061;
  assign n6063 = ~n6059 & n6062;
  assign n6064 = n4674 & n4751;
  assign n6065 = n6063 & ~n6064;
  assign n6291 = n6065 ^ n6057;
  assign n6292 = ~n6290 & n6291;
  assign n6293 = n6292 ^ n6065;
  assign n6294 = n6289 & ~n6293;
  assign n6295 = ~n6046 & ~n6065;
  assign n6296 = n6057 & ~n6295;
  assign n6049 = n6048 ^ n6047;
  assign n6050 = n6049 ^ n6046;
  assign n6058 = n6057 ^ n6050;
  assign n6066 = n6065 ^ n6058;
  assign n6297 = ~n6066 & ~n6289;
  assign n6298 = n6296 & n6297;
  assign n6300 = ~n6057 & ~n6299;
  assign n6301 = n6295 & n6300;
  assign n6302 = ~n6298 & ~n6301;
  assign n6303 = ~n6294 & n6302;
  assign n6286 = n6055 ^ n6053;
  assign n6287 = ~n6056 & ~n6286;
  assign n6288 = n6287 ^ n6053;
  assign n6304 = n6303 ^ n6288;
  assign n6498 = ~n6299 & n6304;
  assign n6499 = ~n6288 & ~n6293;
  assign n6500 = ~n6498 & ~n6499;
  assign n6505 = n6504 ^ n6500;
  assign n4889 = n4888 ^ n4816;
  assign n4584 = n4583 ^ n4578;
  assign n4573 = n4572 ^ n4567;
  assign n4585 = n4584 ^ n4573;
  assign n4607 = n4606 ^ n4601;
  assign n4596 = n4595 ^ n4590;
  assign n4608 = n4607 ^ n4596;
  assign n4754 = n4585 & n4608;
  assign n4890 = n4889 ^ n4754;
  assign n4753 = n4752 ^ n4673;
  assign n6041 = n4754 ^ n4753;
  assign n6042 = n4890 & ~n6041;
  assign n6043 = n6042 ^ n4889;
  assign n6067 = n6066 ^ n6043;
  assign n6305 = n6090 ^ n6066;
  assign n6306 = ~n6067 & n6305;
  assign n6307 = n6306 ^ n6090;
  assign n6324 = n6323 ^ n6307;
  assign n6495 = n6307 ^ n6304;
  assign n6496 = n6324 & ~n6495;
  assign n6497 = n6496 ^ n6323;
  assign n6577 = n6500 ^ n6497;
  assign n6578 = n6505 & ~n6577;
  assign n6579 = n6578 ^ n6504;
  assign n6506 = n6505 ^ n6497;
  assign n6251 = n6250 ^ n6227;
  assign n6284 = n6283 ^ n6251;
  assign n6091 = n6090 ^ n6067;
  assign n5333 = n5332 ^ n5135;
  assign n4562 = n4561 ^ n4522;
  assign n4609 = n4608 ^ n4585;
  assign n4610 = n4609 ^ n4522;
  assign n4611 = n4562 & ~n4610;
  assign n4612 = n4611 ^ n4561;
  assign n4891 = n4890 ^ n4753;
  assign n6036 = ~n4612 & ~n4891;
  assign n6037 = ~n6035 & ~n6036;
  assign n6034 = n4612 & n4891;
  assign n6038 = n6037 ^ n6034;
  assign n6039 = ~n5333 & n6038;
  assign n6040 = n6039 ^ n6037;
  assign n6092 = n6091 ^ n6040;
  assign n6196 = n6195 ^ n6152;
  assign n6222 = n6196 ^ n6040;
  assign n6223 = ~n6092 & ~n6222;
  assign n6224 = n6223 ^ n6196;
  assign n6285 = n6284 ^ n6224;
  assign n6325 = n6324 ^ n6304;
  assign n6492 = n6325 ^ n6224;
  assign n6493 = ~n6285 & n6492;
  assign n6494 = n6493 ^ n6284;
  assign n6507 = n6506 ^ n6494;
  assign n6556 = n6555 ^ n6531;
  assign n6580 = n6556 ^ n6494;
  assign n6581 = ~n6507 & n6580;
  assign n6582 = n6581 ^ n6556;
  assign n6620 = n6579 & n6582;
  assign n6621 = n6615 & n6620;
  assign n6583 = n6582 ^ n6579;
  assign n6616 = n6579 ^ n6576;
  assign n6617 = n6583 & ~n6616;
  assign n6618 = n6617 ^ n6582;
  assign n6619 = ~n6615 & ~n6618;
  assign n5542 = x863 & x864;
  assign n5543 = x861 & x862;
  assign n5544 = ~n5542 & ~n5543;
  assign n5545 = ~x863 & ~x864;
  assign n5546 = ~x861 & ~x862;
  assign n5547 = ~n5545 & ~n5546;
  assign n5548 = ~n5544 & n5547;
  assign n5549 = x860 & n5548;
  assign n5550 = n5542 & n5543;
  assign n5551 = ~n5549 & ~n5550;
  assign n5364 = x860 ^ x859;
  assign n5558 = n5364 & n5548;
  assign n5552 = n5544 & ~n5547;
  assign n5559 = x859 & x860;
  assign n5560 = n5543 & n5559;
  assign n5561 = x864 & n5560;
  assign n5562 = n5561 ^ n5559;
  assign n5563 = ~n5552 & n5562;
  assign n5564 = ~n5558 & ~n5563;
  assign n5956 = n5551 & n5564;
  assign n5513 = x869 & x870;
  assign n5514 = x867 & x868;
  assign n5515 = ~n5513 & ~n5514;
  assign n5516 = ~x869 & ~x870;
  assign n5517 = ~x867 & ~x868;
  assign n5518 = ~n5516 & ~n5517;
  assign n5519 = ~n5515 & n5518;
  assign n5520 = x866 & n5519;
  assign n5521 = n5513 & n5514;
  assign n5522 = ~n5520 & ~n5521;
  assign n5369 = x866 ^ x865;
  assign n5529 = n5369 & n5519;
  assign n5523 = n5515 & ~n5518;
  assign n5530 = x865 & x866;
  assign n5531 = n5514 & n5530;
  assign n5532 = x870 & n5531;
  assign n5533 = n5532 ^ n5530;
  assign n5534 = ~n5523 & n5533;
  assign n5535 = ~n5529 & ~n5534;
  assign n5955 = n5522 & n5535;
  assign n5957 = n5956 ^ n5955;
  assign n5553 = ~x860 & n5552;
  assign n5554 = n5545 & n5546;
  assign n5555 = ~n5553 & ~n5554;
  assign n5556 = n5551 & n5555;
  assign n5557 = ~x859 & ~n5556;
  assign n5565 = ~x860 & ~x864;
  assign n5566 = n5546 & n5565;
  assign n5567 = ~n5560 & ~n5566;
  assign n5568 = ~x863 & ~n5567;
  assign n5569 = n5564 & ~n5568;
  assign n5570 = ~n5557 & n5569;
  assign n5524 = ~x866 & n5523;
  assign n5525 = n5516 & n5517;
  assign n5526 = ~n5524 & ~n5525;
  assign n5527 = n5522 & n5526;
  assign n5528 = ~x865 & ~n5527;
  assign n5536 = ~x866 & ~x870;
  assign n5537 = n5517 & n5536;
  assign n5538 = ~n5531 & ~n5537;
  assign n5539 = ~x869 & ~n5538;
  assign n5540 = n5535 & ~n5539;
  assign n5541 = ~n5528 & n5540;
  assign n5571 = n5570 ^ n5541;
  assign n5363 = x862 ^ x861;
  assign n5365 = n5364 ^ n5363;
  assign n5362 = x864 ^ x863;
  assign n5366 = n5365 ^ n5362;
  assign n5368 = x868 ^ x867;
  assign n5370 = n5369 ^ n5368;
  assign n5367 = x870 ^ x869;
  assign n5371 = n5370 ^ n5367;
  assign n5511 = n5366 & n5371;
  assign n5952 = n5541 ^ n5511;
  assign n5953 = n5571 & ~n5952;
  assign n5954 = n5953 ^ n5570;
  assign n5958 = n5957 ^ n5954;
  assign n5375 = x854 ^ x853;
  assign n5374 = x856 ^ x855;
  assign n5597 = x857 & x858;
  assign n5598 = n5597 ^ x856;
  assign n5599 = n5374 & ~n5598;
  assign n5600 = n5599 ^ x855;
  assign n5601 = n5375 & n5600;
  assign n5602 = ~x855 & ~x856;
  assign n5603 = ~n5597 & n5602;
  assign n5604 = x855 & x856;
  assign n5605 = x853 & x854;
  assign n5606 = ~n5604 & n5605;
  assign n5607 = ~n5603 & n5606;
  assign n5608 = ~n5601 & ~n5607;
  assign n5609 = ~x857 & ~x858;
  assign n5610 = ~n5608 & ~n5609;
  assign n5611 = n5604 & n5605;
  assign n5612 = ~x858 & n5611;
  assign n5613 = ~n5610 & ~n5612;
  assign n5376 = n5375 ^ n5374;
  assign n5614 = ~x854 & ~x858;
  assign n5615 = ~n5604 & n5614;
  assign n5616 = n5376 & n5615;
  assign n5617 = ~n5611 & ~n5616;
  assign n5618 = ~x857 & ~n5617;
  assign n5619 = n5613 & ~n5618;
  assign n5620 = x854 & ~n5609;
  assign n5621 = n5597 & n5604;
  assign n5622 = ~n5620 & ~n5621;
  assign n5623 = n5600 & ~n5622;
  assign n5624 = n5603 & ~n5620;
  assign n5625 = ~n5623 & ~n5624;
  assign n5626 = ~x853 & ~n5625;
  assign n5627 = n5619 & ~n5626;
  assign n5574 = ~x851 & ~x852;
  assign n5575 = ~x849 & ~x850;
  assign n5576 = ~n5574 & ~n5575;
  assign n5577 = x851 & x852;
  assign n5578 = x849 & x850;
  assign n5579 = ~n5577 & ~n5578;
  assign n5580 = n5576 & ~n5579;
  assign n5581 = x848 & n5580;
  assign n5582 = n5577 & n5578;
  assign n5583 = ~n5581 & ~n5582;
  assign n5584 = ~n5576 & n5579;
  assign n5585 = ~x848 & n5584;
  assign n5586 = n5583 & ~n5585;
  assign n5587 = ~x847 & ~n5586;
  assign n5588 = ~n5582 & ~n5584;
  assign n5589 = x848 & ~n5588;
  assign n5590 = ~x848 & ~n5580;
  assign n5591 = x847 & ~n5590;
  assign n5592 = ~n5589 & n5591;
  assign n5380 = x848 ^ x847;
  assign n5593 = n5574 & n5575;
  assign n5594 = n5380 & n5593;
  assign n5595 = ~n5592 & ~n5594;
  assign n5596 = ~n5587 & n5595;
  assign n5628 = n5627 ^ n5596;
  assign n5373 = x858 ^ x857;
  assign n5377 = n5376 ^ n5373;
  assign n5379 = x850 ^ x849;
  assign n5381 = n5380 ^ n5379;
  assign n5378 = x852 ^ x851;
  assign n5382 = n5381 ^ n5378;
  assign n5573 = n5377 & n5382;
  assign n5960 = n5596 ^ n5573;
  assign n5961 = n5628 & ~n5960;
  assign n5962 = n5961 ^ n5627;
  assign n5372 = n5371 ^ n5366;
  assign n5383 = n5382 ^ n5377;
  assign n5510 = n5372 & n5383;
  assign n5512 = ~n5510 & ~n5511;
  assign n5572 = n5571 ^ n5512;
  assign n5629 = n5628 ^ n5573;
  assign n5963 = ~n5572 & n5629;
  assign n5964 = n5510 & n5571;
  assign n5965 = ~n5963 & ~n5964;
  assign n6334 = ~n5962 & n5965;
  assign n6335 = n5958 & ~n6334;
  assign n6336 = n5962 & ~n5965;
  assign n6337 = ~n6335 & ~n6336;
  assign n5949 = n5583 & ~n5592;
  assign n5950 = n5613 & ~n5623;
  assign n6338 = ~n5949 & ~n5950;
  assign n6339 = ~n5958 & ~n6338;
  assign n6340 = n6334 & n6339;
  assign n6341 = n5949 & n5950;
  assign n6342 = ~n6340 & ~n6341;
  assign n6343 = n6337 & ~n6342;
  assign n6344 = n6335 & n6338;
  assign n6345 = n5958 & ~n6341;
  assign n6346 = n6336 & n6345;
  assign n6347 = ~n6344 & ~n6346;
  assign n6348 = ~n6343 & n6347;
  assign n6331 = n5956 ^ n5954;
  assign n6332 = ~n5957 & ~n6331;
  assign n6333 = n6332 ^ n5954;
  assign n6349 = n6348 ^ n6333;
  assign n5966 = n5965 ^ n5962;
  assign n5951 = n5950 ^ n5949;
  assign n5959 = n5958 ^ n5951;
  assign n5967 = n5966 ^ n5959;
  assign n5475 = x875 & x876;
  assign n5476 = x873 & x874;
  assign n5477 = ~n5475 & ~n5476;
  assign n5478 = ~x875 & ~x876;
  assign n5479 = ~x873 & ~x874;
  assign n5480 = ~n5478 & ~n5479;
  assign n5481 = n5477 & ~n5480;
  assign n5482 = x871 & x872;
  assign n5483 = n5476 & n5482;
  assign n5484 = x876 & n5483;
  assign n5485 = n5484 ^ n5482;
  assign n5486 = ~n5481 & n5485;
  assign n5487 = n5475 & n5476;
  assign n5488 = ~n5486 & ~n5487;
  assign n5489 = ~n5477 & n5480;
  assign n5490 = ~x872 & n5489;
  assign n5491 = ~x871 & n5490;
  assign n5492 = n5491 ^ n5489;
  assign n5493 = n5488 & ~n5492;
  assign n5494 = x872 & ~n5478;
  assign n5495 = ~n5475 & n5479;
  assign n5496 = ~n5494 & n5495;
  assign n5497 = n5493 & ~n5496;
  assign n5498 = x871 & ~n5486;
  assign n5499 = ~n5490 & n5498;
  assign n5500 = ~n5497 & ~n5499;
  assign n5348 = x872 ^ x871;
  assign n5347 = x874 ^ x873;
  assign n5349 = n5348 ^ n5347;
  assign n5501 = ~x872 & ~x876;
  assign n5502 = ~n5476 & n5501;
  assign n5503 = n5349 & n5502;
  assign n5504 = ~n5483 & ~n5503;
  assign n5505 = ~x875 & ~n5504;
  assign n5506 = ~n5500 & ~n5505;
  assign n5452 = ~x881 & ~x882;
  assign n5453 = ~x879 & ~x880;
  assign n5454 = ~n5452 & ~n5453;
  assign n5455 = x881 & x882;
  assign n5456 = x879 & x880;
  assign n5457 = ~n5455 & ~n5456;
  assign n5458 = n5454 & ~n5457;
  assign n5459 = x878 & n5458;
  assign n5460 = n5455 & n5456;
  assign n5461 = ~n5459 & ~n5460;
  assign n5462 = ~n5454 & n5457;
  assign n5463 = ~x878 & n5462;
  assign n5464 = n5461 & ~n5463;
  assign n5465 = ~x877 & ~n5464;
  assign n5466 = ~n5460 & ~n5462;
  assign n5467 = x878 & ~n5466;
  assign n5468 = ~x878 & ~n5458;
  assign n5469 = x877 & ~n5468;
  assign n5470 = ~n5467 & n5469;
  assign n5353 = x878 ^ x877;
  assign n5471 = n5452 & n5453;
  assign n5472 = n5353 & n5471;
  assign n5473 = ~n5470 & ~n5472;
  assign n5474 = ~n5465 & n5473;
  assign n5507 = n5506 ^ n5474;
  assign n5420 = x887 & x888;
  assign n5421 = x885 & x886;
  assign n5422 = n5420 & n5421;
  assign n5423 = ~n5420 & ~n5421;
  assign n5424 = ~x887 & ~x888;
  assign n5425 = ~x885 & ~x886;
  assign n5426 = ~n5424 & ~n5425;
  assign n5427 = ~n5423 & n5426;
  assign n5428 = ~x884 & n5427;
  assign n5429 = ~x883 & n5428;
  assign n5430 = n5429 ^ n5427;
  assign n5431 = ~n5422 & ~n5430;
  assign n5432 = x884 & ~n5424;
  assign n5433 = ~n5420 & n5425;
  assign n5434 = ~n5432 & n5433;
  assign n5435 = n5431 & ~n5434;
  assign n5436 = x883 & ~n5428;
  assign n5437 = ~n5435 & ~n5436;
  assign n5342 = x884 ^ x883;
  assign n5341 = x886 ^ x885;
  assign n5343 = n5342 ^ n5341;
  assign n5438 = ~x884 & ~x888;
  assign n5439 = ~n5421 & n5438;
  assign n5440 = n5343 & n5439;
  assign n5441 = x883 & x884;
  assign n5442 = n5421 & n5441;
  assign n5443 = ~n5440 & ~n5442;
  assign n5444 = ~x887 & ~n5443;
  assign n5445 = n5423 & ~n5426;
  assign n5446 = x888 & n5442;
  assign n5447 = n5446 ^ n5441;
  assign n5448 = ~n5445 & n5447;
  assign n5449 = ~n5444 & ~n5448;
  assign n5450 = ~n5437 & n5449;
  assign n5397 = x893 & x894;
  assign n5398 = x891 & x892;
  assign n5399 = ~n5397 & ~n5398;
  assign n5400 = ~x893 & ~x894;
  assign n5401 = ~x891 & ~x892;
  assign n5402 = ~n5400 & ~n5401;
  assign n5403 = ~n5399 & n5402;
  assign n5404 = x890 & n5403;
  assign n5405 = n5397 & n5398;
  assign n5406 = ~n5404 & ~n5405;
  assign n5407 = n5399 & ~n5402;
  assign n5408 = ~x890 & n5407;
  assign n5409 = n5406 & ~n5408;
  assign n5410 = ~x889 & ~n5409;
  assign n5411 = ~n5405 & ~n5407;
  assign n5412 = x890 & ~n5411;
  assign n5413 = ~x890 & ~n5403;
  assign n5414 = x889 & ~n5413;
  assign n5415 = ~n5412 & n5414;
  assign n5337 = x890 ^ x889;
  assign n5416 = n5400 & n5401;
  assign n5417 = n5337 & n5416;
  assign n5418 = ~n5415 & ~n5417;
  assign n5419 = ~n5410 & n5418;
  assign n5451 = n5450 ^ n5419;
  assign n5508 = n5507 ^ n5451;
  assign n5336 = x892 ^ x891;
  assign n5338 = n5337 ^ n5336;
  assign n5335 = x894 ^ x893;
  assign n5339 = n5338 ^ n5335;
  assign n5340 = x888 ^ x887;
  assign n5344 = n5343 ^ n5340;
  assign n5345 = n5339 & n5344;
  assign n5352 = x880 ^ x879;
  assign n5354 = n5353 ^ n5352;
  assign n5351 = x882 ^ x881;
  assign n5355 = n5354 ^ n5351;
  assign n5346 = x876 ^ x875;
  assign n5350 = n5349 ^ n5346;
  assign n5356 = n5355 ^ n5350;
  assign n5357 = n5344 ^ n5339;
  assign n5358 = n5357 ^ n5350;
  assign n5359 = n5356 & ~n5358;
  assign n5360 = n5359 ^ n5355;
  assign n5361 = ~n5345 & ~n5360;
  assign n5384 = n5383 ^ n5372;
  assign n5385 = n5357 ^ n5356;
  assign n5386 = n5384 & n5385;
  assign n5387 = ~n5361 & n5386;
  assign n5388 = ~n5350 & ~n5355;
  assign n5389 = ~n5339 & ~n5344;
  assign n5390 = n5388 & n5389;
  assign n5391 = ~n5387 & ~n5390;
  assign n5392 = n5361 & ~n5384;
  assign n5393 = n5350 & n5355;
  assign n5394 = n5345 & n5393;
  assign n5395 = ~n5392 & ~n5394;
  assign n5396 = n5391 & n5395;
  assign n5509 = n5508 ^ n5396;
  assign n5630 = n5629 ^ n5572;
  assign n5946 = n5630 ^ n5386;
  assign n5947 = ~n5509 & ~n5946;
  assign n5948 = n5947 ^ n5630;
  assign n5968 = n5967 ^ n5948;
  assign n5936 = n5360 & ~n5507;
  assign n5937 = ~n5345 & ~n5451;
  assign n5938 = n5936 & ~n5937;
  assign n5939 = ~n5393 & n5507;
  assign n5940 = ~n5938 & ~n5939;
  assign n5941 = n5361 ^ n5345;
  assign n5942 = ~n5451 & n5941;
  assign n5943 = n5942 ^ n5345;
  assign n5944 = ~n5940 & ~n5943;
  assign n5931 = ~n5345 & n5451;
  assign n5932 = ~n5419 & ~n5450;
  assign n5933 = ~n5931 & ~n5932;
  assign n5928 = n5461 & ~n5470;
  assign n5929 = n5928 ^ n5493;
  assign n5926 = n5406 & ~n5415;
  assign n5925 = n5431 & ~n5448;
  assign n5927 = n5926 ^ n5925;
  assign n5930 = n5929 ^ n5927;
  assign n5934 = n5933 ^ n5930;
  assign n5922 = n5474 ^ n5393;
  assign n5923 = n5507 & ~n5922;
  assign n5924 = n5923 ^ n5506;
  assign n5935 = n5934 ^ n5924;
  assign n5945 = n5944 ^ n5935;
  assign n6328 = n5948 ^ n5945;
  assign n6329 = n5968 & n6328;
  assign n6330 = n6329 ^ n5967;
  assign n6350 = n6349 ^ n6330;
  assign n6351 = ~n5924 & n5928;
  assign n6352 = n5933 ^ n5926;
  assign n6353 = ~n5927 & ~n6352;
  assign n6354 = n6353 ^ n5933;
  assign n6355 = n6351 & ~n6354;
  assign n6356 = ~n5926 & n5933;
  assign n6357 = ~n5925 & n6356;
  assign n6358 = ~n5928 & n6357;
  assign n6359 = ~n6355 & ~n6358;
  assign n6360 = n5493 & ~n6359;
  assign n6361 = ~n5493 & ~n6357;
  assign n6362 = n5925 & n5926;
  assign n6363 = ~n5933 & n6362;
  assign n6364 = n5493 & ~n6363;
  assign n6365 = n5924 & ~n5928;
  assign n6366 = ~n6364 & ~n6365;
  assign n6367 = ~n6361 & n6366;
  assign n6368 = n6351 & n6363;
  assign n6369 = ~n6367 & ~n6368;
  assign n6370 = ~n6360 & n6369;
  assign n6371 = ~n5924 & ~n5944;
  assign n6372 = n6370 & n6371;
  assign n6373 = n5493 & n5928;
  assign n6374 = ~n6357 & ~n6373;
  assign n6375 = n6354 & n6374;
  assign n6376 = ~n5493 & ~n5928;
  assign n6377 = ~n6363 & n6376;
  assign n6378 = ~n6356 & n6377;
  assign n6379 = n6357 & n6373;
  assign n6380 = ~n6378 & ~n6379;
  assign n6381 = ~n6375 & n6380;
  assign n6382 = n5944 & n6381;
  assign n6383 = ~n6372 & ~n6382;
  assign n6384 = n5934 & ~n6383;
  assign n6385 = n5924 & n5944;
  assign n6386 = n6385 ^ n6370;
  assign n6387 = n6381 & n6386;
  assign n6388 = ~n6384 & ~n6387;
  assign n6481 = n6388 ^ n6349;
  assign n6482 = n6350 & ~n6481;
  assign n6483 = n6482 ^ n6388;
  assign n5823 = x909 & x910;
  assign n5824 = x911 & x912;
  assign n5825 = ~n5823 & ~n5824;
  assign n5826 = ~x909 & ~x910;
  assign n5827 = ~x911 & ~x912;
  assign n5828 = ~n5826 & ~n5827;
  assign n5829 = ~n5825 & n5828;
  assign n5830 = x908 & n5829;
  assign n5831 = n5823 & n5824;
  assign n5832 = ~n5830 & ~n5831;
  assign n5833 = n5825 & ~n5828;
  assign n5834 = ~x908 & n5833;
  assign n5835 = n5832 & ~n5834;
  assign n5836 = ~x907 & ~n5835;
  assign n5837 = ~n5831 & ~n5833;
  assign n5838 = x908 & ~n5837;
  assign n5839 = ~x908 & ~n5829;
  assign n5840 = x907 & ~n5839;
  assign n5841 = ~n5838 & n5840;
  assign n5650 = x908 ^ x907;
  assign n5842 = n5826 & n5827;
  assign n5843 = n5650 & n5842;
  assign n5844 = ~n5841 & ~n5843;
  assign n5845 = ~n5836 & n5844;
  assign n5792 = x915 & x916;
  assign n5793 = x917 & x918;
  assign n5794 = ~n5792 & ~n5793;
  assign n5795 = ~x915 & ~x916;
  assign n5796 = ~x917 & ~x918;
  assign n5797 = ~n5795 & ~n5796;
  assign n5798 = ~n5794 & n5797;
  assign n5799 = x914 & n5798;
  assign n5800 = n5792 & n5793;
  assign n5801 = ~n5799 & ~n5800;
  assign n5802 = x914 & ~n5796;
  assign n5803 = ~n5793 & n5795;
  assign n5804 = ~n5802 & n5803;
  assign n5805 = n5801 & ~n5804;
  assign n5806 = ~x913 & ~n5805;
  assign n5807 = x913 & ~n5795;
  assign n5808 = ~x914 & ~x918;
  assign n5809 = ~n5792 & n5808;
  assign n5810 = ~n5807 & n5809;
  assign n5811 = x913 & x914;
  assign n5812 = n5792 & n5811;
  assign n5813 = ~n5810 & ~n5812;
  assign n5814 = ~x917 & ~n5813;
  assign n5645 = x914 ^ x913;
  assign n5815 = n5645 & n5798;
  assign n5816 = n5794 & ~n5797;
  assign n5817 = x918 & n5812;
  assign n5818 = n5817 ^ n5811;
  assign n5819 = ~n5816 & n5818;
  assign n5820 = ~n5815 & ~n5819;
  assign n5821 = ~n5814 & n5820;
  assign n5822 = ~n5806 & n5821;
  assign n5846 = n5845 ^ n5822;
  assign n5878 = x899 & x900;
  assign n5879 = x897 & x898;
  assign n5880 = ~n5878 & ~n5879;
  assign n5881 = ~x899 & ~x900;
  assign n5882 = ~x897 & ~x898;
  assign n5883 = ~n5881 & ~n5882;
  assign n5884 = ~n5880 & n5883;
  assign n5885 = x896 & n5884;
  assign n5886 = n5878 & n5879;
  assign n5887 = ~n5885 & ~n5886;
  assign n5888 = n5880 & ~n5883;
  assign n5889 = ~x896 & n5888;
  assign n5890 = n5887 & ~n5889;
  assign n5891 = ~x895 & ~n5890;
  assign n5892 = ~n5886 & ~n5888;
  assign n5893 = x896 & ~n5892;
  assign n5894 = ~x896 & ~n5884;
  assign n5895 = x895 & ~n5894;
  assign n5896 = ~n5893 & n5895;
  assign n5639 = x896 ^ x895;
  assign n5897 = n5881 & n5882;
  assign n5898 = n5639 & n5897;
  assign n5899 = ~n5896 & ~n5898;
  assign n5900 = ~n5891 & n5899;
  assign n5633 = x904 ^ x903;
  assign n5855 = x905 & x906;
  assign n5856 = n5855 ^ x904;
  assign n5857 = ~n5633 & ~n5856;
  assign n5858 = ~x901 & n5857;
  assign n5859 = x903 & x904;
  assign n5860 = ~x905 & ~x906;
  assign n5861 = ~n5859 & n5860;
  assign n5862 = ~x902 & n5861;
  assign n5863 = ~n5858 & ~n5862;
  assign n5864 = ~x903 & ~x904;
  assign n5865 = x901 & ~n5864;
  assign n5866 = x902 & ~n5860;
  assign n5867 = ~n5865 & ~n5866;
  assign n5868 = ~n5863 & n5867;
  assign n5634 = x902 ^ x901;
  assign n5869 = n5855 & ~n5864;
  assign n5870 = n5859 & ~n5860;
  assign n5871 = ~n5869 & ~n5870;
  assign n5872 = n5634 & ~n5871;
  assign n5873 = x901 & x902;
  assign n5874 = ~n5861 & n5873;
  assign n5875 = ~n5857 & n5874;
  assign n5876 = ~n5872 & ~n5875;
  assign n5877 = ~n5868 & n5876;
  assign n5901 = n5900 ^ n5877;
  assign n5644 = x918 ^ x917;
  assign n5646 = n5645 ^ n5644;
  assign n5643 = x916 ^ x915;
  assign n5647 = n5646 ^ n5643;
  assign n5649 = x912 ^ x911;
  assign n5651 = n5650 ^ n5649;
  assign n5648 = x910 ^ x909;
  assign n5652 = n5651 ^ n5648;
  assign n5847 = n5647 & n5652;
  assign n5635 = n5634 ^ n5633;
  assign n5632 = x906 ^ x905;
  assign n5636 = n5635 ^ n5632;
  assign n5638 = x898 ^ x897;
  assign n5640 = n5639 ^ n5638;
  assign n5637 = x900 ^ x899;
  assign n5641 = n5640 ^ n5637;
  assign n5851 = n5636 & n5641;
  assign n5642 = n5641 ^ n5636;
  assign n5653 = n5652 ^ n5647;
  assign n5848 = n5653 ^ n5641;
  assign n5849 = ~n5642 & n5848;
  assign n5850 = n5849 ^ n5653;
  assign n5852 = n5851 ^ n5850;
  assign n5853 = ~n5847 & ~n5852;
  assign n5854 = n5853 ^ n5851;
  assign n5902 = n5901 ^ n5854;
  assign n5990 = ~n5846 & ~n5902;
  assign n5991 = ~n5850 & ~n5901;
  assign n5992 = n5846 & n5847;
  assign n5993 = ~n5991 & ~n5992;
  assign n5994 = ~n5990 & n5993;
  assign n5995 = n5851 & n5901;
  assign n5996 = n5994 & ~n5995;
  assign n5977 = n5801 & n5820;
  assign n5984 = n5847 ^ n5845;
  assign n5985 = ~n5846 & n5984;
  assign n5986 = n5985 ^ n5847;
  assign n5987 = n5832 & ~n5841;
  assign n6422 = ~n5986 & n5987;
  assign n6423 = n5977 & n6422;
  assign n6424 = n5986 & ~n5987;
  assign n5978 = n5855 & n5859;
  assign n5979 = n5876 & ~n5978;
  assign n5980 = n5887 & ~n5896;
  assign n6425 = ~n5979 & ~n5980;
  assign n6426 = ~n6424 & n6425;
  assign n6427 = ~n6423 & n6426;
  assign n5988 = n5987 ^ n5986;
  assign n5981 = n5980 ^ n5979;
  assign n6428 = ~n5977 & n5981;
  assign n6429 = ~n5988 & n6428;
  assign n6430 = n5979 & n5980;
  assign n6431 = n6430 ^ n5977;
  assign n6432 = n6424 & n6431;
  assign n6433 = ~n6429 & ~n6432;
  assign n6434 = ~n6427 & n6433;
  assign n5974 = n5877 ^ n5851;
  assign n5975 = n5901 & ~n5974;
  assign n5976 = n5975 ^ n5900;
  assign n5982 = n5981 ^ n5977;
  assign n5983 = n5982 ^ n5976;
  assign n5989 = n5988 ^ n5983;
  assign n6435 = ~n5976 & n5989;
  assign n6436 = n6434 & n6435;
  assign n6437 = n6423 & n6430;
  assign n6438 = ~n5977 & n6424;
  assign n6439 = n5981 & n6438;
  assign n6440 = ~n6437 & ~n6439;
  assign n6441 = n5976 & ~n6440;
  assign n6442 = ~n6436 & ~n6441;
  assign n6443 = n5996 & ~n6442;
  assign n6444 = n5989 & n5996;
  assign n6445 = n6440 & ~n6444;
  assign n6446 = n6435 ^ n6434;
  assign n6447 = n6445 & n6446;
  assign n6448 = ~n6443 & ~n6447;
  assign n5997 = n5996 ^ n5989;
  assign n5766 = x941 & x942;
  assign n5767 = x939 & x940;
  assign n5768 = ~n5766 & ~n5767;
  assign n5769 = ~x941 & ~x942;
  assign n5770 = ~x939 & ~x940;
  assign n5771 = ~n5769 & ~n5770;
  assign n5772 = ~n5768 & n5771;
  assign n5773 = x938 & n5772;
  assign n5774 = n5766 & n5767;
  assign n5775 = ~n5773 & ~n5774;
  assign n5776 = n5768 & ~n5771;
  assign n5777 = ~x938 & n5776;
  assign n5778 = n5775 & ~n5777;
  assign n5779 = ~x937 & ~n5778;
  assign n5780 = ~n5774 & ~n5776;
  assign n5781 = x938 & ~n5780;
  assign n5782 = ~x938 & ~n5772;
  assign n5783 = x937 & ~n5782;
  assign n5784 = ~n5781 & n5783;
  assign n5662 = x938 ^ x937;
  assign n5785 = n5769 & n5770;
  assign n5786 = n5662 & n5785;
  assign n5787 = ~n5784 & ~n5786;
  assign n5788 = ~n5779 & n5787;
  assign n5741 = x933 & x934;
  assign n5742 = ~x935 & ~x936;
  assign n5743 = ~n5741 & n5742;
  assign n5744 = ~x932 & n5743;
  assign n5745 = ~x933 & ~x934;
  assign n5746 = x935 & x936;
  assign n5747 = n5745 & ~n5746;
  assign n5748 = x932 & ~n5742;
  assign n5749 = n5747 & ~n5748;
  assign n5750 = ~n5744 & ~n5749;
  assign n5751 = n5741 & n5746;
  assign n5752 = n5750 & ~n5751;
  assign n5753 = ~x931 & ~n5752;
  assign n5754 = x931 & x932;
  assign n5755 = ~n5747 & n5754;
  assign n5756 = ~n5743 & ~n5751;
  assign n5757 = n5755 & n5756;
  assign n5657 = x932 ^ x931;
  assign n5758 = ~n5745 & n5746;
  assign n5759 = n5741 & ~n5742;
  assign n5760 = ~n5758 & ~n5759;
  assign n5761 = n5657 & ~n5760;
  assign n5762 = ~n5757 & ~n5761;
  assign n5763 = n5744 & n5745;
  assign n5764 = n5762 & ~n5763;
  assign n5765 = ~n5753 & n5764;
  assign n5789 = n5788 ^ n5765;
  assign n5710 = ~x929 & ~x930;
  assign n5711 = ~x927 & ~x928;
  assign n5712 = ~n5710 & ~n5711;
  assign n5713 = x929 & x930;
  assign n5714 = x927 & x928;
  assign n5715 = ~n5713 & ~n5714;
  assign n5716 = n5712 & ~n5715;
  assign n5717 = x926 & n5716;
  assign n5718 = n5713 & n5714;
  assign n5719 = ~n5717 & ~n5718;
  assign n5720 = ~n5712 & n5715;
  assign n5721 = n5710 & n5711;
  assign n5722 = x926 & ~n5721;
  assign n5723 = n5720 & ~n5722;
  assign n5724 = n5719 & ~n5723;
  assign n5725 = ~x925 & ~n5724;
  assign n5673 = x926 ^ x925;
  assign n5726 = n5673 & n5716;
  assign n5727 = x925 & x926;
  assign n5728 = n5714 & n5727;
  assign n5729 = x930 & n5728;
  assign n5730 = n5729 ^ n5727;
  assign n5731 = ~n5720 & n5730;
  assign n5732 = ~n5726 & ~n5731;
  assign n5733 = ~x926 & ~x930;
  assign n5734 = n5711 & n5733;
  assign n5735 = ~n5728 & ~n5734;
  assign n5736 = ~x929 & ~n5735;
  assign n5737 = n5732 & ~n5736;
  assign n5738 = ~n5725 & n5737;
  assign n5668 = x920 ^ x919;
  assign n5687 = ~x921 & ~x922;
  assign n5688 = x923 & x924;
  assign n5689 = ~n5687 & n5688;
  assign n5690 = x921 & x922;
  assign n5691 = ~x923 & ~x924;
  assign n5692 = n5690 & ~n5691;
  assign n5693 = ~n5689 & ~n5692;
  assign n5694 = n5668 & ~n5693;
  assign n5695 = ~n5690 & n5691;
  assign n5696 = x919 & x920;
  assign n5697 = ~n5695 & n5696;
  assign n5667 = x922 ^ x921;
  assign n5698 = n5688 ^ x922;
  assign n5699 = ~n5667 & ~n5698;
  assign n5700 = n5697 & ~n5699;
  assign n5701 = ~n5694 & ~n5700;
  assign n5702 = ~x919 & n5699;
  assign n5703 = ~x920 & n5695;
  assign n5704 = ~n5702 & ~n5703;
  assign n5705 = x919 & ~n5687;
  assign n5706 = x920 & ~n5691;
  assign n5707 = ~n5705 & ~n5706;
  assign n5708 = ~n5704 & n5707;
  assign n5709 = n5701 & ~n5708;
  assign n5739 = n5738 ^ n5709;
  assign n5656 = x934 ^ x933;
  assign n5658 = n5657 ^ n5656;
  assign n5655 = x936 ^ x935;
  assign n5659 = n5658 ^ n5655;
  assign n5661 = x940 ^ x939;
  assign n5663 = n5662 ^ n5661;
  assign n5660 = x942 ^ x941;
  assign n5664 = n5663 ^ n5660;
  assign n5679 = n5659 & n5664;
  assign n5669 = n5668 ^ n5667;
  assign n5666 = x924 ^ x923;
  assign n5670 = n5669 ^ n5666;
  assign n5672 = x928 ^ x927;
  assign n5674 = n5673 ^ n5672;
  assign n5671 = x930 ^ x929;
  assign n5675 = n5674 ^ n5671;
  assign n5683 = n5670 & n5675;
  assign n5676 = n5675 ^ n5670;
  assign n5665 = n5664 ^ n5659;
  assign n5680 = n5670 ^ n5665;
  assign n5681 = n5676 & ~n5680;
  assign n5682 = n5681 ^ n5675;
  assign n5684 = n5683 ^ n5682;
  assign n5685 = ~n5679 & ~n5684;
  assign n5686 = n5685 ^ n5683;
  assign n5740 = n5739 ^ n5686;
  assign n5790 = n5789 ^ n5740;
  assign n5654 = n5653 ^ n5642;
  assign n5677 = n5676 ^ n5665;
  assign n5678 = n5654 & n5677;
  assign n5791 = n5790 ^ n5678;
  assign n5903 = n5902 ^ n5846;
  assign n5971 = n5903 ^ n5678;
  assign n5972 = ~n5791 & n5971;
  assign n5973 = n5972 ^ n5790;
  assign n5998 = n5997 ^ n5973;
  assign n6013 = n5775 & ~n5784;
  assign n6014 = ~n5751 & n5762;
  assign n6015 = ~n6013 & ~n6014;
  assign n6016 = n5765 ^ n5679;
  assign n6017 = n5789 & ~n6016;
  assign n6018 = n6017 ^ n5788;
  assign n6019 = n6015 & n6018;
  assign n6020 = n6018 ^ n6013;
  assign n6021 = n6014 ^ n6013;
  assign n6022 = ~n6020 & ~n6021;
  assign n6023 = n6022 ^ n6018;
  assign n6024 = ~n6019 & n6023;
  assign n6025 = n6013 & n6014;
  assign n6026 = ~n6018 & n6025;
  assign n6027 = ~n6024 & ~n6026;
  assign n6011 = n5719 & n5732;
  assign n6009 = n5688 & n5690;
  assign n6010 = n5701 & ~n6009;
  assign n6012 = n6011 ^ n6010;
  assign n6028 = n6027 ^ n6012;
  assign n6006 = n5709 ^ n5683;
  assign n6007 = n5739 & ~n6006;
  assign n6008 = n6007 ^ n5738;
  assign n6029 = n6028 ^ n6008;
  assign n5999 = n5683 & n5739;
  assign n6000 = ~n5740 & ~n5789;
  assign n6001 = n5679 & n5789;
  assign n6002 = ~n5682 & ~n5739;
  assign n6003 = ~n6001 & ~n6002;
  assign n6004 = ~n6000 & n6003;
  assign n6005 = ~n5999 & n6004;
  assign n6030 = n6029 ^ n6005;
  assign n6419 = n6030 ^ n5997;
  assign n6420 = n5998 & n6419;
  assign n6421 = n6420 ^ n6030;
  assign n6449 = n6448 ^ n6421;
  assign n6393 = n6026 ^ n6019;
  assign n6394 = n6011 & n6393;
  assign n6395 = n6394 ^ n6019;
  assign n6396 = n6029 & n6395;
  assign n6397 = ~n6008 & n6010;
  assign n6398 = ~n6023 & n6397;
  assign n6399 = ~n6011 & ~n6026;
  assign n6400 = n6398 & ~n6399;
  assign n6401 = n6012 & n6019;
  assign n6402 = ~n6400 & ~n6401;
  assign n6403 = ~n6396 & n6402;
  assign n6404 = n6005 & n6029;
  assign n6405 = ~n6008 & n6028;
  assign n6406 = n6010 & n6011;
  assign n6407 = n6024 & ~n6406;
  assign n6408 = ~n6010 & ~n6011;
  assign n6409 = ~n6015 & n6408;
  assign n6410 = ~n6026 & n6409;
  assign n6411 = n6019 & n6406;
  assign n6412 = ~n6410 & ~n6411;
  assign n6413 = ~n6407 & n6412;
  assign n6414 = ~n6405 & ~n6413;
  assign n6415 = ~n6404 & ~n6414;
  assign n6416 = n6415 ^ n6404;
  assign n6417 = n6403 & n6416;
  assign n6418 = n6417 ^ n6404;
  assign n6450 = n6449 ^ n6418;
  assign n5969 = n5968 ^ n5945;
  assign n5907 = n5677 ^ n5654;
  assign n5908 = n5385 ^ n5384;
  assign n5913 = n5907 & n5908;
  assign n5904 = n5903 ^ n5791;
  assign n5918 = n5913 ^ n5904;
  assign n5631 = n5630 ^ n5509;
  assign n5919 = n5913 ^ n5631;
  assign n5920 = n5918 & n5919;
  assign n5921 = n5920 ^ n5904;
  assign n5970 = n5969 ^ n5921;
  assign n6031 = n6030 ^ n5998;
  assign n6390 = n6031 ^ n5969;
  assign n6391 = ~n5970 & ~n6390;
  assign n6392 = n6391 ^ n6031;
  assign n6451 = n6450 ^ n6392;
  assign n6389 = n6388 ^ n6350;
  assign n6484 = n6392 ^ n6389;
  assign n6485 = n6451 & n6484;
  assign n6486 = n6485 ^ n6450;
  assign n6589 = n6483 & n6486;
  assign n6474 = ~n6438 & ~n6448;
  assign n6475 = ~n5976 & n6430;
  assign n6476 = ~n6423 & ~n6475;
  assign n6477 = ~n6474 & n6476;
  assign n6471 = n6448 ^ n6418;
  assign n6472 = ~n6449 & n6471;
  assign n6473 = n6472 ^ n6421;
  assign n6478 = n6477 ^ n6473;
  assign n6467 = ~n6011 & n6018;
  assign n6468 = n6418 & ~n6467;
  assign n6469 = ~n6015 & n6415;
  assign n6470 = ~n6468 & ~n6469;
  assign n6479 = n6478 ^ n6470;
  assign n6459 = ~n6338 & n6349;
  assign n6460 = ~n6333 & n6337;
  assign n6461 = ~n6459 & ~n6460;
  assign n6462 = ~n6376 & n6387;
  assign n6463 = ~n6355 & ~n6363;
  assign n6464 = ~n6462 & n6463;
  assign n6465 = ~n6384 & n6464;
  assign n6595 = n6461 & n6465;
  assign n6597 = ~n6479 & ~n6595;
  assign n6598 = n6589 & n6597;
  assign n6590 = n6479 & ~n6589;
  assign n6596 = n6590 & n6595;
  assign n6591 = ~n6483 & ~n6486;
  assign n6592 = ~n6590 & ~n6591;
  assign n6593 = ~n6461 & ~n6465;
  assign n6594 = n6592 & n6593;
  assign n6586 = n6477 ^ n6470;
  assign n6587 = n6478 & ~n6586;
  assign n6588 = n6587 ^ n6473;
  assign n6599 = n6479 & ~n6593;
  assign n6600 = n6591 & n6599;
  assign n6623 = ~n6588 & ~n6600;
  assign n6624 = ~n6594 & ~n6623;
  assign n6625 = ~n6596 & ~n6624;
  assign n6626 = ~n6598 & ~n6625;
  assign n6637 = ~n6619 & n6626;
  assign n6638 = ~n6621 & ~n6637;
  assign n6584 = n6583 ^ n6576;
  assign n6557 = n6556 ^ n6507;
  assign n6326 = n6325 ^ n6285;
  assign n6032 = n6031 ^ n5970;
  assign n4892 = n4891 ^ n4612;
  assign n5334 = n5333 ^ n4892;
  assign n5905 = n5904 ^ n5631;
  assign n5906 = n4609 ^ n4562;
  assign n5909 = n5908 ^ n5907;
  assign n5910 = n5906 & n5909;
  assign n5911 = ~n5905 & n5910;
  assign n5912 = ~n5334 & ~n5911;
  assign n5914 = ~n5910 & ~n5913;
  assign n5915 = n5914 ^ n5905;
  assign n5916 = ~n5910 & ~n5915;
  assign n5917 = ~n5912 & ~n5916;
  assign n6033 = n6032 ^ n5917;
  assign n6197 = n6196 ^ n6092;
  assign n6219 = n6197 ^ n5917;
  assign n6220 = ~n6033 & n6219;
  assign n6221 = n6220 ^ n6032;
  assign n6327 = n6326 ^ n6221;
  assign n6452 = n6451 ^ n6389;
  assign n6489 = n6452 ^ n6221;
  assign n6490 = n6327 & n6489;
  assign n6491 = n6490 ^ n6326;
  assign n6558 = n6557 ^ n6491;
  assign n6487 = n6486 ^ n6483;
  assign n6466 = n6465 ^ n6461;
  assign n6480 = n6479 ^ n6466;
  assign n6488 = n6487 ^ n6480;
  assign n6565 = n6491 ^ n6488;
  assign n6566 = ~n6558 & n6565;
  assign n6567 = n6566 ^ n6557;
  assign n6585 = n6584 ^ n6567;
  assign n6601 = ~n6598 & ~n6600;
  assign n6602 = ~n6596 & n6601;
  assign n6603 = ~n6594 & n6602;
  assign n6604 = n6603 ^ n6588;
  assign n6611 = n6604 ^ n6584;
  assign n6612 = ~n6585 & n6611;
  assign n6613 = n6612 ^ n6604;
  assign n6639 = n6619 & ~n6626;
  assign n6640 = n6613 & ~n6639;
  assign n6641 = n6638 & ~n6640;
  assign n6622 = ~n6619 & ~n6621;
  assign n6627 = n6626 ^ n6622;
  assign n6628 = n6627 ^ n6613;
  assign n6605 = n6604 ^ n6585;
  assign n6559 = n6558 ^ n6488;
  assign n6453 = n6452 ^ n6327;
  assign n6199 = n4427 ^ n4425;
  assign n6200 = n5909 ^ n5906;
  assign n6201 = n6199 & n6200;
  assign n6202 = n5915 ^ n5334;
  assign n6203 = ~n6201 & ~n6202;
  assign n6204 = n4424 & n6199;
  assign n6205 = ~n6203 & ~n6204;
  assign n6206 = ~n6199 & ~n6200;
  assign n6207 = ~n4423 & n6206;
  assign n6208 = n6205 & ~n6207;
  assign n6209 = n4423 & ~n6206;
  assign n6210 = n6199 & n6202;
  assign n6211 = ~n4421 & ~n6210;
  assign n6212 = ~n6209 & n6211;
  assign n6213 = n6208 & ~n6212;
  assign n6198 = n6197 ^ n6033;
  assign n6214 = n6213 ^ n6198;
  assign n6215 = n4433 ^ n4432;
  assign n6216 = n6215 ^ n6198;
  assign n6217 = n6214 & n6216;
  assign n6218 = n6217 ^ n6213;
  assign n6454 = n6453 ^ n6218;
  assign n6455 = n4439 ^ n4438;
  assign n6456 = n6455 ^ n6218;
  assign n6457 = n6454 & n6456;
  assign n6458 = n6457 ^ n6453;
  assign n6560 = n6559 ^ n6458;
  assign n6561 = n4442 ^ n4420;
  assign n6562 = n6561 ^ n6559;
  assign n6563 = n6560 & ~n6562;
  assign n6564 = n6563 ^ n6561;
  assign n6606 = n6605 ^ n6564;
  assign n6607 = n4450 ^ n4447;
  assign n6608 = n6607 ^ n6564;
  assign n6609 = ~n6606 & n6608;
  assign n6610 = n6609 ^ n6607;
  assign n6629 = n6628 ^ n6610;
  assign n6632 = n4453 ^ n4416;
  assign n6630 = n2681 ^ n2678;
  assign n6631 = n6630 ^ n4465;
  assign n6633 = n6632 ^ n6631;
  assign n6634 = n6633 ^ n6628;
  assign n6635 = n6629 & n6634;
  assign n6636 = n6635 ^ n6610;
  assign n6642 = n6641 ^ n6636;
  assign n6643 = n2682 & ~n4463;
  assign n6644 = n4453 & ~n6630;
  assign n6645 = ~n6643 & ~n6644;
  assign n6646 = n4465 & ~n6645;
  assign n6647 = ~n1851 & ~n4465;
  assign n6648 = n1849 & ~n2675;
  assign n6649 = ~n6647 & ~n6648;
  assign n6650 = n1851 & n2635;
  assign n6651 = n2551 & n6650;
  assign n6652 = ~n6649 & ~n6651;
  assign n6653 = ~n1851 & ~n2646;
  assign n6654 = n4465 & ~n6653;
  assign n6655 = ~n1849 & n2675;
  assign n6656 = ~n6654 & ~n6655;
  assign n6657 = ~n6652 & ~n6656;
  assign n6658 = n1846 & ~n6657;
  assign n6659 = n4416 & ~n6658;
  assign n6660 = ~n2602 & ~n2642;
  assign n6661 = ~n6649 & n6656;
  assign n6662 = ~n6660 & ~n6661;
  assign n6663 = n6659 & n6662;
  assign n6664 = ~n6646 & ~n6663;
  assign n6665 = ~n4463 & ~n4465;
  assign n6666 = ~n4453 & n4471;
  assign n6667 = n6665 & ~n6666;
  assign n6668 = ~n4455 & n6667;
  assign n6669 = n6664 & ~n6668;
  assign n6670 = n6669 ^ n4460;
  assign n6671 = n6670 ^ n6636;
  assign n6672 = n6642 & ~n6671;
  assign n6673 = n6672 ^ n6670;
  assign n6674 = ~n4475 & n6673;
  assign n10136 = n6670 ^ n6642;
  assign n8137 = x659 & x660;
  assign n8138 = x657 & x658;
  assign n8139 = ~n8137 & ~n8138;
  assign n8140 = ~x659 & ~x660;
  assign n8141 = ~x657 & ~x658;
  assign n8142 = ~n8140 & ~n8141;
  assign n8143 = ~n8139 & n8142;
  assign n8144 = x656 & n8143;
  assign n8145 = n8137 & n8138;
  assign n8146 = ~n8144 & ~n8145;
  assign n8147 = n8139 & ~n8142;
  assign n8148 = ~x656 & n8147;
  assign n8149 = n8146 & ~n8148;
  assign n8150 = ~x655 & ~n8149;
  assign n8151 = ~n8145 & ~n8147;
  assign n8152 = x656 & ~n8151;
  assign n8153 = ~x656 & ~n8143;
  assign n8154 = x655 & ~n8153;
  assign n8155 = ~n8152 & n8154;
  assign n7885 = x656 ^ x655;
  assign n8156 = n8140 & n8141;
  assign n8157 = n7885 & n8156;
  assign n8158 = ~n8155 & ~n8157;
  assign n8159 = ~n8150 & n8158;
  assign n8112 = x665 & x666;
  assign n8113 = ~x663 & ~x664;
  assign n8114 = ~n8112 & n8113;
  assign n8115 = ~x665 & ~x666;
  assign n8116 = x662 & ~n8115;
  assign n8117 = n8114 & ~n8116;
  assign n8118 = x663 & x664;
  assign n8119 = n8112 & n8118;
  assign n8120 = ~n8117 & ~n8119;
  assign n8121 = n8115 & ~n8118;
  assign n8122 = ~x662 & n8121;
  assign n8123 = n8120 & ~n8122;
  assign n8124 = ~x661 & ~n8123;
  assign n8125 = ~n8114 & ~n8119;
  assign n8126 = x661 & x662;
  assign n8127 = ~n8121 & n8126;
  assign n8128 = n8125 & n8127;
  assign n7880 = x662 ^ x661;
  assign n8129 = n8112 & ~n8113;
  assign n8130 = ~n8115 & n8118;
  assign n8131 = ~n8129 & ~n8130;
  assign n8132 = n7880 & ~n8131;
  assign n8133 = ~n8128 & ~n8132;
  assign n8134 = n8113 & n8122;
  assign n8135 = n8133 & ~n8134;
  assign n8136 = ~n8124 & n8135;
  assign n8160 = n8159 ^ n8136;
  assign n7879 = x664 ^ x663;
  assign n7881 = n7880 ^ n7879;
  assign n7878 = x666 ^ x665;
  assign n7882 = n7881 ^ n7878;
  assign n7884 = x658 ^ x657;
  assign n7886 = n7885 ^ n7884;
  assign n7883 = x660 ^ x659;
  assign n7887 = n7886 ^ n7883;
  assign n8108 = n7882 & n7887;
  assign n9122 = n8136 ^ n8108;
  assign n9123 = n8160 & ~n9122;
  assign n9124 = n9123 ^ n8159;
  assign n9125 = ~n8119 & n8133;
  assign n9711 = n9124 & ~n9125;
  assign n8161 = n8160 ^ n8108;
  assign n7891 = x674 ^ x673;
  assign n7890 = x676 ^ x675;
  assign n7892 = n7891 ^ n7890;
  assign n7889 = x678 ^ x677;
  assign n7893 = n7892 ^ n7889;
  assign n7896 = x672 ^ x671;
  assign n7895 = x670 ^ x669;
  assign n7897 = n7896 ^ n7895;
  assign n7894 = x668 ^ x667;
  assign n7898 = n7897 ^ n7894;
  assign n8109 = n7893 & n7898;
  assign n8162 = n8161 ^ n8109;
  assign n7888 = n7887 ^ n7882;
  assign n7899 = n7898 ^ n7893;
  assign n8107 = n7888 & n7899;
  assign n8110 = ~n8108 & ~n8109;
  assign n8111 = n8107 & n8110;
  assign n8163 = n8162 ^ n8111;
  assign n8197 = ~x671 & ~x672;
  assign n8198 = x668 & ~n8197;
  assign n8199 = x671 & x672;
  assign n8200 = x669 & x670;
  assign n8201 = n8199 & n8200;
  assign n8202 = ~n8198 & ~n8201;
  assign n8203 = n8199 ^ x670;
  assign n8204 = n7895 & ~n8203;
  assign n8205 = n8204 ^ x669;
  assign n8206 = ~n8202 & n8205;
  assign n8207 = ~x669 & ~x670;
  assign n8208 = ~n8199 & n8207;
  assign n8209 = ~n8198 & n8208;
  assign n8210 = ~n8206 & ~n8209;
  assign n8211 = ~x667 & ~n8210;
  assign n8212 = x667 & ~n8197;
  assign n8213 = n8205 & n8212;
  assign n8214 = x667 & x668;
  assign n8215 = ~n8213 & ~n8214;
  assign n8216 = ~n8197 & ~n8200;
  assign n8217 = ~n8208 & n8216;
  assign n8218 = ~x672 & n8200;
  assign n8219 = x668 & ~n8218;
  assign n8220 = ~n8217 & n8219;
  assign n8221 = ~n8215 & ~n8220;
  assign n8222 = ~n8211 & ~n8221;
  assign n8223 = x667 & ~n8207;
  assign n8224 = ~x668 & ~x672;
  assign n8225 = ~n8200 & n8224;
  assign n8226 = ~n8223 & n8225;
  assign n8227 = n8200 & n8214;
  assign n8228 = ~n8226 & ~n8227;
  assign n8229 = ~x671 & ~n8228;
  assign n8230 = n8222 & ~n8229;
  assign n8164 = ~x677 & ~x678;
  assign n8165 = x673 & ~n8164;
  assign n8166 = x677 & x678;
  assign n8167 = n8166 ^ x676;
  assign n8168 = n7890 & ~n8167;
  assign n8169 = n8168 ^ x675;
  assign n8170 = n8165 & n8169;
  assign n8171 = x673 & x674;
  assign n8172 = ~n8170 & ~n8171;
  assign n8173 = ~x675 & ~x676;
  assign n8174 = ~n8166 & n8173;
  assign n8175 = x675 & x676;
  assign n8176 = ~n8164 & ~n8175;
  assign n8177 = ~n8174 & n8176;
  assign n8178 = ~x678 & n8175;
  assign n8179 = x674 & ~n8178;
  assign n8180 = ~n8177 & n8179;
  assign n8181 = ~n8172 & ~n8180;
  assign n8182 = x674 & ~n8164;
  assign n8183 = n8166 & n8175;
  assign n8184 = ~n8182 & ~n8183;
  assign n8185 = n8169 & ~n8184;
  assign n8186 = n8174 & ~n8182;
  assign n8187 = ~n8185 & ~n8186;
  assign n8188 = ~x673 & ~n8187;
  assign n8189 = ~n8181 & ~n8188;
  assign n8190 = ~x674 & ~x678;
  assign n8191 = ~n8175 & n8190;
  assign n8192 = n7892 & n8191;
  assign n8193 = n8171 & n8175;
  assign n8194 = ~n8192 & ~n8193;
  assign n8195 = ~x677 & ~n8194;
  assign n8196 = n8189 & ~n8195;
  assign n8231 = n8230 ^ n8196;
  assign n9136 = n8163 & ~n8231;
  assign n9137 = n8108 & n8160;
  assign n9138 = ~n8107 & n8110;
  assign n9139 = ~n8160 & n9138;
  assign n9140 = ~n9137 & ~n9139;
  assign n9141 = ~n9136 & n9140;
  assign n9142 = n8109 & n8231;
  assign n9143 = n9141 & ~n9142;
  assign n9133 = ~n8181 & ~n8185;
  assign n9132 = ~n8206 & ~n8221;
  assign n9134 = n9133 ^ n9132;
  assign n9129 = n8230 ^ n8109;
  assign n9130 = ~n8231 & n9129;
  assign n9131 = n9130 ^ n8109;
  assign n9135 = n9134 ^ n9131;
  assign n9144 = n9143 ^ n9135;
  assign n9127 = n8146 & ~n8155;
  assign n9712 = n9135 ^ n9127;
  assign n9713 = n9144 & n9712;
  assign n9714 = n9713 ^ n9143;
  assign n9715 = n9711 & ~n9714;
  assign n9716 = ~n9135 & ~n9143;
  assign n9126 = n9125 ^ n9124;
  assign n9717 = ~n9126 & n9127;
  assign n9718 = ~n9716 & n9717;
  assign n9719 = ~n9715 & ~n9718;
  assign n9720 = ~n9124 & n9125;
  assign n9721 = n9714 & n9720;
  assign n9722 = n9135 & n9143;
  assign n9723 = ~n9126 & ~n9127;
  assign n9724 = ~n9722 & n9723;
  assign n9725 = ~n9721 & ~n9724;
  assign n9726 = n9719 & n9725;
  assign n9708 = n9133 ^ n9131;
  assign n9709 = ~n9134 & ~n9708;
  assign n9710 = n9709 ^ n9131;
  assign n9727 = n9726 ^ n9710;
  assign n9947 = ~n9711 & ~n9727;
  assign n9948 = ~n9710 & ~n9714;
  assign n9949 = ~n9947 & ~n9948;
  assign n8069 = x695 & x696;
  assign n8070 = x693 & x694;
  assign n8071 = n8069 & n8070;
  assign n8072 = ~x695 & ~x696;
  assign n8073 = x692 & ~n8072;
  assign n8074 = ~n8071 & ~n8073;
  assign n7919 = x694 ^ x693;
  assign n8075 = n8069 ^ x694;
  assign n8076 = n7919 & ~n8075;
  assign n8077 = n8076 ^ x693;
  assign n8078 = ~n8074 & n8077;
  assign n8087 = x691 & ~n8072;
  assign n8088 = n8077 & n8087;
  assign n8089 = x691 & x692;
  assign n8090 = ~n8088 & ~n8089;
  assign n8079 = ~x693 & ~x694;
  assign n8080 = ~n8069 & n8079;
  assign n8091 = ~n8070 & ~n8072;
  assign n8092 = ~n8080 & n8091;
  assign n8093 = ~x696 & n8070;
  assign n8094 = x692 & ~n8093;
  assign n8095 = ~n8092 & n8094;
  assign n8096 = ~n8090 & ~n8095;
  assign n9161 = ~n8078 & ~n8096;
  assign n8039 = ~x699 & ~x700;
  assign n8040 = ~x701 & ~x702;
  assign n8041 = ~n8039 & ~n8040;
  assign n8042 = x699 & x700;
  assign n8043 = x701 & x702;
  assign n8044 = ~n8042 & ~n8043;
  assign n8045 = n8041 & ~n8044;
  assign n8046 = x698 & n8045;
  assign n8047 = n8042 & n8043;
  assign n8048 = ~n8046 & ~n8047;
  assign n8055 = ~x698 & n8045;
  assign n8049 = ~n8041 & n8044;
  assign n8056 = x702 & n8042;
  assign n8057 = x698 & ~n8056;
  assign n8058 = ~n8049 & n8057;
  assign n8059 = ~n8055 & ~n8058;
  assign n8060 = x697 & ~n8059;
  assign n9160 = n8048 & ~n8060;
  assign n9162 = n9161 ^ n9160;
  assign n8081 = ~n8073 & n8080;
  assign n8082 = ~x692 & ~n8070;
  assign n8083 = n8072 & n8082;
  assign n8084 = ~n8081 & ~n8083;
  assign n8085 = ~n8078 & n8084;
  assign n8086 = ~x691 & ~n8085;
  assign n8097 = ~n8086 & ~n8096;
  assign n8098 = n8070 & n8089;
  assign n8099 = ~x692 & ~x696;
  assign n8100 = n8079 & n8099;
  assign n8101 = ~n8098 & ~n8100;
  assign n8102 = ~x695 & ~n8101;
  assign n8103 = n8097 & ~n8102;
  assign n8050 = ~x698 & n8049;
  assign n8051 = n8039 & n8040;
  assign n8052 = ~n8050 & ~n8051;
  assign n8053 = n8048 & n8052;
  assign n8054 = ~x697 & ~n8053;
  assign n8061 = x697 & x698;
  assign n8062 = n8042 & n8061;
  assign n8063 = ~x698 & ~x702;
  assign n8064 = n8039 & n8063;
  assign n8065 = ~n8062 & ~n8064;
  assign n8066 = ~x701 & ~n8065;
  assign n8067 = ~n8060 & ~n8066;
  assign n8068 = ~n8054 & n8067;
  assign n8104 = n8103 ^ n8068;
  assign n7914 = x700 ^ x699;
  assign n7913 = x702 ^ x701;
  assign n7915 = n7914 ^ n7913;
  assign n7912 = x698 ^ x697;
  assign n7916 = n7915 ^ n7912;
  assign n7918 = x696 ^ x695;
  assign n7920 = n7919 ^ n7918;
  assign n7917 = x692 ^ x691;
  assign n7921 = n7920 ^ n7917;
  assign n8038 = n7916 & n7921;
  assign n9157 = n8068 ^ n8038;
  assign n9158 = n8104 & ~n9157;
  assign n9159 = n9158 ^ n8103;
  assign n9163 = n9162 ^ n9159;
  assign n7985 = x687 & x688;
  assign n7986 = ~x689 & ~x690;
  assign n7987 = ~n7985 & n7986;
  assign n7988 = x685 & ~n7987;
  assign n7989 = x689 & x690;
  assign n7990 = ~x687 & ~x688;
  assign n7991 = ~n7989 & n7990;
  assign n7992 = n7985 & n7989;
  assign n7993 = ~n7991 & ~n7992;
  assign n7994 = n7988 & n7993;
  assign n7995 = x685 & ~x686;
  assign n7996 = ~n7994 & ~n7995;
  assign n7907 = x688 ^ x687;
  assign n7997 = n7989 ^ x688;
  assign n7998 = n7907 & ~n7997;
  assign n7999 = n7998 ^ x687;
  assign n8000 = ~n7986 & n7999;
  assign n8001 = ~x686 & ~n8000;
  assign n8002 = ~n7996 & ~n8001;
  assign n8003 = x686 & ~n7986;
  assign n8004 = ~n7992 & ~n8003;
  assign n8005 = n7999 & ~n8004;
  assign n8006 = n7991 & ~n8003;
  assign n8007 = ~n8005 & ~n8006;
  assign n8008 = ~x685 & ~n8007;
  assign n8009 = ~n8002 & ~n8008;
  assign n7908 = x690 ^ x689;
  assign n7909 = n7908 ^ n7907;
  assign n7906 = x686 ^ x685;
  assign n7910 = n7909 ^ n7906;
  assign n8010 = ~x686 & n7987;
  assign n8011 = n7910 & n8010;
  assign n8012 = n8009 & ~n8011;
  assign n8013 = x681 & x682;
  assign n8014 = x683 & x684;
  assign n8015 = ~n8013 & ~n8014;
  assign n8016 = ~x681 & ~x682;
  assign n8017 = ~x683 & ~x684;
  assign n8018 = ~n8016 & ~n8017;
  assign n8019 = ~n8015 & n8018;
  assign n8020 = x680 & n8019;
  assign n8021 = n8013 & n8014;
  assign n8022 = ~n8020 & ~n8021;
  assign n8023 = n8015 & ~n8018;
  assign n8024 = ~x680 & n8023;
  assign n8025 = n8022 & ~n8024;
  assign n8026 = ~x679 & ~n8025;
  assign n8027 = ~n8021 & ~n8023;
  assign n8028 = x680 & ~n8027;
  assign n8029 = ~x680 & ~n8019;
  assign n8030 = x679 & ~n8029;
  assign n8031 = ~n8028 & n8030;
  assign n7903 = x680 ^ x679;
  assign n8032 = n8016 & n8017;
  assign n8033 = n7903 & n8032;
  assign n8034 = ~n8031 & ~n8033;
  assign n8035 = ~n8026 & n8034;
  assign n9155 = n8012 & n8035;
  assign n9153 = ~n8002 & ~n8005;
  assign n9152 = n8022 & ~n8031;
  assign n9154 = n9153 ^ n9152;
  assign n9156 = n9155 ^ n9154;
  assign n9164 = n9163 ^ n9156;
  assign n8036 = n8035 ^ n8012;
  assign n7922 = n7921 ^ n7916;
  assign n7981 = n7922 ^ n7910;
  assign n7902 = x684 ^ x683;
  assign n7904 = n7903 ^ n7902;
  assign n7901 = x682 ^ x681;
  assign n7905 = n7904 ^ n7901;
  assign n7982 = n7922 ^ n7905;
  assign n7983 = n7981 & ~n7982;
  assign n7984 = n7983 ^ n7910;
  assign n8037 = n8036 ^ n7984;
  assign n8105 = n8104 ^ n8038;
  assign n9149 = n8105 ^ n8036;
  assign n9150 = ~n8037 & n9149;
  assign n9151 = n9150 ^ n8105;
  assign n9165 = n9164 ^ n9151;
  assign n9691 = ~n9152 & ~n9153;
  assign n9692 = ~n9165 & n9691;
  assign n9693 = n9154 & n9155;
  assign n9694 = n9151 & n9693;
  assign n9695 = ~n9692 & ~n9694;
  assign n9696 = n9163 & ~n9695;
  assign n9688 = n9161 ^ n9159;
  assign n9689 = ~n9162 & ~n9688;
  assign n9690 = n9689 ^ n9159;
  assign n9697 = ~n9151 & n9164;
  assign n9698 = n9153 & ~n9693;
  assign n9699 = n9697 & n9698;
  assign n9700 = n9152 & ~n9155;
  assign n9701 = ~n9163 & n9700;
  assign n9702 = ~n9699 & ~n9701;
  assign n9703 = n9151 & ~n9153;
  assign n9704 = ~n9702 & ~n9703;
  assign n9705 = ~n9696 & ~n9704;
  assign n9945 = n9690 & n9705;
  assign n9946 = ~n9696 & ~n9945;
  assign n9950 = n9949 ^ n9946;
  assign n9706 = n9705 ^ n9690;
  assign n8232 = n8231 ^ n8163;
  assign n8106 = n8105 ^ n8037;
  assign n8233 = n8232 ^ n8106;
  assign n7900 = n7899 ^ n7888;
  assign n7911 = n7910 ^ n7905;
  assign n7923 = n7922 ^ n7911;
  assign n7978 = n7900 & n7923;
  assign n9146 = n8106 ^ n7978;
  assign n9147 = n8233 & ~n9146;
  assign n9148 = n9147 ^ n8232;
  assign n9166 = n9165 ^ n9148;
  assign n9128 = n9127 ^ n9126;
  assign n9145 = n9144 ^ n9128;
  assign n9685 = n9148 ^ n9145;
  assign n9686 = n9166 & ~n9685;
  assign n9687 = n9686 ^ n9165;
  assign n9707 = n9706 ^ n9687;
  assign n9942 = n9727 ^ n9706;
  assign n9943 = ~n9707 & ~n9942;
  assign n9944 = n9943 ^ n9727;
  assign n9951 = n9950 ^ n9944;
  assign n8406 = x731 & x732;
  assign n8407 = x729 & x730;
  assign n8408 = ~n8406 & ~n8407;
  assign n8409 = x728 & ~n8408;
  assign n8410 = ~x731 & ~x732;
  assign n8411 = ~x729 & ~x730;
  assign n8412 = ~n8410 & ~n8411;
  assign n8413 = n8409 & n8412;
  assign n8414 = n8406 & n8407;
  assign n8415 = ~n8413 & ~n8414;
  assign n8416 = n8408 & ~n8412;
  assign n7966 = x732 ^ x731;
  assign n7965 = x730 ^ x729;
  assign n7967 = n7966 ^ n7965;
  assign n7964 = x728 ^ x727;
  assign n7968 = n7967 ^ n7964;
  assign n8421 = x727 & ~n7968;
  assign n8423 = ~n8416 & n8421;
  assign n9207 = n8415 & ~n8423;
  assign n7955 = x746 ^ x745;
  assign n7954 = x748 ^ x747;
  assign n8458 = x749 & x750;
  assign n8459 = n8458 ^ x748;
  assign n8460 = n7954 & ~n8459;
  assign n8461 = n8460 ^ x747;
  assign n8462 = n7955 & n8461;
  assign n8463 = ~x747 & ~x748;
  assign n8464 = ~n8458 & n8463;
  assign n8465 = x747 & x748;
  assign n8466 = x745 & x746;
  assign n8467 = ~n8465 & n8466;
  assign n8468 = ~n8464 & n8467;
  assign n8469 = ~n8462 & ~n8468;
  assign n8470 = ~x749 & ~x750;
  assign n8471 = ~n8469 & ~n8470;
  assign n8472 = n8465 & n8466;
  assign n8473 = ~x750 & n8472;
  assign n8474 = ~n8471 & ~n8473;
  assign n8475 = x746 & ~n8470;
  assign n8476 = n8458 & n8465;
  assign n8477 = ~n8475 & ~n8476;
  assign n8478 = n8461 & ~n8477;
  assign n9212 = n8474 & ~n8478;
  assign n8428 = ~x741 & ~x742;
  assign n8429 = ~x743 & ~x744;
  assign n8430 = ~n8428 & ~n8429;
  assign n8431 = x741 & x742;
  assign n8432 = x743 & x744;
  assign n8433 = ~n8431 & ~n8432;
  assign n8434 = n8430 & ~n8433;
  assign n8435 = x740 & n8434;
  assign n8436 = n8431 & n8432;
  assign n8437 = ~n8435 & ~n8436;
  assign n8444 = ~x740 & n8434;
  assign n8438 = ~n8430 & n8433;
  assign n8445 = x744 & n8431;
  assign n8446 = x740 & ~n8445;
  assign n8447 = ~n8438 & n8446;
  assign n8448 = ~n8444 & ~n8447;
  assign n8449 = x739 & ~n8448;
  assign n9211 = n8437 & ~n8449;
  assign n9213 = n9212 ^ n9211;
  assign n8479 = n8464 & ~n8475;
  assign n8480 = ~x746 & ~n8465;
  assign n8481 = n8470 & n8480;
  assign n8482 = ~n8479 & ~n8481;
  assign n8483 = ~n8478 & n8482;
  assign n8484 = ~x745 & ~n8483;
  assign n8485 = n8474 & ~n8484;
  assign n8486 = ~x746 & ~x750;
  assign n8487 = n8463 & n8486;
  assign n8488 = ~n8472 & ~n8487;
  assign n8489 = ~x749 & ~n8488;
  assign n8490 = n8485 & ~n8489;
  assign n8439 = ~x740 & n8438;
  assign n8440 = n8428 & n8429;
  assign n8441 = ~n8439 & ~n8440;
  assign n8442 = n8437 & n8441;
  assign n8443 = ~x739 & ~n8442;
  assign n8450 = x739 & x740;
  assign n8451 = n8431 & n8450;
  assign n8452 = ~x740 & ~x744;
  assign n8453 = n8428 & n8452;
  assign n8454 = ~n8451 & ~n8453;
  assign n8455 = ~x743 & ~n8454;
  assign n8456 = ~n8449 & ~n8455;
  assign n8457 = ~n8443 & n8456;
  assign n8491 = n8490 ^ n8457;
  assign n7950 = x742 ^ x741;
  assign n7949 = x744 ^ x743;
  assign n7951 = n7950 ^ n7949;
  assign n7948 = x740 ^ x739;
  assign n7952 = n7951 ^ n7948;
  assign n7956 = n7955 ^ n7954;
  assign n7953 = x750 ^ x749;
  assign n7957 = n7956 ^ n7953;
  assign n8368 = n7952 & n7957;
  assign n9208 = n8457 ^ n8368;
  assign n9209 = n8491 & ~n9208;
  assign n9210 = n9209 ^ n8490;
  assign n9214 = n9213 ^ n9210;
  assign n9735 = n9207 & ~n9214;
  assign n7961 = x734 ^ x733;
  assign n7960 = x736 ^ x735;
  assign n7962 = n7961 ^ n7960;
  assign n7959 = x738 ^ x737;
  assign n7963 = n7962 ^ n7959;
  assign n8372 = n7963 & n7968;
  assign n8417 = ~x728 & n8416;
  assign n8418 = n8410 & n8411;
  assign n8419 = ~n8417 & ~n8418;
  assign n8420 = n8415 & n8419;
  assign n8422 = ~n8420 & ~n8421;
  assign n8424 = ~n8414 & n8423;
  assign n8425 = ~n8422 & ~n8424;
  assign n8376 = x737 & x738;
  assign n8377 = x735 & x736;
  assign n8378 = ~n8376 & ~n8377;
  assign n8379 = ~x737 & ~x738;
  assign n8380 = ~x735 & ~x736;
  assign n8381 = ~n8379 & ~n8380;
  assign n8382 = ~n8378 & n8381;
  assign n8383 = x734 & n8382;
  assign n8384 = n8376 & n8377;
  assign n8385 = ~n8383 & ~n8384;
  assign n8386 = x734 & ~n8379;
  assign n8387 = ~n8376 & n8380;
  assign n8388 = ~n8386 & n8387;
  assign n8389 = n8385 & ~n8388;
  assign n8390 = ~x733 & ~n8389;
  assign n8391 = ~x734 & n8379;
  assign n8392 = ~n8377 & n8391;
  assign n8393 = n7962 & n8392;
  assign n8394 = x733 & x734;
  assign n8395 = ~x737 & n8394;
  assign n8396 = n8377 & n8395;
  assign n8397 = ~n8393 & ~n8396;
  assign n8398 = n7961 & n8382;
  assign n8399 = n8378 & ~n8381;
  assign n8400 = x738 & n8377;
  assign n8401 = n8394 & ~n8400;
  assign n8402 = ~n8399 & n8401;
  assign n8403 = ~n8398 & ~n8402;
  assign n8404 = n8397 & n8403;
  assign n8405 = ~n8390 & n8404;
  assign n8426 = n8425 ^ n8405;
  assign n9197 = ~n8372 & n8426;
  assign n9198 = ~n8405 & ~n8425;
  assign n9199 = ~n9197 & ~n9198;
  assign n9196 = n8385 & n8403;
  assign n9200 = n9199 ^ n9196;
  assign n7969 = n7968 ^ n7963;
  assign n7958 = n7957 ^ n7952;
  assign n8369 = n7963 ^ n7958;
  assign n8370 = n7969 & ~n8369;
  assign n8371 = n8370 ^ n7968;
  assign n8373 = n8372 ^ n8371;
  assign n8374 = ~n8368 & ~n8373;
  assign n8375 = n8374 ^ n8372;
  assign n8427 = n8426 ^ n8375;
  assign n8492 = n8491 ^ n8427;
  assign n9201 = ~n8368 & n8491;
  assign n9202 = ~n8492 & ~n9201;
  assign n9203 = ~n8373 & ~n8426;
  assign n9204 = n9203 ^ n8372;
  assign n9205 = ~n9202 & ~n9204;
  assign n9736 = n9205 ^ n9199;
  assign n9737 = n9200 & n9736;
  assign n9738 = n9737 ^ n9205;
  assign n9739 = n9735 & ~n9738;
  assign n9215 = n9214 ^ n9207;
  assign n9740 = n9196 & ~n9199;
  assign n9741 = ~n9205 & n9740;
  assign n9742 = ~n9215 & n9741;
  assign n9743 = ~n9739 & ~n9742;
  assign n9732 = n9212 ^ n9210;
  assign n9733 = ~n9213 & ~n9732;
  assign n9734 = n9733 ^ n9210;
  assign n9206 = n9205 ^ n9200;
  assign n9216 = n9215 ^ n9206;
  assign n9744 = n9214 & n9738;
  assign n9745 = ~n9216 & n9744;
  assign n9938 = ~n9734 & ~n9745;
  assign n9939 = n9743 & ~n9938;
  assign n8335 = x705 & x706;
  assign n8336 = x707 & x708;
  assign n8337 = ~n8335 & ~n8336;
  assign n8338 = ~x705 & ~x706;
  assign n8339 = ~x707 & ~x708;
  assign n8340 = ~n8338 & ~n8339;
  assign n8341 = ~n8337 & n8340;
  assign n8342 = x704 & n8341;
  assign n8343 = n8335 & n8336;
  assign n8344 = ~n8342 & ~n8343;
  assign n8357 = n8337 & ~n8340;
  assign n8353 = x703 & x704;
  assign n8354 = n8335 & n8353;
  assign n8358 = x708 & n8354;
  assign n8359 = n8358 ^ n8353;
  assign n8360 = ~n8357 & n8359;
  assign n7943 = x704 ^ x703;
  assign n8361 = n7943 & n8341;
  assign n8362 = ~n8360 & ~n8361;
  assign n9175 = n8344 & n8362;
  assign n8305 = x711 & x712;
  assign n8306 = x713 & x714;
  assign n8307 = ~n8305 & ~n8306;
  assign n8308 = ~x711 & ~x712;
  assign n8309 = ~x713 & ~x714;
  assign n8310 = ~n8308 & ~n8309;
  assign n8311 = ~n8307 & n8310;
  assign n8312 = x710 & n8311;
  assign n8313 = n8305 & n8306;
  assign n8314 = ~n8312 & ~n8313;
  assign n8327 = n8307 & ~n8310;
  assign n8323 = x709 & x710;
  assign n8324 = n8305 & n8323;
  assign n8328 = x714 & n8324;
  assign n8329 = n8328 ^ n8323;
  assign n8330 = ~n8327 & n8329;
  assign n7938 = x710 ^ x709;
  assign n8331 = n7938 & n8311;
  assign n8332 = ~n8330 & ~n8331;
  assign n9174 = n8314 & n8332;
  assign n9176 = n9175 ^ n9174;
  assign n8345 = x704 & ~n8339;
  assign n8346 = ~n8336 & n8338;
  assign n8347 = ~n8345 & n8346;
  assign n8348 = n8344 & ~n8347;
  assign n8349 = ~x703 & ~n8348;
  assign n7942 = x706 ^ x705;
  assign n7944 = n7943 ^ n7942;
  assign n8350 = ~x704 & ~x708;
  assign n8351 = ~n8335 & n8350;
  assign n8352 = n7944 & n8351;
  assign n8355 = ~n8352 & ~n8354;
  assign n8356 = ~x707 & ~n8355;
  assign n8363 = ~n8356 & n8362;
  assign n8364 = ~n8349 & n8363;
  assign n8315 = x710 & ~n8309;
  assign n8316 = ~n8306 & n8308;
  assign n8317 = ~n8315 & n8316;
  assign n8318 = n8314 & ~n8317;
  assign n8319 = ~x709 & ~n8318;
  assign n7937 = x712 ^ x711;
  assign n7939 = n7938 ^ n7937;
  assign n8320 = ~x710 & ~x714;
  assign n8321 = ~n8305 & n8320;
  assign n8322 = n7939 & n8321;
  assign n8325 = ~n8322 & ~n8324;
  assign n8326 = ~x713 & ~n8325;
  assign n8333 = ~n8326 & n8332;
  assign n8334 = ~n8319 & n8333;
  assign n8365 = n8364 ^ n8334;
  assign n7936 = x714 ^ x713;
  assign n7940 = n7939 ^ n7936;
  assign n7941 = x708 ^ x707;
  assign n7945 = n7944 ^ n7941;
  assign n8237 = n7940 & n7945;
  assign n9171 = n8364 ^ n8237;
  assign n9172 = ~n8365 & n9171;
  assign n9173 = n9172 ^ n8237;
  assign n9177 = n9176 ^ n9173;
  assign n8271 = x723 & x724;
  assign n8272 = x725 & x726;
  assign n8273 = ~n8271 & ~n8272;
  assign n8274 = ~x723 & ~x724;
  assign n8275 = ~x725 & ~x726;
  assign n8276 = ~n8274 & ~n8275;
  assign n8277 = ~n8273 & n8276;
  assign n8278 = x722 & n8277;
  assign n8279 = n8271 & n8272;
  assign n8280 = ~n8278 & ~n8279;
  assign n8281 = x722 & ~n8275;
  assign n8282 = ~n8272 & n8274;
  assign n8283 = ~n8281 & n8282;
  assign n8284 = n8280 & ~n8283;
  assign n8285 = ~x721 & ~n8284;
  assign n7932 = x722 ^ x721;
  assign n7931 = x724 ^ x723;
  assign n7933 = n7932 ^ n7931;
  assign n8286 = ~x722 & ~x726;
  assign n8287 = ~n8271 & n8286;
  assign n8288 = n7933 & n8287;
  assign n8289 = x721 & x722;
  assign n8290 = n8271 & n8289;
  assign n8291 = ~n8288 & ~n8290;
  assign n8292 = ~x725 & ~n8291;
  assign n8293 = n8273 & ~n8276;
  assign n8294 = x726 & n8290;
  assign n8295 = n8294 ^ n8289;
  assign n8296 = ~n8293 & n8295;
  assign n8297 = n7932 & n8277;
  assign n8298 = ~n8296 & ~n8297;
  assign n8299 = ~n8292 & n8298;
  assign n8300 = ~n8285 & n8299;
  assign n8241 = x717 & x718;
  assign n8242 = x719 & x720;
  assign n8243 = ~n8241 & ~n8242;
  assign n8244 = ~x717 & ~x718;
  assign n8245 = ~x719 & ~x720;
  assign n8246 = ~n8244 & ~n8245;
  assign n8247 = ~n8243 & n8246;
  assign n8248 = x716 & n8247;
  assign n8249 = n8241 & n8242;
  assign n8250 = ~n8248 & ~n8249;
  assign n8251 = x716 & ~n8245;
  assign n8252 = ~n8242 & n8244;
  assign n8253 = ~n8251 & n8252;
  assign n8254 = n8250 & ~n8253;
  assign n8255 = ~x715 & ~n8254;
  assign n7927 = x716 ^ x715;
  assign n7926 = x718 ^ x717;
  assign n7928 = n7927 ^ n7926;
  assign n8256 = ~x716 & ~x720;
  assign n8257 = ~n8241 & n8256;
  assign n8258 = n7928 & n8257;
  assign n8259 = x715 & x716;
  assign n8260 = n8241 & n8259;
  assign n8261 = ~n8258 & ~n8260;
  assign n8262 = ~x719 & ~n8261;
  assign n8263 = n8243 & ~n8246;
  assign n8264 = x720 & n8260;
  assign n8265 = n8264 ^ n8259;
  assign n8266 = ~n8263 & n8265;
  assign n8267 = n7927 & n8247;
  assign n8268 = ~n8266 & ~n8267;
  assign n8269 = ~n8262 & n8268;
  assign n8270 = ~n8255 & n8269;
  assign n8301 = n8300 ^ n8270;
  assign n8302 = n8301 ^ n8237;
  assign n7925 = x720 ^ x719;
  assign n7929 = n7928 ^ n7925;
  assign n7930 = x726 ^ x725;
  assign n7934 = n7933 ^ n7930;
  assign n8238 = n7929 & n7934;
  assign n8303 = n8302 ^ n8238;
  assign n7935 = n7934 ^ n7929;
  assign n7946 = n7945 ^ n7940;
  assign n8236 = n7935 & n7946;
  assign n8239 = ~n8237 & ~n8238;
  assign n8240 = n8236 & n8239;
  assign n8304 = n8303 ^ n8240;
  assign n9185 = n8304 & ~n8365;
  assign n9186 = ~n8236 & n8239;
  assign n9187 = n9186 ^ n8238;
  assign n9188 = ~n8301 & n9187;
  assign n9189 = n9188 ^ n8238;
  assign n9190 = ~n9185 & ~n9189;
  assign n9191 = n8237 & n8365;
  assign n9192 = n9190 & ~n9191;
  assign n9181 = n8238 & n8301;
  assign n9182 = n8270 & n8300;
  assign n9183 = ~n9181 & ~n9182;
  assign n9179 = n8280 & n8298;
  assign n9178 = n8250 & n8268;
  assign n9180 = n9179 ^ n9178;
  assign n9184 = n9183 ^ n9180;
  assign n9193 = n9192 ^ n9184;
  assign n9754 = n9177 & ~n9193;
  assign n9755 = ~n9184 & n9192;
  assign n9756 = n9175 ^ n9173;
  assign n9757 = ~n9176 & ~n9756;
  assign n9758 = n9757 ^ n9173;
  assign n9759 = ~n9755 & ~n9758;
  assign n9760 = ~n9754 & n9759;
  assign n9751 = n9183 ^ n9179;
  assign n9752 = ~n9180 & n9751;
  assign n9753 = n9752 ^ n9183;
  assign n9194 = n9193 ^ n9177;
  assign n9761 = ~n9184 & n9758;
  assign n9762 = n9194 & n9761;
  assign n9763 = ~n9760 & ~n9762;
  assign n9936 = n9753 & n9763;
  assign n9937 = ~n9760 & ~n9936;
  assign n9940 = n9939 ^ n9937;
  assign n9764 = n9763 ^ n9753;
  assign n8366 = n8365 ^ n8304;
  assign n7947 = n7946 ^ n7935;
  assign n7970 = n7969 ^ n7958;
  assign n8235 = n7947 & n7970;
  assign n8367 = n8366 ^ n8235;
  assign n9168 = n8492 ^ n8235;
  assign n9169 = n8367 & n9168;
  assign n9170 = n9169 ^ n8366;
  assign n9195 = n9194 ^ n9170;
  assign n9748 = n9216 ^ n9170;
  assign n9749 = ~n9195 & ~n9748;
  assign n9750 = n9749 ^ n9194;
  assign n9765 = n9764 ^ n9750;
  assign n9746 = n9743 & ~n9745;
  assign n9747 = n9746 ^ n9734;
  assign n9933 = n9750 ^ n9747;
  assign n9934 = n9765 & n9933;
  assign n9935 = n9934 ^ n9764;
  assign n9941 = n9940 ^ n9935;
  assign n9952 = n9951 ^ n9941;
  assign n9766 = n9765 ^ n9747;
  assign n9217 = n9216 ^ n9195;
  assign n9167 = n9166 ^ n9145;
  assign n9218 = n9217 ^ n9167;
  assign n8493 = n8492 ^ n8367;
  assign n7924 = n7923 ^ n7900;
  assign n7971 = n7970 ^ n7947;
  assign n7979 = n7924 & n7971;
  assign n9116 = n7979 & n8233;
  assign n9117 = n8493 & ~n9116;
  assign n9118 = n7978 & n8233;
  assign n7980 = ~n7978 & ~n7979;
  assign n9119 = n7980 & ~n8233;
  assign n9120 = ~n9118 & ~n9119;
  assign n9121 = ~n9117 & n9120;
  assign n9729 = n9167 ^ n9121;
  assign n9730 = ~n9218 & ~n9729;
  assign n9731 = n9730 ^ n9217;
  assign n9767 = n9766 ^ n9731;
  assign n9728 = n9727 ^ n9707;
  assign n9930 = n9731 ^ n9728;
  assign n9931 = ~n9767 & ~n9930;
  assign n9932 = n9931 ^ n9766;
  assign n9985 = n9941 ^ n9932;
  assign n9986 = ~n9952 & n9985;
  assign n9987 = n9986 ^ n9951;
  assign n9991 = n9939 ^ n9935;
  assign n9992 = ~n9940 & ~n9991;
  assign n9993 = n9992 ^ n9935;
  assign n10081 = ~n9987 & n9993;
  assign n8534 = x789 & x790;
  assign n8535 = x791 & x792;
  assign n8536 = ~n8534 & ~n8535;
  assign n8537 = ~x789 & ~x790;
  assign n8538 = ~x791 & ~x792;
  assign n8539 = ~n8537 & ~n8538;
  assign n8540 = ~n8536 & n8539;
  assign n8541 = x788 & n8540;
  assign n8542 = n8534 & n8535;
  assign n8543 = ~n8541 & ~n8542;
  assign n7855 = x788 ^ x787;
  assign n8550 = n7855 & n8540;
  assign n8544 = n8536 & ~n8539;
  assign n8551 = x787 & x788;
  assign n8552 = n8534 & n8551;
  assign n8553 = x792 & n8552;
  assign n8554 = n8553 ^ n8551;
  assign n8555 = ~n8544 & n8554;
  assign n8556 = ~n8550 & ~n8555;
  assign n9041 = n8543 & n8556;
  assign n8505 = ~x795 & ~x796;
  assign n8506 = ~x797 & ~x798;
  assign n8507 = ~n8505 & ~n8506;
  assign n8508 = x795 & x796;
  assign n8509 = x797 & x798;
  assign n8510 = ~n8508 & ~n8509;
  assign n8511 = n8507 & ~n8510;
  assign n8512 = x794 & n8511;
  assign n8513 = n8508 & n8509;
  assign n8514 = ~n8512 & ~n8513;
  assign n7860 = x794 ^ x793;
  assign n8521 = n7860 & n8511;
  assign n8515 = ~n8507 & n8510;
  assign n8522 = x793 & x794;
  assign n8523 = n8508 & n8522;
  assign n8524 = x798 & n8523;
  assign n8525 = n8524 ^ n8522;
  assign n8526 = ~n8515 & n8525;
  assign n8527 = ~n8521 & ~n8526;
  assign n9040 = n8514 & n8527;
  assign n9042 = n9041 ^ n9040;
  assign n8545 = ~x788 & n8544;
  assign n8546 = n8537 & n8538;
  assign n8547 = ~n8545 & ~n8546;
  assign n8548 = n8543 & n8547;
  assign n8549 = ~x787 & ~n8548;
  assign n8557 = ~x788 & ~x792;
  assign n8558 = n8537 & n8557;
  assign n8559 = ~n8552 & ~n8558;
  assign n8560 = ~x791 & ~n8559;
  assign n8561 = n8556 & ~n8560;
  assign n8562 = ~n8549 & n8561;
  assign n8516 = ~x794 & n8515;
  assign n8517 = n8505 & n8506;
  assign n8518 = ~n8516 & ~n8517;
  assign n8519 = n8514 & n8518;
  assign n8520 = ~x793 & ~n8519;
  assign n8528 = ~x794 & ~x798;
  assign n8529 = n8505 & n8528;
  assign n8530 = ~n8523 & ~n8529;
  assign n8531 = ~x797 & ~n8530;
  assign n8532 = n8527 & ~n8531;
  assign n8533 = ~n8520 & n8532;
  assign n8563 = n8562 ^ n8533;
  assign n7854 = x790 ^ x789;
  assign n7856 = n7855 ^ n7854;
  assign n7853 = x792 ^ x791;
  assign n7857 = n7856 ^ n7853;
  assign n7859 = x796 ^ x795;
  assign n7861 = n7860 ^ n7859;
  assign n7858 = x798 ^ x797;
  assign n7862 = n7861 ^ n7858;
  assign n8504 = n7857 & n7862;
  assign n9037 = n8533 ^ n8504;
  assign n9038 = n8563 & ~n9037;
  assign n9039 = n9038 ^ n8562;
  assign n9835 = n9041 ^ n9039;
  assign n9836 = ~n9042 & ~n9835;
  assign n9837 = n9836 ^ n9039;
  assign n9043 = n9042 ^ n9039;
  assign n8594 = x779 & x780;
  assign n8595 = x777 & x778;
  assign n8596 = ~n8594 & ~n8595;
  assign n8597 = ~x779 & ~x780;
  assign n8598 = ~x777 & ~x778;
  assign n8599 = ~n8597 & ~n8598;
  assign n8600 = ~n8596 & n8599;
  assign n8601 = x776 & n8600;
  assign n8602 = n8594 & n8595;
  assign n8603 = ~n8601 & ~n8602;
  assign n8604 = n8596 & ~n8599;
  assign n8605 = ~x776 & n8604;
  assign n8606 = n8603 & ~n8605;
  assign n8607 = ~x775 & ~n8606;
  assign n8608 = ~n8602 & ~n8604;
  assign n8609 = x776 & ~n8608;
  assign n8610 = ~x776 & ~n8600;
  assign n8611 = x775 & ~n8610;
  assign n8612 = ~n8609 & n8611;
  assign n7866 = x776 ^ x775;
  assign n8613 = n8597 & n8598;
  assign n8614 = n7866 & n8613;
  assign n8615 = ~n8612 & ~n8614;
  assign n8616 = ~n8607 & n8615;
  assign n8565 = ~x785 & ~x786;
  assign n8566 = ~x783 & ~x784;
  assign n8567 = ~n8565 & ~n8566;
  assign n8568 = x785 & x786;
  assign n8569 = x783 & x784;
  assign n8570 = ~n8568 & ~n8569;
  assign n8571 = n8567 & ~n8570;
  assign n8572 = x782 & n8571;
  assign n8573 = n8568 & n8569;
  assign n8574 = ~n8572 & ~n8573;
  assign n8575 = ~n8567 & n8570;
  assign n8576 = ~x782 & n8575;
  assign n8577 = n8565 & n8566;
  assign n8578 = ~n8576 & ~n8577;
  assign n8579 = n8574 & n8578;
  assign n8580 = ~x781 & ~n8579;
  assign n7871 = x782 ^ x781;
  assign n8581 = n7871 & n8571;
  assign n8582 = x781 & x782;
  assign n8583 = n8569 & n8582;
  assign n8584 = x786 & n8583;
  assign n8585 = n8584 ^ n8582;
  assign n8586 = ~n8575 & n8585;
  assign n8587 = ~n8581 & ~n8586;
  assign n8588 = ~x782 & ~x786;
  assign n8589 = n8566 & n8588;
  assign n8590 = ~n8583 & ~n8589;
  assign n8591 = ~x785 & ~n8590;
  assign n8592 = n8587 & ~n8591;
  assign n8593 = ~n8580 & n8592;
  assign n8617 = n8616 ^ n8593;
  assign n7865 = x778 ^ x777;
  assign n7867 = n7866 ^ n7865;
  assign n7864 = x780 ^ x779;
  assign n7868 = n7867 ^ n7864;
  assign n7870 = x784 ^ x783;
  assign n7872 = n7871 ^ n7870;
  assign n7869 = x786 ^ x785;
  assign n7873 = n7872 ^ n7869;
  assign n9045 = ~n7868 & ~n7873;
  assign n8500 = n7868 & n7873;
  assign n9046 = n9045 ^ n8500;
  assign n9047 = n8617 & n9046;
  assign n9048 = n9047 ^ n9045;
  assign n9053 = ~n8500 & ~n8617;
  assign n7874 = n7873 ^ n7868;
  assign n9054 = ~n7862 & ~n7874;
  assign n9055 = ~n8563 & ~n9054;
  assign n9056 = ~n9053 & n9055;
  assign n9057 = ~n8504 & n8563;
  assign n9058 = ~n9056 & ~n9057;
  assign n9059 = n8563 & ~n9053;
  assign n7863 = n7862 ^ n7857;
  assign n7875 = n7874 ^ n7863;
  assign n9060 = ~n7857 & n7875;
  assign n9061 = ~n9059 & n9060;
  assign n9062 = ~n9058 & ~n9061;
  assign n9063 = ~n9048 & n9062;
  assign n9049 = ~n8616 & ~n9048;
  assign n9050 = ~n8500 & ~n8593;
  assign n9051 = ~n9049 & ~n9050;
  assign n9034 = n8574 & n8587;
  assign n9035 = n8603 & ~n8612;
  assign n9838 = ~n9034 & ~n9035;
  assign n9839 = n9051 & n9838;
  assign n9840 = ~n9063 & ~n9839;
  assign n9841 = n9043 & ~n9840;
  assign n9842 = ~n9051 & ~n9838;
  assign n9843 = n9841 & ~n9842;
  assign n9844 = ~n9837 & ~n9843;
  assign n9036 = n9035 ^ n9034;
  assign n9044 = n9043 ^ n9036;
  assign n9052 = n9051 ^ n9044;
  assign n9064 = n9063 ^ n9052;
  assign n9845 = n9034 & n9035;
  assign n9846 = n9064 & n9845;
  assign n9847 = ~n9844 & ~n9846;
  assign n9849 = ~n9043 & n9842;
  assign n9850 = ~n9846 & ~n9849;
  assign n9851 = ~n9063 & ~n9850;
  assign n9976 = n9847 & ~n9851;
  assign n8707 = x767 & x768;
  assign n8708 = x765 & x766;
  assign n8709 = ~n8707 & ~n8708;
  assign n8710 = ~x767 & ~x768;
  assign n8711 = ~x765 & ~x766;
  assign n8712 = ~n8710 & ~n8711;
  assign n8713 = n8709 & ~n8712;
  assign n8714 = x763 & x764;
  assign n8715 = n8708 & n8714;
  assign n8716 = x768 & n8715;
  assign n8717 = n8716 ^ n8714;
  assign n8718 = ~n8713 & n8717;
  assign n8719 = ~n8709 & n8712;
  assign n8720 = ~x764 & n8719;
  assign n8721 = ~x763 & n8720;
  assign n8722 = n8721 ^ n8719;
  assign n8723 = ~n8718 & ~n8722;
  assign n8724 = n8707 & n8708;
  assign n8725 = n8723 & ~n8724;
  assign n8726 = x764 & ~n8710;
  assign n8727 = ~n8707 & n8711;
  assign n8728 = ~n8726 & n8727;
  assign n8729 = n8725 & ~n8728;
  assign n8730 = x763 & ~n8718;
  assign n8731 = ~n8720 & n8730;
  assign n8732 = ~n8729 & ~n8731;
  assign n7832 = x764 ^ x763;
  assign n7831 = x766 ^ x765;
  assign n7833 = n7832 ^ n7831;
  assign n8733 = ~x764 & ~x768;
  assign n8734 = ~n8708 & n8733;
  assign n8735 = n7833 & n8734;
  assign n8736 = ~n8715 & ~n8735;
  assign n8737 = ~x767 & ~n8736;
  assign n8738 = ~n8732 & ~n8737;
  assign n8684 = x773 & x774;
  assign n8685 = x771 & x772;
  assign n8686 = ~n8684 & ~n8685;
  assign n8687 = ~x773 & ~x774;
  assign n8688 = ~x771 & ~x772;
  assign n8689 = ~n8687 & ~n8688;
  assign n8690 = ~n8686 & n8689;
  assign n8691 = x770 & n8690;
  assign n8692 = n8684 & n8685;
  assign n8693 = ~n8691 & ~n8692;
  assign n8694 = n8686 & ~n8689;
  assign n8695 = ~x770 & n8694;
  assign n8696 = n8693 & ~n8695;
  assign n8697 = ~x769 & ~n8696;
  assign n8698 = ~n8692 & ~n8694;
  assign n8699 = x770 & ~n8698;
  assign n8700 = ~x770 & ~n8690;
  assign n8701 = x769 & ~n8700;
  assign n8702 = ~n8699 & n8701;
  assign n7837 = x770 ^ x769;
  assign n8703 = n8687 & n8688;
  assign n8704 = n7837 & n8703;
  assign n8705 = ~n8702 & ~n8704;
  assign n8706 = ~n8697 & n8705;
  assign n8739 = n8738 ^ n8706;
  assign n7830 = x768 ^ x767;
  assign n7834 = n7833 ^ n7830;
  assign n7836 = x772 ^ x771;
  assign n7838 = n7837 ^ n7836;
  assign n7835 = x774 ^ x773;
  assign n7839 = n7838 ^ n7835;
  assign n8620 = n7834 & n7839;
  assign n9008 = n8706 ^ n8620;
  assign n9009 = n8739 & ~n9008;
  assign n9010 = n9009 ^ n8738;
  assign n9817 = n9010 ^ n8725;
  assign n9011 = n8693 & ~n8702;
  assign n9818 = n9011 ^ n9010;
  assign n9819 = ~n9817 & n9818;
  assign n9820 = n9819 ^ n8725;
  assign n9012 = n9011 ^ n8725;
  assign n9013 = n9012 ^ n9010;
  assign n8628 = x761 & x762;
  assign n8629 = x759 & x760;
  assign n8630 = ~n8628 & ~n8629;
  assign n8631 = ~x761 & ~x762;
  assign n8632 = ~x759 & ~x760;
  assign n8633 = ~n8631 & ~n8632;
  assign n8634 = ~n8630 & n8633;
  assign n8635 = x758 & n8634;
  assign n8636 = n8628 & n8629;
  assign n8637 = ~n8635 & ~n8636;
  assign n8638 = n8630 & ~n8633;
  assign n8642 = ~n8636 & ~n8638;
  assign n8643 = x758 & ~n8642;
  assign n8644 = ~x758 & ~n8634;
  assign n8645 = x757 & ~n8644;
  assign n8646 = ~n8643 & n8645;
  assign n9015 = n8637 & ~n8646;
  assign n8651 = x755 & x756;
  assign n8652 = x753 & x754;
  assign n8653 = n8651 & n8652;
  assign n8654 = ~n8651 & ~n8652;
  assign n8655 = ~x755 & ~x756;
  assign n8656 = ~x753 & ~x754;
  assign n8657 = ~n8655 & ~n8656;
  assign n8658 = ~n8654 & n8657;
  assign n8659 = ~x752 & n8658;
  assign n8660 = ~x751 & n8659;
  assign n8661 = n8660 ^ n8658;
  assign n8662 = ~n8653 & ~n8661;
  assign n8676 = n8654 & ~n8657;
  assign n8672 = x751 & x752;
  assign n8673 = n8652 & n8672;
  assign n8677 = x756 & n8673;
  assign n8678 = n8677 ^ n8672;
  assign n8679 = ~n8676 & n8678;
  assign n9014 = n8662 & ~n8679;
  assign n9016 = n9015 ^ n9014;
  assign n8663 = x752 & ~n8655;
  assign n8664 = ~n8651 & n8656;
  assign n8665 = ~n8663 & n8664;
  assign n8666 = n8662 & ~n8665;
  assign n8667 = x751 & ~n8659;
  assign n8668 = ~n8666 & ~n8667;
  assign n7843 = x752 ^ x751;
  assign n7842 = x754 ^ x753;
  assign n7844 = n7843 ^ n7842;
  assign n8669 = ~x752 & ~x756;
  assign n8670 = ~n8652 & n8669;
  assign n8671 = n7844 & n8670;
  assign n8674 = ~n8671 & ~n8673;
  assign n8675 = ~x755 & ~n8674;
  assign n8680 = ~n8675 & ~n8679;
  assign n8681 = ~n8668 & n8680;
  assign n8639 = ~x758 & n8638;
  assign n8640 = n8637 & ~n8639;
  assign n8641 = ~x757 & ~n8640;
  assign n7848 = x758 ^ x757;
  assign n8647 = n8631 & n8632;
  assign n8648 = n7848 & n8647;
  assign n8649 = ~n8646 & ~n8648;
  assign n8650 = ~n8641 & n8649;
  assign n8682 = n8681 ^ n8650;
  assign n7841 = x756 ^ x755;
  assign n7845 = n7844 ^ n7841;
  assign n7847 = x760 ^ x759;
  assign n7849 = n7848 ^ n7847;
  assign n7846 = x762 ^ x761;
  assign n7850 = n7849 ^ n7846;
  assign n8624 = n7845 & n7850;
  assign n7851 = n7850 ^ n7845;
  assign n7840 = n7839 ^ n7834;
  assign n8621 = n7845 ^ n7840;
  assign n8622 = n7851 & ~n8621;
  assign n8623 = n8622 ^ n7850;
  assign n8625 = n8624 ^ n8623;
  assign n8626 = ~n8620 & ~n8625;
  assign n8627 = n8626 ^ n8624;
  assign n8683 = n8682 ^ n8627;
  assign n8740 = n8739 ^ n8683;
  assign n9021 = ~n8620 & n8739;
  assign n9022 = ~n8740 & ~n9021;
  assign n9023 = ~n8625 & ~n8682;
  assign n9024 = n9023 ^ n8624;
  assign n9025 = ~n9022 & ~n9024;
  assign n9018 = ~n8624 & n8682;
  assign n9019 = ~n8650 & ~n8681;
  assign n9020 = ~n9018 & ~n9019;
  assign n9026 = n9025 ^ n9020;
  assign n9821 = n9016 & n9026;
  assign n9822 = n9013 & ~n9821;
  assign n9824 = ~n9020 & ~n9025;
  assign n9823 = n9014 & n9015;
  assign n9825 = n9824 ^ n9823;
  assign n9826 = n9822 & ~n9825;
  assign n9827 = ~n9823 & ~n9824;
  assign n9828 = n9020 & n9025;
  assign n9829 = ~n9014 & ~n9015;
  assign n9830 = ~n9013 & ~n9829;
  assign n9831 = ~n9828 & n9830;
  assign n9832 = ~n9827 & n9831;
  assign n9833 = ~n9826 & ~n9832;
  assign n9973 = ~n9820 & n9833;
  assign n9974 = n9822 & n9827;
  assign n9975 = ~n9973 & ~n9974;
  assign n9977 = n9976 ^ n9975;
  assign n8900 = x813 & x814;
  assign n8901 = x815 & x816;
  assign n8902 = ~n8900 & ~n8901;
  assign n8903 = ~x813 & ~x814;
  assign n8904 = ~x815 & ~x816;
  assign n8905 = ~n8903 & ~n8904;
  assign n8906 = ~n8902 & n8905;
  assign n8907 = x812 & n8906;
  assign n8908 = n8900 & n8901;
  assign n8909 = ~n8907 & ~n8908;
  assign n8910 = x812 & ~n8904;
  assign n8911 = ~n8901 & n8903;
  assign n8912 = ~n8910 & n8911;
  assign n8913 = n8909 & ~n8912;
  assign n8914 = ~x811 & ~n8913;
  assign n8915 = x811 & ~n8903;
  assign n8916 = ~x812 & ~x816;
  assign n8917 = ~n8900 & n8916;
  assign n8918 = ~n8915 & n8917;
  assign n8919 = x811 & x812;
  assign n8920 = n8900 & n8919;
  assign n8921 = ~n8918 & ~n8920;
  assign n8922 = ~x815 & ~n8921;
  assign n7801 = x812 ^ x811;
  assign n8923 = n7801 & n8906;
  assign n8924 = n8902 & ~n8905;
  assign n8925 = x816 & n8920;
  assign n8926 = n8925 ^ n8919;
  assign n8927 = ~n8924 & n8926;
  assign n8928 = ~n8923 & ~n8927;
  assign n8929 = ~n8922 & n8928;
  assign n8930 = ~n8914 & n8929;
  assign n8869 = x819 & x820;
  assign n8870 = x821 & x822;
  assign n8871 = ~n8869 & ~n8870;
  assign n8872 = ~x819 & ~x820;
  assign n8873 = ~x821 & ~x822;
  assign n8874 = ~n8872 & ~n8873;
  assign n8875 = ~n8871 & n8874;
  assign n8876 = x818 & n8875;
  assign n8877 = n8869 & n8870;
  assign n8878 = ~n8876 & ~n8877;
  assign n8879 = x818 & ~n8873;
  assign n8880 = ~n8870 & n8872;
  assign n8881 = ~n8879 & n8880;
  assign n8882 = n8878 & ~n8881;
  assign n8883 = ~x817 & ~n8882;
  assign n8884 = x817 & ~n8872;
  assign n8885 = ~x818 & ~x822;
  assign n8886 = ~n8869 & n8885;
  assign n8887 = ~n8884 & n8886;
  assign n8888 = x817 & x818;
  assign n8889 = n8869 & n8888;
  assign n8890 = ~n8887 & ~n8889;
  assign n8891 = ~x821 & ~n8890;
  assign n7796 = x818 ^ x817;
  assign n8892 = n7796 & n8875;
  assign n8893 = n8871 & ~n8874;
  assign n8894 = x822 & n8889;
  assign n8895 = n8894 ^ n8888;
  assign n8896 = ~n8893 & n8895;
  assign n8897 = ~n8892 & ~n8896;
  assign n8898 = ~n8891 & n8897;
  assign n8899 = ~n8883 & n8898;
  assign n8931 = n8930 ^ n8899;
  assign n7795 = x822 ^ x821;
  assign n7797 = n7796 ^ n7795;
  assign n7794 = x820 ^ x819;
  assign n7798 = n7797 ^ n7794;
  assign n7800 = x816 ^ x815;
  assign n7802 = n7801 ^ n7800;
  assign n7799 = x814 ^ x813;
  assign n7803 = n7802 ^ n7799;
  assign n8934 = n7798 & n7803;
  assign n9094 = n8931 & n8934;
  assign n9095 = n8899 & n8930;
  assign n9096 = ~n9094 & ~n9095;
  assign n9092 = n8878 & n8897;
  assign n9091 = n8909 & n8928;
  assign n9093 = n9092 ^ n9091;
  assign n9097 = n9096 ^ n9093;
  assign n8937 = x803 & x804;
  assign n8938 = x801 & x802;
  assign n8939 = ~n8937 & ~n8938;
  assign n8940 = ~x803 & ~x804;
  assign n8941 = ~x801 & ~x802;
  assign n8942 = ~n8940 & ~n8941;
  assign n8943 = ~n8939 & n8942;
  assign n8944 = x800 & n8943;
  assign n8945 = n8937 & n8938;
  assign n8946 = ~n8944 & ~n8945;
  assign n8947 = n8939 & ~n8942;
  assign n8948 = ~x800 & n8947;
  assign n8949 = n8946 & ~n8948;
  assign n8950 = ~x799 & ~n8949;
  assign n8951 = ~n8945 & ~n8947;
  assign n8952 = x800 & ~n8951;
  assign n8953 = ~x800 & ~n8943;
  assign n8954 = x799 & ~n8953;
  assign n8955 = ~n8952 & n8954;
  assign n7785 = x800 ^ x799;
  assign n8956 = n8940 & n8941;
  assign n8957 = n7785 & n8956;
  assign n8958 = ~n8955 & ~n8957;
  assign n8959 = ~n8950 & n8958;
  assign n8960 = ~x809 & ~x810;
  assign n8961 = ~x807 & ~x808;
  assign n8962 = ~n8960 & ~n8961;
  assign n8963 = x809 & x810;
  assign n8964 = x807 & x808;
  assign n8965 = ~n8963 & ~n8964;
  assign n8966 = n8962 & ~n8965;
  assign n8967 = x806 & n8966;
  assign n8968 = n8963 & n8964;
  assign n8969 = ~n8967 & ~n8968;
  assign n8970 = ~n8962 & n8965;
  assign n8971 = n8960 & n8961;
  assign n8972 = x806 & ~n8971;
  assign n8973 = n8970 & ~n8972;
  assign n8974 = n8969 & ~n8973;
  assign n8975 = ~x805 & ~n8974;
  assign n7790 = x806 ^ x805;
  assign n8976 = n7790 & n8966;
  assign n8977 = x805 & x806;
  assign n8978 = n8964 & n8977;
  assign n8979 = x810 & n8978;
  assign n8980 = n8979 ^ n8977;
  assign n8981 = ~n8970 & n8980;
  assign n8982 = ~n8976 & ~n8981;
  assign n8983 = ~x806 & ~x810;
  assign n8984 = n8961 & n8983;
  assign n8985 = ~n8978 & ~n8984;
  assign n8986 = ~x809 & ~n8985;
  assign n8987 = n8982 & ~n8986;
  assign n8988 = ~n8975 & n8987;
  assign n9102 = ~n8959 & ~n8988;
  assign n7789 = x808 ^ x807;
  assign n7791 = n7790 ^ n7789;
  assign n7788 = x810 ^ x809;
  assign n7792 = n7791 ^ n7788;
  assign n7784 = x802 ^ x801;
  assign n7786 = n7785 ^ n7784;
  assign n7783 = x804 ^ x803;
  assign n7787 = n7786 ^ n7783;
  assign n7793 = n7792 ^ n7787;
  assign n7804 = n7803 ^ n7798;
  assign n8932 = n7793 & n7804;
  assign n8933 = n7787 & n7792;
  assign n9103 = ~n8932 & ~n8933;
  assign n9104 = n9102 & n9103;
  assign n9105 = n8959 & n8988;
  assign n8989 = n8988 ^ n8959;
  assign n8935 = n8934 ^ n8933;
  assign n8936 = ~n8932 & ~n8935;
  assign n8990 = n8989 ^ n8936;
  assign n8991 = n8990 ^ n8931;
  assign n9106 = n8934 ^ n8931;
  assign n9107 = ~n8991 & ~n9106;
  assign n9108 = ~n9105 & n9107;
  assign n9109 = ~n9104 & ~n9108;
  assign n9098 = n8969 & n8982;
  assign n9099 = n8946 & ~n8955;
  assign n9796 = n9098 & n9099;
  assign n9797 = n9109 & n9796;
  assign n9100 = n9099 ^ n9098;
  assign n9110 = ~n9103 & n9105;
  assign n9111 = n8991 & n9110;
  assign n9798 = n9100 & ~n9111;
  assign n9799 = ~n9797 & ~n9798;
  assign n9800 = ~n9097 & ~n9799;
  assign n9801 = n9099 ^ n9097;
  assign n9802 = n9109 & ~n9801;
  assign n9803 = n9802 ^ n9099;
  assign n9804 = ~n9098 & ~n9803;
  assign n9805 = ~n9800 & ~n9804;
  assign n9806 = n9097 & n9109;
  assign n9807 = n9099 & ~n9111;
  assign n9808 = n9806 & ~n9807;
  assign n9809 = n9805 & ~n9808;
  assign n9793 = n9096 ^ n9092;
  assign n9794 = ~n9093 & n9793;
  assign n9795 = n9794 ^ n9096;
  assign n9810 = n9809 ^ n9795;
  assign n8776 = x839 & x840;
  assign n8777 = x837 & x838;
  assign n8778 = ~n8776 & ~n8777;
  assign n8779 = ~x839 & ~x840;
  assign n8780 = ~x837 & ~x838;
  assign n8781 = ~n8779 & ~n8780;
  assign n8782 = ~n8778 & n8781;
  assign n8783 = x836 & n8782;
  assign n8784 = n8776 & n8777;
  assign n8785 = ~n8783 & ~n8784;
  assign n8786 = x836 & ~n8779;
  assign n8787 = ~n8776 & n8780;
  assign n8788 = ~n8786 & n8787;
  assign n8789 = n8785 & ~n8788;
  assign n8790 = ~x835 & ~n8789;
  assign n7813 = x838 ^ x837;
  assign n7812 = x836 ^ x835;
  assign n7814 = n7813 ^ n7812;
  assign n8791 = ~x836 & ~x840;
  assign n8792 = ~n8777 & n8791;
  assign n8793 = n7814 & n8792;
  assign n8794 = x835 & x836;
  assign n8795 = n8777 & n8794;
  assign n8796 = ~n8793 & ~n8795;
  assign n8797 = ~x839 & ~n8796;
  assign n8798 = n8778 & ~n8781;
  assign n8799 = x840 & n8795;
  assign n8800 = n8799 ^ n8794;
  assign n8801 = ~n8798 & n8800;
  assign n8802 = n7812 & n8782;
  assign n8803 = ~n8801 & ~n8802;
  assign n8804 = ~n8797 & n8803;
  assign n8805 = ~n8790 & n8804;
  assign n8746 = x845 & x846;
  assign n8747 = x843 & x844;
  assign n8748 = ~n8746 & ~n8747;
  assign n8749 = ~x845 & ~x846;
  assign n8750 = ~x843 & ~x844;
  assign n8751 = ~n8749 & ~n8750;
  assign n8752 = ~n8748 & n8751;
  assign n8753 = x842 & n8752;
  assign n8754 = n8746 & n8747;
  assign n8755 = ~n8753 & ~n8754;
  assign n8756 = x842 & ~n8749;
  assign n8757 = ~n8746 & n8750;
  assign n8758 = ~n8756 & n8757;
  assign n8759 = n8755 & ~n8758;
  assign n8760 = ~x841 & ~n8759;
  assign n7808 = x844 ^ x843;
  assign n7807 = x842 ^ x841;
  assign n7809 = n7808 ^ n7807;
  assign n8761 = ~x842 & ~x846;
  assign n8762 = ~n8747 & n8761;
  assign n8763 = n7809 & n8762;
  assign n8764 = x841 & x842;
  assign n8765 = n8747 & n8764;
  assign n8766 = ~n8763 & ~n8765;
  assign n8767 = ~x845 & ~n8766;
  assign n8768 = n8748 & ~n8751;
  assign n8769 = x846 & n8765;
  assign n8770 = n8769 ^ n8764;
  assign n8771 = ~n8768 & n8770;
  assign n8772 = n7807 & n8752;
  assign n8773 = ~n8771 & ~n8772;
  assign n8774 = ~n8767 & n8773;
  assign n8775 = ~n8760 & n8774;
  assign n8806 = n8805 ^ n8775;
  assign n7811 = x840 ^ x839;
  assign n7815 = n7814 ^ n7811;
  assign n7806 = x846 ^ x845;
  assign n7810 = n7809 ^ n7806;
  assign n7816 = n7815 ^ n7810;
  assign n7824 = x824 ^ x823;
  assign n7823 = x826 ^ x825;
  assign n7825 = n7824 ^ n7823;
  assign n7822 = x828 ^ x827;
  assign n7826 = n7825 ^ n7822;
  assign n7819 = x830 ^ x829;
  assign n7818 = x832 ^ x831;
  assign n7820 = n7819 ^ n7818;
  assign n7817 = x834 ^ x833;
  assign n7821 = n7820 ^ n7817;
  assign n7827 = n7826 ^ n7821;
  assign n8743 = n7816 & n7827;
  assign n8744 = n7810 & n7815;
  assign n8745 = ~n8743 & ~n8744;
  assign n8807 = n8806 ^ n8745;
  assign n8834 = x827 & x828;
  assign n8835 = n8834 ^ x826;
  assign n8836 = n7823 & ~n8835;
  assign n8837 = n8836 ^ x825;
  assign n8838 = n7824 & n8837;
  assign n8839 = ~x825 & ~x826;
  assign n8840 = ~n8834 & n8839;
  assign n8841 = x825 & x826;
  assign n8842 = x823 & x824;
  assign n8843 = ~n8841 & n8842;
  assign n8844 = ~n8840 & n8843;
  assign n8845 = ~n8838 & ~n8844;
  assign n8846 = ~x827 & ~x828;
  assign n8847 = ~n8845 & ~n8846;
  assign n8848 = n8841 & n8842;
  assign n8849 = ~x828 & n8848;
  assign n8850 = ~n8847 & ~n8849;
  assign n8851 = n8834 & n8841;
  assign n8852 = x824 & ~n8846;
  assign n8853 = ~n8851 & ~n8852;
  assign n8854 = n8837 & ~n8853;
  assign n8855 = n8840 & ~n8852;
  assign n8856 = ~n8854 & ~n8855;
  assign n8857 = ~x823 & ~n8856;
  assign n8858 = ~x824 & ~x828;
  assign n8859 = ~n8841 & n8858;
  assign n8860 = n7825 & n8859;
  assign n8861 = ~n8848 & ~n8860;
  assign n8862 = ~x827 & ~n8861;
  assign n8863 = ~n8857 & ~n8862;
  assign n8864 = n8850 & n8863;
  assign n8833 = n7821 & n7826;
  assign n8865 = n8864 ^ n8833;
  assign n8808 = x831 & x832;
  assign n8809 = x833 & x834;
  assign n8810 = n8808 & n8809;
  assign n8811 = ~x833 & ~x834;
  assign n8812 = ~n8808 & n8811;
  assign n8813 = ~n8810 & ~n8812;
  assign n8814 = ~x831 & ~x832;
  assign n8815 = ~n8809 & n8814;
  assign n8816 = x829 & x830;
  assign n8817 = ~n8815 & n8816;
  assign n8818 = n8813 & n8817;
  assign n8819 = n7819 & ~n8811;
  assign n8820 = n8809 ^ x832;
  assign n8821 = n7818 & ~n8820;
  assign n8822 = n8821 ^ x831;
  assign n8823 = n8819 & n8822;
  assign n8824 = ~n8818 & ~n8823;
  assign n8825 = x830 & ~n8811;
  assign n8826 = n8815 & ~n8825;
  assign n8827 = ~n8810 & ~n8826;
  assign n8828 = ~x829 & ~n8827;
  assign n8829 = n8824 & ~n8828;
  assign n8830 = ~x830 & n8812;
  assign n8831 = n7820 & n8830;
  assign n8832 = n8829 & ~n8831;
  assign n8866 = n8865 ^ n8832;
  assign n9085 = ~n8807 & n8866;
  assign n9086 = n8743 & n8806;
  assign n9087 = ~n9085 & ~n9086;
  assign n9082 = n8785 & n8803;
  assign n9081 = n8755 & n8773;
  assign n9083 = n9082 ^ n9081;
  assign n9078 = n8775 ^ n8744;
  assign n9079 = n8806 & ~n9078;
  assign n9080 = n9079 ^ n8805;
  assign n9084 = n9083 ^ n9080;
  assign n9088 = n9087 ^ n9084;
  assign n9075 = n8850 & ~n8854;
  assign n9074 = ~n8810 & n8824;
  assign n9076 = n9075 ^ n9074;
  assign n9071 = n8833 ^ n8832;
  assign n9072 = n8865 & ~n9071;
  assign n9073 = n9072 ^ n8864;
  assign n9077 = n9076 ^ n9073;
  assign n9089 = n9088 ^ n9077;
  assign n8867 = n8866 ^ n8807;
  assign n7805 = n7804 ^ n7793;
  assign n7828 = n7827 ^ n7816;
  assign n8742 = n7805 & n7828;
  assign n8868 = n8867 ^ n8742;
  assign n9068 = n8991 ^ n8867;
  assign n9069 = n8868 & n9068;
  assign n9070 = n9069 ^ n8991;
  assign n9090 = n9089 ^ n9070;
  assign n9112 = n9109 & ~n9111;
  assign n9101 = n9100 ^ n9097;
  assign n9113 = n9112 ^ n9101;
  assign n9790 = n9113 ^ n9089;
  assign n9791 = ~n9090 & n9790;
  assign n9792 = n9791 ^ n9113;
  assign n9811 = n9810 ^ n9792;
  assign n9776 = ~n9084 & n9087;
  assign n9777 = n9073 & ~n9776;
  assign n9778 = ~n9074 & ~n9075;
  assign n9779 = ~n9777 & ~n9778;
  assign n9780 = n9074 & n9075;
  assign n9781 = n9089 & ~n9780;
  assign n9782 = n9779 & ~n9781;
  assign n9783 = n9084 & ~n9087;
  assign n9784 = ~n9777 & ~n9783;
  assign n9785 = n9781 & ~n9784;
  assign n9786 = ~n9782 & ~n9785;
  assign n9773 = n9082 ^ n9080;
  assign n9774 = ~n9083 & ~n9773;
  assign n9775 = n9774 ^ n9080;
  assign n9787 = n9786 ^ n9775;
  assign n9788 = n9779 & n9783;
  assign n9789 = ~n9787 & ~n9788;
  assign n9812 = n9811 ^ n9789;
  assign n8564 = n8563 ^ n8504;
  assign n8618 = n8617 ^ n8564;
  assign n7852 = n7851 ^ n7840;
  assign n8495 = n7852 & n7875;
  assign n8496 = n7868 ^ n7863;
  assign n8497 = n7874 & ~n8496;
  assign n8498 = n8497 ^ n7873;
  assign n8499 = ~n8495 & ~n8498;
  assign n8501 = n7863 & n8500;
  assign n8502 = n7852 & n8501;
  assign n8503 = ~n8499 & ~n8502;
  assign n8619 = n8618 ^ n8503;
  assign n9028 = n8619 & n8740;
  assign n9029 = n8498 & ~n8502;
  assign n9030 = n9029 ^ n8499;
  assign n9031 = n8618 & n9030;
  assign n9032 = n9031 ^ n8499;
  assign n9033 = ~n9028 & ~n9032;
  assign n9065 = n9064 ^ n9033;
  assign n9017 = n9016 ^ n9013;
  assign n9027 = n9026 ^ n9017;
  assign n9066 = n9065 ^ n9027;
  assign n7829 = n7828 ^ n7805;
  assign n7876 = n7875 ^ n7852;
  assign n8995 = n7829 & n7876;
  assign n8992 = n8991 ^ n8868;
  assign n9004 = n8995 ^ n8992;
  assign n8741 = n8740 ^ n8619;
  assign n9005 = n8995 ^ n8741;
  assign n9006 = n9004 & n9005;
  assign n9007 = n9006 ^ n8992;
  assign n9067 = n9066 ^ n9007;
  assign n9114 = n9113 ^ n9090;
  assign n9770 = n9114 ^ n9007;
  assign n9771 = n9067 & n9770;
  assign n9772 = n9771 ^ n9066;
  assign n9813 = n9812 ^ n9772;
  assign n9848 = n9841 & n9847;
  assign n9852 = ~n9051 & n9846;
  assign n9853 = ~n9851 & ~n9852;
  assign n9854 = ~n9848 & n9853;
  assign n9855 = n9854 ^ n9837;
  assign n9834 = n9833 ^ n9820;
  assign n9856 = n9855 ^ n9834;
  assign n9814 = n9033 ^ n9027;
  assign n9815 = n9065 & ~n9814;
  assign n9816 = n9815 ^ n9064;
  assign n9857 = n9856 ^ n9816;
  assign n9970 = n9857 ^ n9812;
  assign n9971 = ~n9813 & ~n9970;
  assign n9972 = n9971 ^ n9857;
  assign n9978 = n9977 ^ n9972;
  assign n9962 = ~n9098 & ~n9099;
  assign n9963 = n9810 & ~n9962;
  assign n9964 = n9803 & ~n9807;
  assign n9965 = n9795 & ~n9964;
  assign n9966 = ~n9963 & ~n9965;
  assign n9960 = ~n9775 & ~n9785;
  assign n9961 = ~n9782 & ~n9960;
  assign n9967 = n9966 ^ n9961;
  assign n9957 = n9792 ^ n9789;
  assign n9958 = ~n9811 & ~n9957;
  assign n9959 = n9958 ^ n9810;
  assign n9968 = n9967 ^ n9959;
  assign n9954 = n9834 ^ n9816;
  assign n9955 = ~n9856 & n9954;
  assign n9956 = n9955 ^ n9855;
  assign n9969 = n9968 ^ n9956;
  assign n9979 = n9978 ^ n9969;
  assign n10002 = n9956 & n9968;
  assign n10003 = n9975 & ~n9976;
  assign n10004 = n10002 & ~n10003;
  assign n10005 = ~n9972 & n10004;
  assign n10010 = ~n9975 & n9976;
  assign n10061 = ~n10005 & ~n10010;
  assign n10062 = ~n9956 & n10061;
  assign n10063 = n9979 & n10062;
  assign n10006 = ~n9968 & n10003;
  assign n10064 = n9972 & n10006;
  assign n10065 = ~n9961 & ~n9966;
  assign n10066 = ~n9959 & n10065;
  assign n10067 = ~n10064 & ~n10066;
  assign n10068 = ~n10063 & n10067;
  assign n9999 = n9966 ^ n9959;
  assign n10000 = ~n9967 & n9999;
  assign n10001 = n10000 ^ n9959;
  assign n10009 = ~n9956 & n9972;
  assign n10069 = ~n10009 & ~n10061;
  assign n10070 = ~n10001 & ~n10069;
  assign n10071 = n10068 & ~n10070;
  assign n9988 = n9946 ^ n9944;
  assign n9989 = ~n9950 & ~n9988;
  assign n9990 = n9989 ^ n9949;
  assign n10007 = ~n9956 & n10006;
  assign n10008 = ~n10005 & ~n10007;
  assign n10011 = n9968 & n10010;
  assign n10012 = ~n10009 & n10011;
  assign n10013 = n10008 & ~n10012;
  assign n10014 = ~n10002 & n10003;
  assign n10015 = ~n9956 & ~n9968;
  assign n10016 = ~n10010 & n10015;
  assign n10017 = ~n10014 & ~n10016;
  assign n10018 = n9972 & ~n10017;
  assign n10019 = n10013 & ~n10018;
  assign n10020 = n10019 ^ n10001;
  assign n9953 = n9952 ^ n9932;
  assign n9980 = n9979 ^ n9953;
  assign n9768 = n9767 ^ n9728;
  assign n9219 = n9218 ^ n9121;
  assign n9115 = n9114 ^ n9067;
  assign n9220 = n9219 ^ n9115;
  assign n8993 = n8992 ^ n8741;
  assign n8234 = n8233 ^ n7980;
  assign n8494 = n8493 ^ n8234;
  assign n8994 = n8993 ^ n8494;
  assign n8996 = n8995 ^ n8994;
  assign n7877 = n7876 ^ n7829;
  assign n7972 = n7971 ^ n7924;
  assign n8997 = n7877 & n7972;
  assign n9221 = ~n8996 & ~n8997;
  assign n9222 = ~n8993 & n8997;
  assign n9223 = ~n8494 & ~n9222;
  assign n9224 = ~n9221 & ~n9223;
  assign n9682 = n9224 ^ n9115;
  assign n9683 = n9220 & n9682;
  assign n9684 = n9683 ^ n9219;
  assign n9769 = n9768 ^ n9684;
  assign n9858 = n9857 ^ n9813;
  assign n9927 = n9858 ^ n9768;
  assign n9928 = n9769 & ~n9927;
  assign n9929 = n9928 ^ n9858;
  assign n9996 = n9953 ^ n9929;
  assign n9997 = ~n9980 & ~n9996;
  assign n9998 = n9997 ^ n9979;
  assign n10021 = n10020 ^ n9998;
  assign n10122 = n9990 & n10021;
  assign n10123 = n10071 & n10122;
  assign n10124 = n10081 & ~n10123;
  assign n10078 = n9990 & n10020;
  assign n10125 = n9998 & n10020;
  assign n10126 = ~n10071 & ~n10125;
  assign n10127 = ~n10078 & n10126;
  assign n10128 = ~n10124 & ~n10127;
  assign n10077 = n9987 & ~n9993;
  assign n10129 = ~n9990 & ~n10021;
  assign n10130 = ~n9998 & ~n10071;
  assign n10131 = ~n10129 & ~n10130;
  assign n10132 = ~n10077 & ~n10131;
  assign n10133 = n10128 & ~n10132;
  assign n7316 = ~x615 & ~x616;
  assign n7317 = ~x617 & ~x618;
  assign n7318 = ~n7316 & ~n7317;
  assign n7319 = x615 & x616;
  assign n7320 = x617 & x618;
  assign n7321 = ~n7319 & ~n7320;
  assign n7322 = n7318 & ~n7321;
  assign n7323 = x614 & n7322;
  assign n7324 = n7319 & n7320;
  assign n7325 = ~n7323 & ~n7324;
  assign n7326 = ~n7318 & n7321;
  assign n7327 = n7316 & n7317;
  assign n7328 = x614 & ~n7327;
  assign n7329 = n7326 & ~n7328;
  assign n7330 = n7325 & ~n7329;
  assign n7331 = ~x613 & ~n7330;
  assign n6811 = x614 ^ x613;
  assign n7332 = n6811 & n7322;
  assign n7333 = x613 & x614;
  assign n7334 = n7319 & n7333;
  assign n7335 = x618 & n7334;
  assign n7336 = n7335 ^ n7333;
  assign n7337 = ~n7326 & n7336;
  assign n7338 = ~n7332 & ~n7337;
  assign n7339 = ~x614 & ~x618;
  assign n7340 = n7316 & n7339;
  assign n7341 = ~n7334 & ~n7340;
  assign n7342 = ~x617 & ~n7341;
  assign n7343 = n7338 & ~n7342;
  assign n7344 = ~n7331 & n7343;
  assign n7286 = x609 & x610;
  assign n7287 = x611 & x612;
  assign n7288 = ~n7286 & ~n7287;
  assign n7289 = ~x609 & ~x610;
  assign n7290 = ~x611 & ~x612;
  assign n7291 = ~n7289 & ~n7290;
  assign n7292 = ~n7288 & n7291;
  assign n7293 = x608 & n7292;
  assign n7294 = n7286 & n7287;
  assign n7295 = ~n7293 & ~n7294;
  assign n7296 = x608 & ~n7290;
  assign n7297 = ~n7287 & n7289;
  assign n7298 = ~n7296 & n7297;
  assign n7299 = n7295 & ~n7298;
  assign n7300 = ~x607 & ~n7299;
  assign n6806 = x608 ^ x607;
  assign n7301 = n6806 & n7292;
  assign n7302 = n7288 & ~n7291;
  assign n7303 = x612 & n7286;
  assign n7304 = x607 & x608;
  assign n7305 = ~n7303 & n7304;
  assign n7306 = ~n7302 & n7305;
  assign n7307 = ~n7301 & ~n7306;
  assign n6805 = x610 ^ x609;
  assign n6807 = n6806 ^ n6805;
  assign n7308 = ~x608 & ~n7286;
  assign n7309 = n7290 & n7308;
  assign n7310 = n6807 & n7309;
  assign n7311 = ~x611 & n7286;
  assign n7312 = n7304 & n7311;
  assign n7313 = ~n7310 & ~n7312;
  assign n7314 = n7307 & n7313;
  assign n7315 = ~n7300 & n7314;
  assign n7345 = n7344 ^ n7315;
  assign n6793 = x628 ^ x627;
  assign n7261 = x629 & x630;
  assign n7262 = n7261 ^ x628;
  assign n7263 = ~n6793 & ~n7262;
  assign n7264 = ~x625 & n7263;
  assign n7265 = x627 & x628;
  assign n7266 = ~x629 & ~x630;
  assign n7267 = ~n7265 & n7266;
  assign n7268 = ~x626 & n7267;
  assign n7269 = ~n7264 & ~n7268;
  assign n7270 = ~x627 & ~x628;
  assign n7271 = x625 & ~n7270;
  assign n7272 = x626 & ~n7266;
  assign n7273 = ~n7271 & ~n7272;
  assign n7274 = ~n7269 & n7273;
  assign n6795 = x626 ^ x625;
  assign n7275 = n7261 & ~n7270;
  assign n7276 = n7265 & ~n7266;
  assign n7277 = ~n7275 & ~n7276;
  assign n7278 = n6795 & ~n7277;
  assign n7279 = x625 & x626;
  assign n7280 = ~n7267 & n7279;
  assign n7281 = ~n7263 & n7280;
  assign n7282 = ~n7278 & ~n7281;
  assign n7283 = ~n7274 & n7282;
  assign n6798 = x622 ^ x621;
  assign n7238 = x623 & x624;
  assign n7239 = n7238 ^ x622;
  assign n7240 = ~n6798 & ~n7239;
  assign n7241 = ~x619 & n7240;
  assign n7242 = x621 & x622;
  assign n7243 = ~x623 & ~x624;
  assign n7244 = ~n7242 & n7243;
  assign n7245 = ~x620 & n7244;
  assign n7246 = ~n7241 & ~n7245;
  assign n7247 = ~x621 & ~x622;
  assign n7248 = x619 & ~n7247;
  assign n7249 = x620 & ~n7243;
  assign n7250 = ~n7248 & ~n7249;
  assign n7251 = ~n7246 & n7250;
  assign n6800 = x620 ^ x619;
  assign n7252 = n7238 & ~n7247;
  assign n7253 = n7242 & ~n7243;
  assign n7254 = ~n7252 & ~n7253;
  assign n7255 = n6800 & ~n7254;
  assign n7256 = x619 & x620;
  assign n7257 = ~n7244 & n7256;
  assign n7258 = ~n7240 & n7257;
  assign n7259 = ~n7255 & ~n7258;
  assign n7260 = ~n7251 & n7259;
  assign n7284 = n7283 ^ n7260;
  assign n6799 = x624 ^ x623;
  assign n6801 = n6800 ^ n6799;
  assign n6802 = n6801 ^ n6798;
  assign n6794 = x630 ^ x629;
  assign n6796 = n6795 ^ n6794;
  assign n6797 = n6796 ^ n6793;
  assign n6803 = n6802 ^ n6797;
  assign n6810 = x616 ^ x615;
  assign n6812 = n6811 ^ n6810;
  assign n6809 = x618 ^ x617;
  assign n6813 = n6812 ^ n6809;
  assign n6804 = x612 ^ x611;
  assign n6808 = n6807 ^ n6804;
  assign n6814 = n6813 ^ n6808;
  assign n7233 = n6803 & n6814;
  assign n7235 = n6808 & n6813;
  assign n7234 = n6797 & n6802;
  assign n7236 = n7235 ^ n7234;
  assign n7237 = ~n7233 & ~n7236;
  assign n7285 = n7284 ^ n7237;
  assign n7346 = n7345 ^ n7285;
  assign n9472 = ~n7234 & n7284;
  assign n9473 = ~n7346 & ~n9472;
  assign n9474 = n7345 ^ n7235;
  assign n9475 = ~n7233 & ~n9474;
  assign n9476 = ~n9473 & ~n9475;
  assign n9471 = n7325 & n7338;
  assign n9477 = n9476 ^ n9471;
  assign n9468 = n7295 & n7307;
  assign n9465 = n7315 ^ n7235;
  assign n9466 = n7345 & ~n9465;
  assign n9467 = n9466 ^ n7344;
  assign n9469 = n9468 ^ n9467;
  assign n9461 = n7261 & n7265;
  assign n9462 = n7282 & ~n9461;
  assign n9459 = n7238 & n7242;
  assign n9460 = n7259 & ~n9459;
  assign n9463 = n9462 ^ n9460;
  assign n9456 = n7260 ^ n7234;
  assign n9457 = n7284 & ~n9456;
  assign n9458 = n9457 ^ n7283;
  assign n9464 = n9463 ^ n9458;
  assign n9470 = n9469 ^ n9464;
  assign n9478 = n9477 ^ n9470;
  assign n9519 = n9471 & ~n9476;
  assign n9520 = ~n9467 & n9468;
  assign n9521 = ~n9519 & ~n9520;
  assign n9522 = n9464 & n9521;
  assign n9523 = ~n9478 & n9522;
  assign n9524 = ~n9464 & n9478;
  assign n9525 = n9524 ^ n9519;
  assign n9526 = n9520 ^ n9519;
  assign n9527 = n9525 & ~n9526;
  assign n9528 = n9527 ^ n9524;
  assign n9529 = ~n9523 & ~n9528;
  assign n9516 = n9462 ^ n9458;
  assign n9517 = ~n9463 & ~n9516;
  assign n9518 = n9517 ^ n9458;
  assign n9530 = n9529 ^ n9518;
  assign n6772 = x638 ^ x637;
  assign n6771 = x640 ^ x639;
  assign n7200 = x641 & x642;
  assign n7201 = n7200 ^ x640;
  assign n7202 = n6771 & ~n7201;
  assign n7203 = n7202 ^ x639;
  assign n7204 = n6772 & n7203;
  assign n7205 = ~x639 & ~x640;
  assign n7206 = ~n7200 & n7205;
  assign n7207 = x639 & x640;
  assign n7208 = x637 & x638;
  assign n7209 = ~n7207 & n7208;
  assign n7210 = ~n7206 & n7209;
  assign n7211 = ~n7204 & ~n7210;
  assign n7212 = ~x641 & ~x642;
  assign n7213 = ~n7211 & ~n7212;
  assign n7214 = n7207 & n7208;
  assign n7215 = ~x642 & n7214;
  assign n7216 = ~n7213 & ~n7215;
  assign n7217 = x638 & ~n7212;
  assign n7218 = n7200 & n7207;
  assign n7219 = ~n7217 & ~n7218;
  assign n7220 = n7203 & ~n7219;
  assign n7221 = n7206 & ~n7217;
  assign n7222 = ~n7220 & ~n7221;
  assign n7223 = ~x637 & ~n7222;
  assign n7224 = n7216 & ~n7223;
  assign n6773 = n6772 ^ n6771;
  assign n7225 = ~x638 & ~x642;
  assign n7226 = ~n7207 & n7225;
  assign n7227 = n6773 & n7226;
  assign n7228 = ~n7214 & ~n7227;
  assign n7229 = ~x641 & ~n7228;
  assign n7230 = n7224 & ~n7229;
  assign n7171 = x633 & x634;
  assign n7172 = x635 & x636;
  assign n7173 = ~n7171 & ~n7172;
  assign n7174 = ~x633 & ~x634;
  assign n7175 = ~x635 & ~x636;
  assign n7176 = ~n7174 & ~n7175;
  assign n7177 = ~n7173 & n7176;
  assign n7178 = x632 & n7177;
  assign n7179 = n7171 & n7172;
  assign n7180 = ~n7178 & ~n7179;
  assign n7181 = n7173 & ~n7176;
  assign n7182 = ~x632 & n7181;
  assign n7183 = n7174 & n7175;
  assign n7184 = ~n7182 & ~n7183;
  assign n7185 = n7180 & n7184;
  assign n7186 = ~x631 & ~n7185;
  assign n6777 = x632 ^ x631;
  assign n7187 = n6777 & n7177;
  assign n7188 = x631 & x632;
  assign n7189 = n7171 & n7188;
  assign n7190 = x636 & n7189;
  assign n7191 = n7190 ^ n7188;
  assign n7192 = ~n7181 & n7191;
  assign n7193 = ~n7187 & ~n7192;
  assign n7194 = ~x632 & ~x636;
  assign n7195 = n7174 & n7194;
  assign n7196 = ~n7189 & ~n7195;
  assign n7197 = ~x635 & ~n7196;
  assign n7198 = n7193 & ~n7197;
  assign n7199 = ~n7186 & n7198;
  assign n7231 = n7230 ^ n7199;
  assign n7139 = x651 & x652;
  assign n7140 = x653 & x654;
  assign n7141 = ~n7139 & ~n7140;
  assign n7142 = ~x653 & ~x654;
  assign n7143 = ~x651 & ~x652;
  assign n7144 = ~n7142 & ~n7143;
  assign n7145 = ~n7141 & n7144;
  assign n7146 = x650 & n7145;
  assign n7147 = n7139 & n7140;
  assign n7148 = ~n7146 & ~n7147;
  assign n7149 = x650 & ~n7142;
  assign n7150 = ~n7140 & n7143;
  assign n7151 = ~n7149 & n7150;
  assign n7152 = n7148 & ~n7151;
  assign n7153 = ~x649 & ~n7152;
  assign n6783 = x650 ^ x649;
  assign n7154 = n6783 & n7145;
  assign n7155 = n7141 & ~n7144;
  assign n7156 = x654 & n7139;
  assign n7157 = x649 & x650;
  assign n7158 = ~n7156 & n7157;
  assign n7159 = ~n7155 & n7158;
  assign n7160 = ~n7154 & ~n7159;
  assign n6782 = x652 ^ x651;
  assign n6784 = n6783 ^ n6782;
  assign n7161 = ~x650 & ~n7139;
  assign n7162 = n7142 & n7161;
  assign n7163 = n6784 & n7162;
  assign n7164 = ~x653 & n7139;
  assign n7165 = n7157 & n7164;
  assign n7166 = ~n7163 & ~n7165;
  assign n7167 = n7160 & n7166;
  assign n7168 = ~n7153 & n7167;
  assign n6788 = x644 ^ x643;
  assign n7119 = x645 & x646;
  assign n7120 = x647 & x648;
  assign n7121 = ~n7119 & ~n7120;
  assign n7122 = ~x645 & ~x646;
  assign n7123 = ~x647 & ~x648;
  assign n7124 = ~n7122 & ~n7123;
  assign n7125 = n7121 & ~n7124;
  assign n7126 = ~n6788 & n7125;
  assign n7127 = n7119 & n7120;
  assign n7128 = n7122 & n7123;
  assign n7129 = ~n7127 & ~n7128;
  assign n7130 = ~n7126 & n7129;
  assign n7131 = x643 & x644;
  assign n7132 = ~n7130 & ~n7131;
  assign n7133 = n6788 & n7124;
  assign n7134 = ~n7121 & n7133;
  assign n7135 = ~n7127 & n7131;
  assign n7136 = ~n7125 & n7135;
  assign n7137 = ~n7134 & ~n7136;
  assign n7138 = ~n7132 & n7137;
  assign n7169 = n7168 ^ n7138;
  assign n6776 = x634 ^ x633;
  assign n6778 = n6777 ^ n6776;
  assign n6775 = x636 ^ x635;
  assign n6779 = n6778 ^ n6775;
  assign n6787 = x648 ^ x647;
  assign n6789 = n6788 ^ n6787;
  assign n6786 = x646 ^ x645;
  assign n6790 = n6789 ^ n6786;
  assign n6770 = x642 ^ x641;
  assign n6774 = n6773 ^ n6770;
  assign n7114 = n6790 ^ n6774;
  assign n6781 = x654 ^ x653;
  assign n6785 = n6784 ^ n6781;
  assign n7116 = n7114 ^ n6785;
  assign n7117 = ~n6779 & n7116;
  assign n6791 = n6790 ^ n6785;
  assign n7115 = ~n6791 & ~n7114;
  assign n7118 = n7117 ^ n7115;
  assign n7170 = n7169 ^ n7118;
  assign n7232 = n7231 ^ n7170;
  assign n7347 = n7346 ^ n7232;
  assign n6780 = n6779 ^ n6774;
  assign n6792 = n6791 ^ n6780;
  assign n6815 = n6814 ^ n6803;
  assign n6871 = n6792 & n6815;
  assign n9453 = n7232 ^ n6871;
  assign n9454 = n7347 & n9453;
  assign n9455 = n9454 ^ n7346;
  assign n9479 = n9478 ^ n9455;
  assign n9441 = ~n6785 & ~n6790;
  assign n9442 = ~n7169 & ~n9441;
  assign n9443 = n7232 & n9442;
  assign n9431 = n6785 & n6790;
  assign n9444 = n7169 & ~n9431;
  assign n9445 = ~n9443 & ~n9444;
  assign n9446 = ~n6774 & ~n6779;
  assign n9447 = n7170 & ~n9446;
  assign n9427 = n6774 & n6779;
  assign n9448 = n9447 ^ n9427;
  assign n9449 = ~n7231 & ~n9448;
  assign n9450 = n9449 ^ n9427;
  assign n9451 = ~n9445 & ~n9450;
  assign n9436 = ~n7127 & n7137;
  assign n9435 = n7148 & n7160;
  assign n9437 = n9436 ^ n9435;
  assign n9432 = n9431 ^ n7138;
  assign n9433 = n7169 & ~n9432;
  assign n9434 = n9433 ^ n7168;
  assign n9438 = n9437 ^ n9434;
  assign n9428 = n7231 & n9427;
  assign n9429 = n7199 & n7230;
  assign n9430 = ~n9428 & ~n9429;
  assign n9439 = n9438 ^ n9430;
  assign n9425 = n7216 & ~n7220;
  assign n9424 = n7180 & n7193;
  assign n9426 = n9425 ^ n9424;
  assign n9440 = n9439 ^ n9426;
  assign n9452 = n9451 ^ n9440;
  assign n9513 = n9455 ^ n9452;
  assign n9514 = ~n9479 & ~n9513;
  assign n9515 = n9514 ^ n9478;
  assign n9531 = n9530 ^ n9515;
  assign n9496 = n9430 & ~n9438;
  assign n9497 = n9496 ^ n9430;
  assign n9498 = ~n9451 & ~n9497;
  assign n9499 = n9498 ^ n9430;
  assign n9500 = n9426 & n9499;
  assign n9501 = n9424 & n9425;
  assign n9502 = ~n9438 & ~n9501;
  assign n9503 = n9440 & n9502;
  assign n9504 = ~n9500 & ~n9503;
  assign n9505 = ~n9439 & ~n9451;
  assign n9506 = ~n9496 & ~n9505;
  assign n9507 = n9501 & n9506;
  assign n9508 = ~n9424 & ~n9425;
  assign n9509 = n9505 & n9508;
  assign n9510 = ~n9507 & ~n9509;
  assign n9511 = n9504 & n9510;
  assign n9493 = n9436 ^ n9434;
  assign n9494 = ~n9437 & ~n9493;
  assign n9495 = n9494 ^ n9434;
  assign n9512 = n9511 ^ n9495;
  assign n9906 = n9515 ^ n9512;
  assign n9907 = n9531 & n9906;
  assign n9908 = n9907 ^ n9530;
  assign n6853 = x560 ^ x559;
  assign n7037 = x561 & x562;
  assign n7038 = x563 & x564;
  assign n7039 = ~n7037 & ~n7038;
  assign n7040 = ~x561 & ~x562;
  assign n7041 = ~x563 & ~x564;
  assign n7042 = ~n7040 & ~n7041;
  assign n7043 = ~n7039 & n7042;
  assign n7044 = n6853 & n7043;
  assign n7045 = n7037 & n7038;
  assign n7046 = ~n7044 & ~n7045;
  assign n7047 = n7039 & ~n7042;
  assign n7048 = x559 & x560;
  assign n7049 = ~n7045 & n7048;
  assign n7050 = ~n7047 & n7049;
  assign n7051 = n7046 & ~n7050;
  assign n7012 = x569 & x570;
  assign n7018 = x567 & x568;
  assign n7019 = n7012 & n7018;
  assign n7013 = ~x567 & ~x568;
  assign n7014 = ~n7012 & n7013;
  assign n7015 = ~x569 & ~x570;
  assign n7021 = n7015 & ~n7018;
  assign n7025 = ~n7014 & ~n7021;
  assign n7026 = x565 & x566;
  assign n7027 = ~n7019 & n7026;
  assign n7028 = n7025 & n7027;
  assign n6858 = x566 ^ x565;
  assign n7029 = n7012 & ~n7013;
  assign n7030 = ~n7015 & n7018;
  assign n7031 = ~n7029 & ~n7030;
  assign n7032 = n6858 & ~n7031;
  assign n7033 = ~n7028 & ~n7032;
  assign n9392 = ~n7019 & n7033;
  assign n9575 = ~n7051 & ~n9392;
  assign n7016 = x566 & ~n7015;
  assign n7017 = n7014 & ~n7016;
  assign n7020 = ~n7017 & ~n7019;
  assign n7022 = ~x566 & n7021;
  assign n7023 = n7020 & ~n7022;
  assign n7024 = ~x565 & ~n7023;
  assign n7034 = n7013 & n7022;
  assign n7035 = n7033 & ~n7034;
  assign n7036 = ~n7024 & n7035;
  assign n7052 = ~n6853 & n7047;
  assign n7053 = n7040 & n7041;
  assign n7054 = ~n7052 & ~n7053;
  assign n7055 = n7051 & n7054;
  assign n7056 = n7048 & ~n7050;
  assign n7057 = ~n7055 & ~n7056;
  assign n9403 = n7036 & ~n7057;
  assign n6852 = x564 ^ x563;
  assign n6854 = n6853 ^ n6852;
  assign n6851 = x562 ^ x561;
  assign n6855 = n6854 ^ n6851;
  assign n6857 = x568 ^ x567;
  assign n6859 = n6858 ^ n6857;
  assign n6856 = x570 ^ x569;
  assign n6860 = n6859 ^ n6856;
  assign n9404 = n6855 & n6860;
  assign n9405 = ~n9403 & ~n9404;
  assign n7087 = x579 & x580;
  assign n7088 = x581 & x582;
  assign n7089 = ~n7087 & ~n7088;
  assign n7090 = ~x579 & ~x580;
  assign n7091 = ~x581 & ~x582;
  assign n7092 = ~n7090 & ~n7091;
  assign n7093 = ~n7089 & n7092;
  assign n7094 = x578 & n7093;
  assign n7095 = n7087 & n7088;
  assign n7096 = ~n7094 & ~n7095;
  assign n7097 = n7089 & ~n7092;
  assign n7098 = ~x578 & n7097;
  assign n7099 = n7096 & ~n7098;
  assign n7100 = ~x577 & ~n7099;
  assign n7101 = ~n7095 & ~n7097;
  assign n7102 = x578 & ~n7101;
  assign n7103 = ~x578 & ~n7093;
  assign n7104 = x577 & ~n7103;
  assign n7105 = ~n7102 & n7104;
  assign n6847 = x578 ^ x577;
  assign n7106 = n7090 & n7091;
  assign n7107 = n6847 & n7106;
  assign n7108 = ~n7105 & ~n7107;
  assign n7109 = ~n7100 & n7108;
  assign n7064 = x573 & x574;
  assign n7065 = x575 & x576;
  assign n7066 = ~n7064 & ~n7065;
  assign n7067 = ~x573 & ~x574;
  assign n7068 = ~x575 & ~x576;
  assign n7069 = ~n7067 & ~n7068;
  assign n7070 = ~n7066 & n7069;
  assign n7071 = x572 & n7070;
  assign n7072 = n7064 & n7065;
  assign n7073 = ~n7071 & ~n7072;
  assign n7074 = n7066 & ~n7069;
  assign n7075 = ~x572 & n7074;
  assign n7076 = n7073 & ~n7075;
  assign n7077 = ~x571 & ~n7076;
  assign n7078 = ~n7072 & ~n7074;
  assign n7079 = x572 & ~n7078;
  assign n7080 = ~x572 & ~n7070;
  assign n7081 = x571 & ~n7080;
  assign n7082 = ~n7079 & n7081;
  assign n6842 = x572 ^ x571;
  assign n7083 = n7067 & n7068;
  assign n7084 = n6842 & n7083;
  assign n7085 = ~n7082 & ~n7084;
  assign n7086 = ~n7077 & n7085;
  assign n7110 = n7109 ^ n7086;
  assign n6861 = n6860 ^ n6855;
  assign n6846 = x580 ^ x579;
  assign n6848 = n6847 ^ n6846;
  assign n6845 = x582 ^ x581;
  assign n6849 = n6848 ^ n6845;
  assign n6841 = x574 ^ x573;
  assign n6843 = n6842 ^ n6841;
  assign n6840 = x576 ^ x575;
  assign n6844 = n6843 ^ n6840;
  assign n6850 = n6849 ^ n6844;
  assign n6862 = n6861 ^ n6850;
  assign n9397 = n6844 & n6849;
  assign n9406 = ~n6855 & ~n9397;
  assign n9407 = n6862 & n9406;
  assign n9408 = ~n6844 & ~n6849;
  assign n9409 = ~n9407 & ~n9408;
  assign n9410 = n9409 ^ n9397;
  assign n9411 = ~n7110 & ~n9410;
  assign n9412 = n9411 ^ n9397;
  assign n9413 = n9405 & n9412;
  assign n7059 = n6860 ^ n6844;
  assign n7061 = n7059 ^ n6855;
  assign n7062 = ~n6849 & n7061;
  assign n7060 = ~n6861 & ~n7059;
  assign n7063 = n7062 ^ n7060;
  assign n7111 = n7110 ^ n7063;
  assign n9414 = ~n7036 & n7057;
  assign n9415 = ~n7111 & n9414;
  assign n9416 = ~n9413 & ~n9415;
  assign n9398 = n7110 & n9397;
  assign n9399 = n7086 & n7109;
  assign n9400 = ~n9398 & ~n9399;
  assign n9395 = n7073 & ~n7082;
  assign n9394 = n7096 & ~n7105;
  assign n9396 = n9395 ^ n9394;
  assign n9401 = n9400 ^ n9396;
  assign n9557 = n9416 ^ n9401;
  assign n9417 = n7111 & n9403;
  assign n9418 = ~n9412 & n9417;
  assign n9558 = n7051 & ~n9418;
  assign n9559 = n9558 ^ n9401;
  assign n9560 = ~n9557 & ~n9559;
  assign n9561 = n9560 ^ n9416;
  assign n9554 = n9400 ^ n9395;
  assign n9555 = ~n9396 & n9554;
  assign n9556 = n9555 ^ n9400;
  assign n9562 = n9561 ^ n9556;
  assign n9563 = n7045 & n9396;
  assign n9564 = n9418 & n9563;
  assign n9565 = n9392 & ~n9564;
  assign n9566 = ~n9562 & n9565;
  assign n9419 = n9416 & ~n9418;
  assign n9567 = ~n9392 & n9556;
  assign n9568 = n9419 & n9567;
  assign n9569 = n9401 & ~n9416;
  assign n9570 = ~n9556 & n9569;
  assign n9571 = ~n9568 & ~n9570;
  assign n9572 = n7051 & ~n9571;
  assign n9573 = ~n9401 & n9416;
  assign n9574 = ~n9556 & ~n9573;
  assign n9576 = ~n9568 & n9575;
  assign n9577 = ~n9574 & n9576;
  assign n9578 = ~n9557 & n9567;
  assign n9579 = ~n9577 & ~n9578;
  assign n9580 = ~n9572 & n9579;
  assign n9581 = ~n9566 & n9580;
  assign n9911 = ~n9575 & ~n9581;
  assign n9912 = n9556 & ~n9573;
  assign n9913 = ~n9911 & ~n9912;
  assign n6890 = x605 & x606;
  assign n6891 = x603 & x604;
  assign n6892 = ~n6890 & ~n6891;
  assign n6893 = ~x605 & ~x606;
  assign n6894 = ~x603 & ~x604;
  assign n6895 = ~n6893 & ~n6894;
  assign n6896 = ~n6892 & n6895;
  assign n6897 = x602 & n6896;
  assign n6898 = n6890 & n6891;
  assign n6899 = ~n6897 & ~n6898;
  assign n6824 = x602 ^ x601;
  assign n6906 = n6824 & n6896;
  assign n6900 = n6892 & ~n6895;
  assign n6907 = x601 & x602;
  assign n6908 = n6891 & n6907;
  assign n6909 = x606 & n6908;
  assign n6910 = n6909 ^ n6907;
  assign n6911 = ~n6900 & n6910;
  assign n6912 = ~n6906 & ~n6911;
  assign n9368 = n6899 & n6912;
  assign n6919 = x599 & x600;
  assign n6920 = x597 & x598;
  assign n6921 = ~n6919 & ~n6920;
  assign n6922 = ~x599 & ~x600;
  assign n6923 = ~x597 & ~x598;
  assign n6924 = ~n6922 & ~n6923;
  assign n6925 = ~n6921 & n6924;
  assign n6926 = x596 & n6925;
  assign n6927 = n6919 & n6920;
  assign n6928 = ~n6926 & ~n6927;
  assign n6819 = x596 ^ x595;
  assign n6935 = n6819 & n6925;
  assign n6929 = n6921 & ~n6924;
  assign n6936 = x595 & x596;
  assign n6937 = n6920 & n6936;
  assign n6938 = x600 & n6937;
  assign n6939 = n6938 ^ n6936;
  assign n6940 = ~n6929 & n6939;
  assign n6941 = ~n6935 & ~n6940;
  assign n9367 = n6928 & n6941;
  assign n9369 = n9368 ^ n9367;
  assign n6930 = ~x596 & n6929;
  assign n6931 = n6922 & n6923;
  assign n6932 = ~n6930 & ~n6931;
  assign n6933 = n6928 & n6932;
  assign n6934 = ~x595 & ~n6933;
  assign n6942 = ~x596 & ~x600;
  assign n6943 = n6923 & n6942;
  assign n6944 = ~n6937 & ~n6943;
  assign n6945 = ~x599 & ~n6944;
  assign n6946 = n6941 & ~n6945;
  assign n6947 = ~n6934 & n6946;
  assign n6901 = ~x602 & n6900;
  assign n6902 = n6893 & n6894;
  assign n6903 = ~n6901 & ~n6902;
  assign n6904 = n6899 & n6903;
  assign n6905 = ~x601 & ~n6904;
  assign n6913 = ~x602 & ~x606;
  assign n6914 = n6894 & n6913;
  assign n6915 = ~n6908 & ~n6914;
  assign n6916 = ~x605 & ~n6915;
  assign n6917 = n6912 & ~n6916;
  assign n6918 = ~n6905 & n6917;
  assign n6948 = n6947 ^ n6918;
  assign n6818 = x598 ^ x597;
  assign n6820 = n6819 ^ n6818;
  assign n6817 = x600 ^ x599;
  assign n6821 = n6820 ^ n6817;
  assign n6823 = x604 ^ x603;
  assign n6825 = n6824 ^ n6823;
  assign n6822 = x606 ^ x605;
  assign n6826 = n6825 ^ n6822;
  assign n6875 = n6821 & n6826;
  assign n9364 = n6918 ^ n6875;
  assign n9365 = n6948 & ~n9364;
  assign n9366 = n9365 ^ n6947;
  assign n9370 = n9369 ^ n9366;
  assign n6830 = x586 ^ x585;
  assign n6829 = x588 ^ x587;
  assign n6831 = n6830 ^ n6829;
  assign n6828 = x584 ^ x583;
  assign n6832 = n6831 ^ n6828;
  assign n6835 = x590 ^ x589;
  assign n6834 = x592 ^ x591;
  assign n6836 = n6835 ^ n6834;
  assign n6833 = x594 ^ x593;
  assign n6837 = n6836 ^ n6833;
  assign n6878 = n6832 & n6837;
  assign n6980 = ~x585 & ~x586;
  assign n6981 = ~x587 & ~x588;
  assign n6982 = ~n6980 & ~n6981;
  assign n6983 = x585 & x586;
  assign n6984 = x587 & x588;
  assign n6985 = ~n6983 & ~n6984;
  assign n6986 = n6982 & ~n6985;
  assign n6987 = x584 & n6986;
  assign n6988 = n6983 & n6984;
  assign n6989 = ~n6987 & ~n6988;
  assign n6990 = ~n6982 & n6985;
  assign n6991 = ~x584 & n6990;
  assign n6992 = n6980 & n6981;
  assign n6993 = ~n6991 & ~n6992;
  assign n6994 = n6989 & n6993;
  assign n6995 = ~x583 & ~n6994;
  assign n6996 = ~x584 & n6986;
  assign n6997 = x588 & n6983;
  assign n6998 = x584 & ~n6997;
  assign n6999 = ~n6990 & n6998;
  assign n7000 = ~n6996 & ~n6999;
  assign n7001 = x583 & ~n7000;
  assign n7002 = x583 & x584;
  assign n7003 = n6983 & n7002;
  assign n7004 = ~x584 & ~x588;
  assign n7005 = n6980 & n7004;
  assign n7006 = ~n7003 & ~n7005;
  assign n7007 = ~x587 & ~n7006;
  assign n7008 = ~n7001 & ~n7007;
  assign n7009 = ~n6995 & n7008;
  assign n6950 = x591 & x592;
  assign n6951 = x593 & x594;
  assign n6952 = ~n6950 & ~n6951;
  assign n6953 = ~x591 & ~x592;
  assign n6954 = ~x593 & ~x594;
  assign n6955 = ~n6953 & ~n6954;
  assign n6956 = ~n6952 & n6955;
  assign n6957 = x590 & n6956;
  assign n6958 = n6950 & n6951;
  assign n6959 = ~n6957 & ~n6958;
  assign n6960 = x590 & ~n6954;
  assign n6961 = ~n6951 & n6953;
  assign n6962 = ~n6960 & n6961;
  assign n6963 = n6959 & ~n6962;
  assign n6964 = ~x589 & ~n6963;
  assign n6965 = ~x590 & ~x594;
  assign n6966 = ~n6950 & n6965;
  assign n6967 = n6836 & n6966;
  assign n6968 = x589 & x590;
  assign n6969 = n6950 & n6968;
  assign n6970 = ~n6967 & ~n6969;
  assign n6971 = ~x593 & ~n6970;
  assign n6972 = n6952 & ~n6955;
  assign n6973 = x594 & n6969;
  assign n6974 = n6973 ^ n6968;
  assign n6975 = ~n6972 & n6974;
  assign n6976 = n6835 & n6956;
  assign n6977 = ~n6975 & ~n6976;
  assign n6978 = ~n6971 & n6977;
  assign n6979 = ~n6964 & n6978;
  assign n7010 = n7009 ^ n6979;
  assign n9379 = ~n6878 & ~n7010;
  assign n6827 = n6826 ^ n6821;
  assign n6838 = n6837 ^ n6832;
  assign n9380 = n6838 ^ n6821;
  assign n9381 = n6827 & ~n9380;
  assign n9382 = n9381 ^ n6826;
  assign n9383 = ~n6948 & n9382;
  assign n9384 = ~n9379 & n9383;
  assign n9385 = ~n6875 & n6948;
  assign n9386 = ~n9384 & ~n9385;
  assign n6876 = ~n6832 & ~n6837;
  assign n6877 = ~n6875 & n6876;
  assign n6879 = ~n6821 & ~n6826;
  assign n6880 = ~n6878 & n6879;
  assign n6881 = ~n6877 & ~n6880;
  assign n9387 = n6881 ^ n6878;
  assign n9388 = ~n7010 & ~n9387;
  assign n9389 = n9388 ^ n6878;
  assign n9390 = ~n9386 & ~n9389;
  assign n9540 = ~n9370 & ~n9390;
  assign n9372 = n6989 & ~n7001;
  assign n9371 = n6959 & n6977;
  assign n9373 = n9372 ^ n9371;
  assign n9374 = ~n6878 & n7010;
  assign n9375 = ~n6979 & ~n7009;
  assign n9376 = ~n9374 & ~n9375;
  assign n9541 = n9376 ^ n9372;
  assign n9542 = ~n9373 & ~n9541;
  assign n9543 = n9542 ^ n9376;
  assign n9544 = n9540 & ~n9543;
  assign n9377 = n9376 ^ n9373;
  assign n9378 = n9377 ^ n9370;
  assign n9391 = n9390 ^ n9378;
  assign n9545 = n9371 & n9372;
  assign n9546 = ~n9376 & n9545;
  assign n9547 = n9391 & n9546;
  assign n9548 = ~n9544 & ~n9547;
  assign n9549 = n9370 & n9543;
  assign n9550 = ~n9391 & n9549;
  assign n9551 = n9548 & ~n9550;
  assign n9537 = n9368 ^ n9366;
  assign n9538 = ~n9369 & ~n9537;
  assign n9539 = n9538 ^ n9366;
  assign n9552 = n9551 ^ n9539;
  assign n9393 = n9392 ^ n7051;
  assign n9402 = n9401 ^ n9393;
  assign n9420 = n9419 ^ n9402;
  assign n9421 = n9420 ^ n9391;
  assign n6882 = ~n6862 & ~n6881;
  assign n6883 = ~n6878 & ~n6879;
  assign n6884 = ~n6875 & ~n6876;
  assign n6885 = ~n6883 & ~n6884;
  assign n6886 = ~n6882 & ~n6885;
  assign n6839 = n6838 ^ n6827;
  assign n6887 = n6839 & n6862;
  assign n6888 = n6881 & n6887;
  assign n6889 = n6886 & ~n6888;
  assign n6949 = n6948 ^ n6889;
  assign n7011 = n7010 ^ n6949;
  assign n7058 = n7057 ^ n7036;
  assign n7112 = n7111 ^ n7058;
  assign n9361 = n7112 ^ n6887;
  assign n9362 = ~n7011 & n9361;
  assign n9363 = n9362 ^ n7112;
  assign n9534 = n9391 ^ n9363;
  assign n9535 = ~n9421 & ~n9534;
  assign n9536 = n9535 ^ n9420;
  assign n9553 = n9552 ^ n9536;
  assign n9914 = n9581 ^ n9536;
  assign n9915 = n9553 & n9914;
  assign n9916 = n9915 ^ n9581;
  assign n9917 = ~n9913 & n9916;
  assign n9918 = n9536 & n9581;
  assign n9919 = n9552 & ~n9918;
  assign n9920 = n9913 & n9919;
  assign n9921 = ~n9917 & ~n9920;
  assign n9909 = ~n9539 & ~n9550;
  assign n9910 = n9548 & ~n9909;
  assign n9922 = n9921 ^ n9910;
  assign n10042 = ~n9908 & ~n9922;
  assign n9901 = ~n9508 & ~n9512;
  assign n9902 = ~n9495 & ~n9506;
  assign n9903 = ~n9901 & ~n9902;
  assign n9899 = ~n9518 & ~n9523;
  assign n9900 = ~n9528 & ~n9899;
  assign n9904 = n9903 ^ n9900;
  assign n9532 = n9531 ^ n9512;
  assign n9480 = n9479 ^ n9452;
  assign n9422 = n9421 ^ n9363;
  assign n9489 = n9480 ^ n9422;
  assign n6816 = n6815 ^ n6792;
  assign n6863 = n6862 ^ n6839;
  assign n6864 = n6863 ^ n6792;
  assign n6865 = n6816 & ~n6864;
  assign n6866 = n6865 ^ n6815;
  assign n7113 = n7112 ^ n7011;
  assign n9355 = n7113 & n7347;
  assign n9356 = ~n6866 & ~n9355;
  assign n9357 = n6871 & n7347;
  assign n9358 = ~n7113 & ~n7347;
  assign n9359 = ~n9357 & ~n9358;
  assign n9360 = ~n9356 & n9359;
  assign n9490 = n9480 ^ n9360;
  assign n9491 = ~n9489 & ~n9490;
  assign n9492 = n9491 ^ n9422;
  assign n9533 = n9532 ^ n9492;
  assign n9582 = n9581 ^ n9553;
  assign n9896 = n9582 ^ n9492;
  assign n9897 = n9533 & n9896;
  assign n9898 = n9897 ^ n9532;
  assign n10043 = n9903 ^ n9898;
  assign n10044 = ~n9904 & ~n10043;
  assign n10045 = n10044 ^ n9898;
  assign n10046 = n10042 & n10045;
  assign n10047 = ~n9900 & ~n9903;
  assign n10048 = n9898 & n10047;
  assign n9923 = n9922 ^ n9908;
  assign n9905 = n9904 ^ n9898;
  assign n9924 = n9923 ^ n9905;
  assign n10049 = n9898 & ~n9908;
  assign n10050 = n9924 & ~n10049;
  assign n10051 = n10048 & ~n10050;
  assign n10052 = ~n10046 & ~n10051;
  assign n10053 = n9922 & ~n10045;
  assign n10054 = n9924 & n10053;
  assign n10055 = n10052 & ~n10054;
  assign n10040 = ~n9910 & ~n9920;
  assign n10041 = ~n9917 & ~n10040;
  assign n10056 = n10055 ^ n10041;
  assign n7754 = x515 & x516;
  assign n7755 = x513 & x514;
  assign n7756 = ~n7754 & ~n7755;
  assign n7757 = ~x515 & ~x516;
  assign n7758 = ~x513 & ~x514;
  assign n7759 = ~n7757 & ~n7758;
  assign n7760 = ~n7756 & n7759;
  assign n7761 = x512 & n7760;
  assign n7762 = n7754 & n7755;
  assign n7763 = ~n7761 & ~n7762;
  assign n7764 = n7756 & ~n7759;
  assign n7768 = ~n7762 & ~n7764;
  assign n7769 = x512 & ~n7768;
  assign n7770 = ~x512 & ~n7760;
  assign n7771 = x511 & ~n7770;
  assign n7772 = ~n7769 & n7771;
  assign n9306 = n7763 & ~n7772;
  assign n7731 = x521 & x522;
  assign n7732 = x519 & x520;
  assign n7733 = ~n7731 & ~n7732;
  assign n7734 = ~x521 & ~x522;
  assign n7735 = ~x519 & ~x520;
  assign n7736 = ~n7734 & ~n7735;
  assign n7737 = ~n7733 & n7736;
  assign n7738 = x518 & n7737;
  assign n7739 = n7731 & n7732;
  assign n7740 = ~n7738 & ~n7739;
  assign n7741 = n7733 & ~n7736;
  assign n7745 = ~n7739 & ~n7741;
  assign n7746 = x518 & ~n7745;
  assign n7747 = ~x518 & ~n7737;
  assign n7748 = x517 & ~n7747;
  assign n7749 = ~n7746 & n7748;
  assign n9307 = n7740 & ~n7749;
  assign n9647 = ~n9306 & ~n9307;
  assign n7699 = x527 & x528;
  assign n7700 = x525 & x526;
  assign n7701 = ~n7699 & ~n7700;
  assign n7702 = ~x527 & ~x528;
  assign n7703 = ~x525 & ~x526;
  assign n7704 = ~n7702 & ~n7703;
  assign n7705 = ~n7701 & n7704;
  assign n7706 = x524 & n7705;
  assign n7707 = n7699 & n7700;
  assign n7708 = ~n7706 & ~n7707;
  assign n7709 = n7701 & ~n7704;
  assign n7713 = ~n7707 & ~n7709;
  assign n7714 = x524 & ~n7713;
  assign n7715 = ~x524 & ~n7705;
  assign n7716 = x523 & ~n7715;
  assign n7717 = ~n7714 & n7716;
  assign n9314 = n7708 & ~n7717;
  assign n7676 = x531 & x532;
  assign n7677 = x533 & x534;
  assign n7678 = ~n7676 & ~n7677;
  assign n7679 = ~x531 & ~x532;
  assign n7680 = ~x533 & ~x534;
  assign n7681 = ~n7679 & ~n7680;
  assign n7682 = ~n7678 & n7681;
  assign n7683 = x530 & n7682;
  assign n7684 = n7676 & n7677;
  assign n7685 = ~n7683 & ~n7684;
  assign n7686 = n7678 & ~n7681;
  assign n7690 = ~n7684 & ~n7686;
  assign n7691 = x530 & ~n7690;
  assign n7692 = ~x530 & ~n7682;
  assign n7693 = x529 & ~n7692;
  assign n7694 = ~n7691 & n7693;
  assign n9313 = n7685 & ~n7694;
  assign n9315 = n9314 ^ n9313;
  assign n7710 = ~x524 & n7709;
  assign n7711 = n7708 & ~n7710;
  assign n7712 = ~x523 & ~n7711;
  assign n6758 = x524 ^ x523;
  assign n7718 = n7702 & n7703;
  assign n7719 = n6758 & n7718;
  assign n7720 = ~n7717 & ~n7719;
  assign n7721 = ~n7712 & n7720;
  assign n7687 = ~x530 & n7686;
  assign n7688 = n7685 & ~n7687;
  assign n7689 = ~x529 & ~n7688;
  assign n6763 = x530 ^ x529;
  assign n7695 = n7679 & n7680;
  assign n7696 = n6763 & n7695;
  assign n7697 = ~n7694 & ~n7696;
  assign n7698 = ~n7689 & n7697;
  assign n7722 = n7721 ^ n7698;
  assign n6757 = x526 ^ x525;
  assign n6759 = n6758 ^ n6757;
  assign n6756 = x528 ^ x527;
  assign n6760 = n6759 ^ n6756;
  assign n6762 = x532 ^ x531;
  assign n6764 = n6763 ^ n6762;
  assign n6761 = x534 ^ x533;
  assign n6765 = n6764 ^ n6761;
  assign n7723 = n6760 & n6765;
  assign n9310 = n7723 ^ n7721;
  assign n9311 = ~n7722 & n9310;
  assign n9312 = n9311 ^ n7723;
  assign n9316 = n9315 ^ n9312;
  assign n7765 = ~x512 & n7764;
  assign n7766 = n7763 & ~n7765;
  assign n7767 = ~x511 & ~n7766;
  assign n6747 = x512 ^ x511;
  assign n7773 = n7757 & n7758;
  assign n7774 = n6747 & n7773;
  assign n7775 = ~n7772 & ~n7774;
  assign n7776 = ~n7767 & n7775;
  assign n7742 = ~x518 & n7741;
  assign n7743 = n7740 & ~n7742;
  assign n7744 = ~x517 & ~n7743;
  assign n6752 = x518 ^ x517;
  assign n7750 = n7734 & n7735;
  assign n7751 = n6752 & n7750;
  assign n7752 = ~n7749 & ~n7751;
  assign n7753 = ~n7744 & n7752;
  assign n7777 = n7776 ^ n7753;
  assign n6746 = x514 ^ x513;
  assign n6748 = n6747 ^ n6746;
  assign n6745 = x516 ^ x515;
  assign n6749 = n6748 ^ n6745;
  assign n6751 = x520 ^ x519;
  assign n6753 = n6752 ^ n6751;
  assign n6750 = x522 ^ x521;
  assign n6754 = n6753 ^ n6750;
  assign n7727 = n6749 & n6754;
  assign n9303 = n7753 ^ n7727;
  assign n9304 = n7777 & ~n9303;
  assign n9305 = n9304 ^ n7776;
  assign n6755 = n6754 ^ n6749;
  assign n6766 = n6765 ^ n6760;
  assign n7724 = n6766 ^ n6754;
  assign n7725 = ~n6755 & n7724;
  assign n7726 = n7725 ^ n6766;
  assign n7728 = n7727 ^ n7726;
  assign n7729 = ~n7723 & ~n7728;
  assign n7730 = n7729 ^ n7727;
  assign n7778 = n7777 ^ n7730;
  assign n9318 = ~n7722 & ~n7778;
  assign n9319 = n7722 & n7723;
  assign n9320 = n7727 & n7777;
  assign n9321 = ~n9319 & ~n9320;
  assign n9322 = ~n9318 & n9321;
  assign n9323 = ~n7726 & ~n7777;
  assign n9324 = n9322 & ~n9323;
  assign n9637 = ~n9305 & ~n9324;
  assign n9638 = n9316 & ~n9637;
  assign n9639 = n9305 & n9324;
  assign n9640 = n9306 & n9307;
  assign n9641 = ~n9639 & n9640;
  assign n9642 = ~n9638 & n9641;
  assign n9643 = n9316 & ~n9640;
  assign n9644 = n9639 & n9643;
  assign n9645 = ~n9642 & ~n9644;
  assign n9646 = n9637 ^ n9316;
  assign n9648 = n9647 ^ n9316;
  assign n9649 = n9646 & ~n9648;
  assign n9650 = n9645 & ~n9649;
  assign n9634 = n9314 ^ n9312;
  assign n9635 = ~n9315 & ~n9634;
  assign n9636 = n9635 ^ n9312;
  assign n9651 = n9650 ^ n9636;
  assign n9872 = ~n9647 & n9651;
  assign n9873 = ~n9636 & ~n9638;
  assign n9874 = ~n9872 & ~n9873;
  assign n7660 = x551 & x552;
  assign n7661 = x549 & x550;
  assign n7662 = n7660 & n7661;
  assign n7651 = ~x551 & ~x552;
  assign n7652 = ~x550 & n7651;
  assign n7653 = x549 & ~n7652;
  assign n6738 = x552 ^ x551;
  assign n7654 = x551 ^ x550;
  assign n7655 = ~n6738 & n7654;
  assign n7656 = n7655 ^ x550;
  assign n7657 = ~n7653 & ~n7656;
  assign n7665 = x547 & x548;
  assign n7667 = ~n7662 & n7665;
  assign n7668 = ~n7657 & n7667;
  assign n6739 = x550 ^ x549;
  assign n6740 = n6739 ^ n6738;
  assign n6741 = x548 ^ x547;
  assign n7669 = n6740 & n6741;
  assign n7670 = n7656 & n7669;
  assign n7671 = ~n7668 & ~n7670;
  assign n9334 = ~n7662 & n7671;
  assign n6734 = x556 ^ x555;
  assign n7628 = x557 & x558;
  assign n7629 = n7628 ^ x556;
  assign n7630 = ~n6734 & ~n7629;
  assign n7632 = x555 & x556;
  assign n7633 = ~x557 & ~x558;
  assign n7634 = ~n7632 & n7633;
  assign n7642 = x553 & x554;
  assign n7643 = ~n7634 & n7642;
  assign n7644 = ~n7630 & n7643;
  assign n6735 = x554 ^ x553;
  assign n7637 = ~x555 & ~x556;
  assign n7645 = n7628 & ~n7637;
  assign n7646 = n7632 & ~n7633;
  assign n7647 = ~n7645 & ~n7646;
  assign n7648 = n6735 & ~n7647;
  assign n7649 = ~n7644 & ~n7648;
  assign n9332 = n7628 & n7632;
  assign n9333 = n7649 & ~n9332;
  assign n9335 = n9334 ^ n9333;
  assign n6736 = n6735 ^ n6734;
  assign n6733 = x558 ^ x557;
  assign n6737 = n6736 ^ n6733;
  assign n6742 = n6741 ^ n6740;
  assign n7619 = n6737 & n6742;
  assign n7658 = ~n6741 & n7657;
  assign n7659 = ~x549 & n7652;
  assign n7663 = ~n7659 & ~n7662;
  assign n7664 = ~n7658 & n7663;
  assign n7666 = ~n7664 & ~n7665;
  assign n7672 = ~n7666 & n7671;
  assign n7631 = ~x553 & n7630;
  assign n7635 = ~x554 & n7634;
  assign n7636 = ~n7631 & ~n7635;
  assign n7638 = x553 & ~n7637;
  assign n7639 = x554 & ~n7633;
  assign n7640 = ~n7638 & ~n7639;
  assign n7641 = ~n7636 & n7640;
  assign n7650 = ~n7641 & n7649;
  assign n7673 = n7672 ^ n7650;
  assign n9336 = ~n7619 & n7673;
  assign n9337 = ~n7650 & ~n7672;
  assign n9338 = ~n9336 & ~n9337;
  assign n9653 = n9338 ^ n9334;
  assign n9654 = ~n9335 & ~n9653;
  assign n9655 = n9654 ^ n9338;
  assign n7590 = ~x545 & ~x546;
  assign n7591 = x541 & ~n7590;
  assign n6728 = x544 ^ x543;
  assign n7592 = x545 & x546;
  assign n7593 = n7592 ^ x544;
  assign n7594 = n6728 & ~n7593;
  assign n7595 = n7594 ^ x543;
  assign n7596 = n7591 & n7595;
  assign n7597 = x541 & x542;
  assign n7598 = ~n7596 & ~n7597;
  assign n7599 = x543 & x544;
  assign n7600 = n7590 & ~n7599;
  assign n7601 = ~x543 & ~x544;
  assign n7602 = ~n7592 & n7601;
  assign n7603 = ~n7600 & ~n7602;
  assign n7604 = n7592 & n7599;
  assign n7605 = n7603 & ~n7604;
  assign n7606 = x542 & ~n7605;
  assign n7607 = ~n7598 & ~n7606;
  assign n7608 = x542 & ~n7590;
  assign n7609 = ~n7604 & ~n7608;
  assign n7610 = n7595 & ~n7609;
  assign n7611 = n7602 & ~n7608;
  assign n7612 = ~n7610 & ~n7611;
  assign n7613 = ~x541 & ~n7612;
  assign n7614 = ~n7607 & ~n7613;
  assign n6729 = x546 ^ x545;
  assign n6730 = n6729 ^ n6728;
  assign n6727 = x542 ^ x541;
  assign n6731 = n6730 ^ n6727;
  assign n7615 = ~x542 & n7600;
  assign n7616 = n6731 & n7615;
  assign n7617 = n7614 & ~n7616;
  assign n7567 = x539 & x540;
  assign n7568 = x537 & x538;
  assign n7569 = ~n7567 & ~n7568;
  assign n7570 = ~x539 & ~x540;
  assign n7571 = ~x537 & ~x538;
  assign n7572 = ~n7570 & ~n7571;
  assign n7573 = ~n7569 & n7572;
  assign n7574 = x536 & n7573;
  assign n7575 = n7567 & n7568;
  assign n7576 = ~n7574 & ~n7575;
  assign n7577 = n7569 & ~n7572;
  assign n7578 = ~x536 & n7577;
  assign n7579 = n7576 & ~n7578;
  assign n7580 = ~x535 & ~n7579;
  assign n7581 = ~n7575 & ~n7577;
  assign n7582 = x536 & ~n7581;
  assign n7583 = ~x536 & ~n7573;
  assign n7584 = x535 & ~n7583;
  assign n7585 = ~n7582 & n7584;
  assign n6724 = x536 ^ x535;
  assign n7586 = n7570 & n7571;
  assign n7587 = n6724 & n7586;
  assign n7588 = ~n7585 & ~n7587;
  assign n7589 = ~n7580 & n7588;
  assign n7618 = n7617 ^ n7589;
  assign n6723 = x538 ^ x537;
  assign n6725 = n6724 ^ n6723;
  assign n6722 = x540 ^ x539;
  assign n6726 = n6725 ^ n6722;
  assign n7620 = ~n6726 & ~n6731;
  assign n7621 = ~n7619 & n7620;
  assign n7622 = n6726 & n6731;
  assign n7623 = ~n6737 & ~n6742;
  assign n7624 = ~n7622 & n7623;
  assign n7625 = ~n7621 & ~n7624;
  assign n7626 = n7619 & n7622;
  assign n7627 = n7625 & ~n7626;
  assign n7674 = n7673 ^ n7627;
  assign n9341 = ~n7618 & n7674;
  assign n9342 = n7625 ^ n7619;
  assign n9343 = ~n7673 & ~n9342;
  assign n9344 = n9343 ^ n7619;
  assign n9345 = ~n9341 & ~n9344;
  assign n9346 = n7618 & n7622;
  assign n9347 = n9345 & ~n9346;
  assign n9326 = n7576 & ~n7585;
  assign n9327 = ~n7607 & ~n7610;
  assign n9656 = ~n9326 & ~n9327;
  assign n9657 = ~n9347 & ~n9656;
  assign n9329 = n7622 ^ n7617;
  assign n9330 = ~n7618 & n9329;
  assign n9331 = n9330 ^ n7622;
  assign n9339 = n9338 ^ n9335;
  assign n9658 = n9331 & n9339;
  assign n9659 = ~n9657 & n9658;
  assign n9660 = ~n9331 & ~n9339;
  assign n9661 = n9347 & ~n9660;
  assign n9662 = n9656 & n9661;
  assign n9663 = ~n9659 & ~n9662;
  assign n9664 = ~n9655 & n9663;
  assign n9340 = n9339 ^ n9331;
  assign n9348 = n9347 ^ n9340;
  assign n9665 = n9326 & n9327;
  assign n9666 = n9348 & n9665;
  assign n9667 = n9657 & n9660;
  assign n9668 = ~n9666 & ~n9667;
  assign n9669 = ~n9664 & n9668;
  assign n9875 = n9874 ^ n9669;
  assign n9328 = n9327 ^ n9326;
  assign n9349 = n9348 ^ n9328;
  assign n9308 = n9307 ^ n9306;
  assign n9309 = n9308 ^ n9305;
  assign n9317 = n9316 ^ n9309;
  assign n9325 = n9324 ^ n9317;
  assign n9350 = n9349 ^ n9325;
  assign n7779 = n7778 ^ n7722;
  assign n7675 = n7674 ^ n7618;
  assign n7780 = n7779 ^ n7675;
  assign n6743 = n6742 ^ n6737;
  assign n6732 = n6731 ^ n6726;
  assign n6744 = n6743 ^ n6732;
  assign n6767 = n6766 ^ n6755;
  assign n9296 = n6744 & n6767;
  assign n9300 = n9296 ^ n7675;
  assign n9301 = ~n7780 & ~n9300;
  assign n9302 = n9301 ^ n7779;
  assign n9631 = n9325 ^ n9302;
  assign n9632 = n9350 & n9631;
  assign n9633 = n9632 ^ n9349;
  assign n9652 = n9651 ^ n9633;
  assign n9670 = n9339 & n9347;
  assign n9671 = n9669 & n9670;
  assign n9672 = ~n9661 & n9666;
  assign n9673 = n9656 & n9658;
  assign n9674 = ~n9667 & ~n9673;
  assign n9675 = ~n9672 & n9674;
  assign n9676 = ~n9671 & n9675;
  assign n9677 = n9676 ^ n9655;
  assign n9869 = n9677 ^ n9651;
  assign n9870 = ~n9652 & n9869;
  assign n9871 = n9870 ^ n9677;
  assign n9876 = n9875 ^ n9871;
  assign n7401 = x501 & x502;
  assign n7402 = x503 & x504;
  assign n7403 = ~n7401 & ~n7402;
  assign n7404 = ~x501 & ~x502;
  assign n7405 = ~x503 & ~x504;
  assign n7406 = ~n7404 & ~n7405;
  assign n7407 = ~n7403 & n7406;
  assign n7408 = x500 & n7407;
  assign n7409 = n7401 & n7402;
  assign n7410 = ~n7408 & ~n7409;
  assign n7411 = n7403 & ~n7406;
  assign n7415 = ~n7409 & ~n7411;
  assign n7416 = x500 & ~n7415;
  assign n7417 = ~x500 & ~n7407;
  assign n7418 = x499 & ~n7417;
  assign n7419 = ~n7416 & n7418;
  assign n9276 = n7410 & ~n7419;
  assign n7432 = x509 & x510;
  assign n7433 = x508 & n7432;
  assign n7434 = x507 & n7433;
  assign n7424 = ~x509 & ~x510;
  assign n7425 = ~x508 & n7424;
  assign n7426 = x507 & ~n7425;
  assign n6703 = x510 ^ x509;
  assign n7427 = x509 ^ x508;
  assign n7428 = ~n6703 & n7427;
  assign n7429 = n7428 ^ x508;
  assign n7430 = ~n7426 & ~n7429;
  assign n7437 = x505 & x506;
  assign n7438 = ~n7434 & n7437;
  assign n7439 = ~n7430 & n7438;
  assign n6705 = x506 ^ x505;
  assign n7440 = ~x507 & ~n7433;
  assign n7441 = n6705 & ~n7440;
  assign n7442 = n7429 & n7441;
  assign n7443 = ~n7439 & ~n7442;
  assign n9275 = ~n7434 & n7443;
  assign n9277 = n9276 ^ n9275;
  assign n7431 = ~x506 & n7430;
  assign n7435 = ~n7431 & ~n7434;
  assign n7436 = ~x505 & ~n7435;
  assign n7444 = ~x507 & ~n7437;
  assign n7445 = n7425 & n7444;
  assign n7446 = n7443 & ~n7445;
  assign n7447 = ~n7436 & n7446;
  assign n7412 = ~x500 & n7411;
  assign n7413 = n7410 & ~n7412;
  assign n7414 = ~x499 & ~n7413;
  assign n6700 = x500 ^ x499;
  assign n7420 = n7404 & n7405;
  assign n7421 = n6700 & n7420;
  assign n7422 = ~n7419 & ~n7421;
  assign n7423 = ~n7414 & n7422;
  assign n7448 = n7447 ^ n7423;
  assign n6699 = x502 ^ x501;
  assign n6701 = n6700 ^ n6699;
  assign n6698 = x504 ^ x503;
  assign n6702 = n6701 ^ n6698;
  assign n6704 = x508 ^ x507;
  assign n6706 = n6705 ^ n6704;
  assign n6707 = n6706 ^ n6703;
  assign n7358 = n6702 & n6707;
  assign n9272 = n7423 ^ n7358;
  assign n9273 = n7448 & ~n9272;
  assign n9274 = n9273 ^ n7447;
  assign n9278 = n9277 ^ n9274;
  assign n6711 = x494 ^ x493;
  assign n7379 = x495 & x496;
  assign n7380 = x497 & x498;
  assign n7381 = ~n7379 & ~n7380;
  assign n7382 = ~x495 & ~x496;
  assign n7383 = ~x497 & ~x498;
  assign n7384 = ~n7382 & ~n7383;
  assign n7385 = n7381 & ~n7384;
  assign n7386 = ~n6711 & n7385;
  assign n7387 = n7379 & n7380;
  assign n7388 = n7382 & n7383;
  assign n7389 = ~n7387 & ~n7388;
  assign n7390 = ~n7386 & n7389;
  assign n7391 = x493 & x494;
  assign n7392 = ~n7390 & ~n7391;
  assign n7393 = n6711 & n7384;
  assign n7394 = ~n7381 & n7393;
  assign n7395 = ~n7387 & n7391;
  assign n7396 = ~n7385 & n7395;
  assign n7397 = ~n7394 & ~n7396;
  assign n7398 = ~n7392 & n7397;
  assign n6717 = x488 ^ x487;
  assign n7360 = x489 & x490;
  assign n7361 = ~x491 & ~x492;
  assign n7362 = ~n7360 & n7361;
  assign n7363 = ~x489 & ~x490;
  assign n7364 = x491 & x492;
  assign n7365 = n7363 & ~n7364;
  assign n7366 = ~n7362 & ~n7365;
  assign n7367 = ~n6717 & ~n7366;
  assign n7368 = n7360 & n7364;
  assign n7369 = n7361 & n7363;
  assign n7370 = ~n7368 & ~n7369;
  assign n7371 = ~n7367 & n7370;
  assign n7372 = x487 & x488;
  assign n7373 = ~n7371 & ~n7372;
  assign n6715 = x490 ^ x489;
  assign n6714 = x492 ^ x491;
  assign n6716 = n6715 ^ n6714;
  assign n7374 = n6716 & n6717;
  assign n7375 = ~n7368 & n7372;
  assign n7376 = ~n7374 & ~n7375;
  assign n7377 = n7366 & ~n7376;
  assign n7378 = ~n7373 & ~n7377;
  assign n7399 = n7398 ^ n7378;
  assign n6718 = n6717 ^ n6716;
  assign n6710 = x496 ^ x495;
  assign n6712 = n6711 ^ n6710;
  assign n6709 = x498 ^ x497;
  assign n6713 = n6712 ^ n6709;
  assign n6719 = n6718 ^ n6713;
  assign n6708 = n6707 ^ n6702;
  assign n7355 = n6713 ^ n6708;
  assign n7356 = n6719 & ~n7355;
  assign n7357 = n7356 ^ n6718;
  assign n7359 = n7358 ^ n7357;
  assign n7400 = n7399 ^ n7359;
  assign n9281 = n7400 & ~n7448;
  assign n9267 = n6713 & n6718;
  assign n9282 = n9267 ^ n7357;
  assign n9283 = n7399 & ~n9282;
  assign n9284 = n9283 ^ n7357;
  assign n9285 = ~n9281 & n9284;
  assign n9286 = n7358 & n7448;
  assign n9287 = n9285 & ~n9286;
  assign n9280 = ~n7387 & n7397;
  assign n9288 = n9287 ^ n9280;
  assign n9268 = n7399 & n9267;
  assign n9269 = n7378 & n7398;
  assign n9270 = ~n9268 & ~n9269;
  assign n9266 = ~n7368 & ~n7377;
  assign n9271 = n9270 ^ n9266;
  assign n9279 = n9278 ^ n9271;
  assign n9289 = n9288 ^ n9279;
  assign n9615 = n9278 & n9289;
  assign n9616 = ~n9266 & ~n9270;
  assign n9617 = ~n9615 & ~n9616;
  assign n9618 = n9280 & ~n9287;
  assign n9619 = n9617 & n9618;
  assign n9620 = ~n9280 & n9287;
  assign n9621 = ~n9616 & ~n9620;
  assign n9622 = n9615 & ~n9621;
  assign n9623 = n9270 & ~n9278;
  assign n9624 = n9266 & n9623;
  assign n9625 = ~n9620 & n9624;
  assign n9626 = ~n9622 & ~n9625;
  assign n9627 = ~n9619 & n9626;
  assign n9612 = n9276 ^ n9274;
  assign n9613 = ~n9277 & ~n9612;
  assign n9614 = n9613 ^ n9274;
  assign n9628 = n9627 ^ n9614;
  assign n7510 = x479 & x480;
  assign n7511 = x477 & x478;
  assign n7512 = ~n7510 & ~n7511;
  assign n7513 = ~x479 & ~x480;
  assign n7514 = ~x477 & ~x478;
  assign n7515 = ~n7513 & ~n7514;
  assign n7516 = ~n7512 & n7515;
  assign n7517 = x476 & n7516;
  assign n7518 = n7510 & n7511;
  assign n7519 = ~n7517 & ~n7518;
  assign n7520 = n7512 & ~n7515;
  assign n7524 = ~n7518 & ~n7520;
  assign n7525 = x476 & ~n7524;
  assign n7526 = ~x476 & ~n7516;
  assign n7527 = x475 & ~n7526;
  assign n7528 = ~n7525 & n7527;
  assign n9254 = n7519 & ~n7528;
  assign n7533 = x485 & x486;
  assign n7534 = x483 & x484;
  assign n7535 = ~n7533 & ~n7534;
  assign n7536 = ~x485 & ~x486;
  assign n7537 = ~x483 & ~x484;
  assign n7538 = ~n7536 & ~n7537;
  assign n7539 = ~n7535 & n7538;
  assign n7540 = x482 & n7539;
  assign n7541 = n7533 & n7534;
  assign n7542 = ~n7540 & ~n7541;
  assign n6682 = x482 ^ x481;
  assign n7549 = n6682 & n7539;
  assign n7543 = n7535 & ~n7538;
  assign n7550 = x481 & x482;
  assign n7551 = n7534 & n7550;
  assign n7552 = x486 & n7551;
  assign n7553 = n7552 ^ n7550;
  assign n7554 = ~n7543 & n7553;
  assign n7555 = ~n7549 & ~n7554;
  assign n9253 = n7542 & n7555;
  assign n9255 = n9254 ^ n9253;
  assign n7544 = ~x482 & n7543;
  assign n7545 = n7536 & n7537;
  assign n7546 = ~n7544 & ~n7545;
  assign n7547 = n7542 & n7546;
  assign n7548 = ~x481 & ~n7547;
  assign n7556 = ~x482 & ~x486;
  assign n7557 = n7537 & n7556;
  assign n7558 = ~n7551 & ~n7557;
  assign n7559 = ~x485 & ~n7558;
  assign n7560 = n7555 & ~n7559;
  assign n7561 = ~n7548 & n7560;
  assign n7521 = ~x476 & n7520;
  assign n7522 = n7519 & ~n7521;
  assign n7523 = ~x475 & ~n7522;
  assign n6677 = x476 ^ x475;
  assign n7529 = n7513 & n7514;
  assign n7530 = n6677 & n7529;
  assign n7531 = ~n7528 & ~n7530;
  assign n7532 = ~n7523 & n7531;
  assign n7562 = n7561 ^ n7532;
  assign n6676 = x478 ^ x477;
  assign n6678 = n6677 ^ n6676;
  assign n6675 = x480 ^ x479;
  assign n6679 = n6678 ^ n6675;
  assign n6681 = x484 ^ x483;
  assign n6683 = n6682 ^ n6681;
  assign n6680 = x486 ^ x485;
  assign n6684 = n6683 ^ n6680;
  assign n7506 = n6679 & n6684;
  assign n9250 = n7532 ^ n7506;
  assign n9251 = n7562 & ~n9250;
  assign n9252 = n9251 ^ n7561;
  assign n9256 = n9255 ^ n9252;
  assign n7478 = x467 & x468;
  assign n7479 = x465 & x466;
  assign n7480 = ~n7478 & ~n7479;
  assign n7481 = ~x467 & ~x468;
  assign n7482 = ~x465 & ~x466;
  assign n7483 = ~n7481 & ~n7482;
  assign n7484 = ~n7480 & n7483;
  assign n7485 = x464 & n7484;
  assign n7486 = n7478 & n7479;
  assign n7487 = ~n7485 & ~n7486;
  assign n7488 = n7480 & ~n7483;
  assign n7492 = ~n7486 & ~n7488;
  assign n7493 = x464 & ~n7492;
  assign n7494 = ~x464 & ~n7484;
  assign n7495 = x463 & ~n7494;
  assign n7496 = ~n7493 & n7495;
  assign n9247 = n7487 & ~n7496;
  assign n7450 = x471 & x472;
  assign n7451 = x473 & x474;
  assign n7452 = n7450 & n7451;
  assign n7453 = ~x473 & ~x474;
  assign n7454 = x470 & ~n7453;
  assign n7455 = ~n7452 & ~n7454;
  assign n6692 = x472 ^ x471;
  assign n7456 = n7451 ^ x472;
  assign n7457 = n6692 & ~n7456;
  assign n7458 = n7457 ^ x471;
  assign n7459 = ~n7455 & n7458;
  assign n7470 = ~n7453 & n7458;
  assign n7471 = ~x470 & ~n7470;
  assign n7460 = ~x471 & ~x472;
  assign n7461 = ~n7451 & n7460;
  assign n7465 = x469 & ~n7461;
  assign n7466 = ~n7450 & n7453;
  assign n7472 = ~n7452 & ~n7466;
  assign n7473 = n7465 & n7472;
  assign n7474 = x469 & ~x470;
  assign n7475 = ~n7473 & ~n7474;
  assign n7476 = ~n7471 & ~n7475;
  assign n9246 = ~n7459 & ~n7476;
  assign n9248 = n9247 ^ n9246;
  assign n7489 = ~x464 & n7488;
  assign n7490 = n7487 & ~n7489;
  assign n7491 = ~x463 & ~n7490;
  assign n6688 = x464 ^ x463;
  assign n7497 = n7481 & n7482;
  assign n7498 = n6688 & n7497;
  assign n7499 = ~n7496 & ~n7498;
  assign n7500 = ~n7491 & n7499;
  assign n7462 = ~n7454 & n7461;
  assign n7463 = ~n7459 & ~n7462;
  assign n7464 = ~x469 & ~n7463;
  assign n7467 = ~x470 & n7466;
  assign n7468 = ~n7465 & n7467;
  assign n7469 = ~n7464 & ~n7468;
  assign n7477 = n7469 & ~n7476;
  assign n7501 = n7500 ^ n7477;
  assign n6687 = x468 ^ x467;
  assign n6689 = n6688 ^ n6687;
  assign n6686 = x466 ^ x465;
  assign n6690 = n6689 ^ n6686;
  assign n6693 = x474 ^ x473;
  assign n6694 = n6693 ^ n6692;
  assign n6691 = x470 ^ x469;
  assign n6695 = n6694 ^ n6691;
  assign n7502 = n6690 & n6695;
  assign n9243 = n7502 ^ n7500;
  assign n9244 = ~n7501 & n9243;
  assign n9245 = n9244 ^ n7502;
  assign n9249 = n9248 ^ n9245;
  assign n9257 = n9256 ^ n9249;
  assign n6685 = n6684 ^ n6679;
  assign n6696 = n6695 ^ n6690;
  assign n7503 = n6696 ^ n6684;
  assign n7504 = ~n6685 & n7503;
  assign n7505 = n7504 ^ n6696;
  assign n7507 = n7506 ^ n7505;
  assign n7508 = ~n7502 & ~n7507;
  assign n7509 = n7508 ^ n7506;
  assign n7563 = n7562 ^ n7509;
  assign n9258 = ~n7501 & ~n7563;
  assign n9259 = ~n7505 & ~n7562;
  assign n9260 = n7501 & n7502;
  assign n9261 = ~n9259 & ~n9260;
  assign n9262 = ~n9258 & n9261;
  assign n9263 = n7506 & n7562;
  assign n9264 = n9262 & ~n9263;
  assign n9594 = n9257 & n9264;
  assign n9595 = n9245 & n9256;
  assign n9596 = ~n9594 & ~n9595;
  assign n9597 = n9246 & n9247;
  assign n9598 = n9596 & n9597;
  assign n9599 = ~n9246 & ~n9247;
  assign n9600 = ~n9245 & ~n9599;
  assign n9601 = ~n9597 & ~n9600;
  assign n9602 = n9264 & n9601;
  assign n9603 = n9256 & n9602;
  assign n9604 = n9595 & n9599;
  assign n9605 = ~n9256 & n9600;
  assign n9606 = ~n9264 & n9605;
  assign n9607 = ~n9604 & ~n9606;
  assign n9608 = ~n9603 & n9607;
  assign n9609 = ~n9598 & n9608;
  assign n9591 = n9254 ^ n9252;
  assign n9592 = ~n9255 & ~n9591;
  assign n9593 = n9592 ^ n9252;
  assign n9610 = n9609 ^ n9593;
  assign n9265 = n9264 ^ n9257;
  assign n9290 = n9289 ^ n9265;
  assign n7564 = n7563 ^ n7501;
  assign n7449 = n7448 ^ n7400;
  assign n7565 = n7564 ^ n7449;
  assign n6697 = n6696 ^ n6685;
  assign n6720 = n6719 ^ n6708;
  assign n9239 = n6697 & n6720;
  assign n9240 = n9239 ^ n7449;
  assign n9241 = ~n7565 & ~n9240;
  assign n9242 = n9241 ^ n7564;
  assign n9588 = n9265 ^ n9242;
  assign n9589 = ~n9290 & n9588;
  assign n9590 = n9589 ^ n9289;
  assign n9611 = n9610 ^ n9590;
  assign n9629 = n9628 ^ n9611;
  assign n9351 = n9350 ^ n9302;
  assign n9292 = n7565 & n7780;
  assign n6721 = n6720 ^ n6697;
  assign n6768 = n6767 ^ n6744;
  assign n9293 = n6721 & n6768;
  assign n9294 = ~n9292 & n9293;
  assign n9295 = n9239 ^ n7565;
  assign n9297 = n9296 ^ n7780;
  assign n9298 = ~n9295 & ~n9297;
  assign n9299 = ~n9294 & ~n9298;
  assign n9352 = n9351 ^ n9299;
  assign n9291 = n9290 ^ n9242;
  assign n9585 = n9299 ^ n9291;
  assign n9586 = n9352 & n9585;
  assign n9587 = n9586 ^ n9351;
  assign n9630 = n9629 ^ n9587;
  assign n9678 = n9677 ^ n9652;
  assign n9866 = n9678 ^ n9587;
  assign n9867 = ~n9630 & ~n9866;
  assign n9868 = n9867 ^ n9678;
  assign n9877 = n9876 ^ n9868;
  assign n9884 = ~n9266 & ~n9628;
  assign n9885 = n9614 & ~n9623;
  assign n9886 = ~n9884 & ~n9885;
  assign n9887 = ~n9618 & ~n9886;
  assign n9888 = ~n9617 & ~n9628;
  assign n9889 = n9614 & n9620;
  assign n9890 = ~n9888 & ~n9889;
  assign n9891 = ~n9887 & n9890;
  assign n9881 = ~n9599 & n9610;
  assign n9882 = ~n9593 & n9596;
  assign n9883 = ~n9881 & ~n9882;
  assign n9892 = n9891 ^ n9883;
  assign n9878 = n9628 ^ n9610;
  assign n9879 = n9611 & n9878;
  assign n9880 = n9879 ^ n9628;
  assign n9893 = n9892 ^ n9880;
  assign n10027 = n9893 ^ n9876;
  assign n10028 = ~n9877 & ~n10027;
  assign n10029 = n10028 ^ n9893;
  assign n10030 = n9874 ^ n9871;
  assign n10031 = n9871 ^ n9669;
  assign n10032 = ~n10030 & n10031;
  assign n10033 = n10032 ^ n9669;
  assign n10034 = n9883 ^ n9880;
  assign n10035 = ~n9892 & ~n10034;
  assign n10036 = n10035 ^ n9891;
  assign n10103 = ~n10033 & n10036;
  assign n10104 = n10029 & n10103;
  assign n9894 = n9893 ^ n9877;
  assign n9583 = n9582 ^ n9533;
  assign n9353 = n9352 ^ n9291;
  assign n7348 = n7347 ^ n7113;
  assign n6769 = n6768 ^ n6721;
  assign n6867 = ~n6769 & ~n6866;
  assign n6868 = ~n6792 & ~n6815;
  assign n6869 = ~n6863 & n6868;
  assign n6870 = ~n6867 & ~n6869;
  assign n7350 = n6767 ^ n6697;
  assign n7352 = n7350 ^ n6744;
  assign n7353 = ~n6720 & n7352;
  assign n7351 = ~n6768 & ~n7350;
  assign n7354 = n7353 ^ n7351;
  assign n7566 = n7565 ^ n7354;
  assign n7781 = n7780 ^ n7566;
  assign n9227 = n6815 & n6863;
  assign n9228 = n7781 & ~n9227;
  assign n9229 = n6870 & ~n9228;
  assign n9230 = ~n7348 & ~n9229;
  assign n6872 = n6769 & n6863;
  assign n9231 = ~n6816 & n6872;
  assign n9232 = ~n7781 & n9231;
  assign n9233 = n6866 & n7348;
  assign n9234 = ~n9232 & n9233;
  assign n7974 = n6863 ^ n6816;
  assign n9235 = n6769 & n7974;
  assign n9236 = n7781 & ~n9235;
  assign n9237 = ~n9234 & ~n9236;
  assign n9238 = ~n9230 & n9237;
  assign n9354 = n9353 ^ n9238;
  assign n9423 = n9422 ^ n9360;
  assign n9481 = n9480 ^ n9423;
  assign n9486 = n9481 ^ n9238;
  assign n9487 = n9354 & n9486;
  assign n9488 = n9487 ^ n9353;
  assign n9584 = n9583 ^ n9488;
  assign n9679 = n9678 ^ n9630;
  assign n9863 = n9679 ^ n9488;
  assign n9864 = ~n9584 & n9863;
  assign n9865 = n9864 ^ n9679;
  assign n9895 = n9894 ^ n9865;
  assign n10024 = n9924 ^ n9894;
  assign n10025 = n9895 & n10024;
  assign n10026 = n10025 ^ n9924;
  assign n10037 = n10036 ^ n10033;
  assign n10097 = n10036 ^ n10029;
  assign n10098 = n10037 & n10097;
  assign n10099 = n10098 ^ n10029;
  assign n10109 = n10026 & n10099;
  assign n10110 = ~n10104 & ~n10109;
  assign n10111 = n10110 ^ n10052;
  assign n10112 = ~n10056 & n10111;
  assign n10090 = n9900 & n9903;
  assign n10091 = n10056 & ~n10090;
  assign n10092 = ~n10041 & ~n10050;
  assign n10093 = ~n10091 & ~n10092;
  assign n10094 = n10033 & ~n10036;
  assign n10095 = ~n10029 & n10094;
  assign n10096 = ~n10093 & n10095;
  assign n10100 = ~n10026 & ~n10099;
  assign n10101 = ~n10096 & ~n10100;
  assign n10119 = n10093 & ~n10104;
  assign n10120 = n10101 & ~n10119;
  assign n10121 = ~n10112 & ~n10120;
  assign n10134 = n10133 ^ n10121;
  assign n10072 = ~n9998 & ~n10020;
  assign n9994 = n9993 ^ n9990;
  assign n10073 = n9993 ^ n9987;
  assign n10074 = n9994 & ~n10073;
  assign n10075 = n10074 ^ n9987;
  assign n10076 = n10072 & ~n10075;
  assign n10079 = n10077 & n10078;
  assign n10080 = ~n10076 & ~n10079;
  assign n10082 = ~n9990 & n10081;
  assign n10083 = n10082 ^ n10075;
  assign n10084 = n9998 & n10083;
  assign n10085 = n10020 & n10084;
  assign n10086 = n10085 ^ n10082;
  assign n10087 = n10080 & ~n10086;
  assign n10088 = n10087 ^ n10071;
  assign n9995 = n9994 ^ n9987;
  assign n10022 = n10021 ^ n9995;
  assign n9925 = n9924 ^ n9895;
  assign n9680 = n9679 ^ n9584;
  assign n9225 = n9224 ^ n9220;
  assign n6873 = n6871 & n6872;
  assign n6874 = n6870 & ~n6873;
  assign n7349 = n7348 ^ n6874;
  assign n7782 = n7781 ^ n7349;
  assign n7973 = ~n7877 & ~n7972;
  assign n7975 = n7974 ^ n6769;
  assign n7976 = ~n7973 & n7975;
  assign n7977 = n7782 & ~n7976;
  assign n8998 = ~n7976 & ~n8997;
  assign n8999 = ~n7782 & ~n8998;
  assign n9000 = n8999 ^ n8997;
  assign n9001 = n8996 & ~n9000;
  assign n9002 = n9001 ^ n8997;
  assign n9003 = ~n7977 & ~n9002;
  assign n9226 = n9225 ^ n9003;
  assign n9482 = n9481 ^ n9354;
  assign n9483 = n9482 ^ n9003;
  assign n9484 = n9226 & n9483;
  assign n9485 = n9484 ^ n9225;
  assign n9681 = n9680 ^ n9485;
  assign n9859 = n9858 ^ n9769;
  assign n9860 = n9859 ^ n9485;
  assign n9861 = n9681 & ~n9860;
  assign n9862 = n9861 ^ n9680;
  assign n9926 = n9925 ^ n9862;
  assign n9981 = n9980 ^ n9929;
  assign n9982 = n9981 ^ n9925;
  assign n9983 = ~n9926 & n9982;
  assign n9984 = n9983 ^ n9981;
  assign n10023 = n10022 ^ n9984;
  assign n10038 = n10037 ^ n10029;
  assign n10039 = n10038 ^ n10026;
  assign n10057 = n10056 ^ n10039;
  assign n10058 = n10057 ^ n9984;
  assign n10059 = ~n10023 & n10058;
  assign n10060 = n10059 ^ n10022;
  assign n10089 = n10088 ^ n10060;
  assign n10102 = n10056 & n10101;
  assign n10105 = ~n10093 & ~n10104;
  assign n10106 = n10026 & ~n10095;
  assign n10107 = ~n10105 & n10106;
  assign n10108 = n10102 & ~n10107;
  assign n10113 = n10093 & n10104;
  assign n10114 = ~n10112 & ~n10113;
  assign n10115 = ~n10108 & n10114;
  assign n10116 = n10115 ^ n10060;
  assign n10117 = ~n10089 & ~n10116;
  assign n10118 = n10117 ^ n10088;
  assign n10135 = n10134 ^ n10118;
  assign n10137 = n10136 ^ n10135;
  assign n10180 = n6633 ^ n6629;
  assign n10139 = n6607 ^ n6606;
  assign n10138 = n10057 ^ n10023;
  assign n10140 = n10139 ^ n10138;
  assign n10171 = n6561 ^ n6560;
  assign n10141 = n6455 ^ n6454;
  assign n10142 = n9859 ^ n9681;
  assign n10143 = ~n10141 & n10142;
  assign n10145 = n6215 ^ n6214;
  assign n10144 = n9482 ^ n9226;
  assign n10146 = n10145 ^ n10144;
  assign n10151 = n4423 ^ n4421;
  assign n10152 = n6200 ^ n4423;
  assign n10153 = n10151 & ~n10152;
  assign n10154 = n10153 ^ n4421;
  assign n10155 = n10154 ^ n6202;
  assign n10156 = n10155 ^ n6199;
  assign n10147 = n8995 ^ n7976;
  assign n10148 = ~n8997 & ~n10147;
  assign n10149 = n10148 ^ n8994;
  assign n10150 = n10149 ^ n7782;
  assign n10157 = n10156 ^ n10150;
  assign n10158 = n10151 ^ n6200;
  assign n10159 = n7972 ^ n7877;
  assign n10160 = n10159 ^ n7975;
  assign n10161 = n10158 & n10160;
  assign n10162 = n10161 ^ n10150;
  assign n10163 = ~n10157 & n10162;
  assign n10164 = n10163 ^ n10156;
  assign n10165 = n10164 ^ n10144;
  assign n10166 = n10146 & n10165;
  assign n10167 = n10166 ^ n10145;
  assign n10168 = ~n10143 & n10167;
  assign n10169 = n10141 & ~n10142;
  assign n10170 = ~n10168 & ~n10169;
  assign n10172 = n10171 ^ n10170;
  assign n10173 = n9981 ^ n9926;
  assign n10174 = n10173 ^ n10170;
  assign n10175 = ~n10172 & ~n10174;
  assign n10176 = n10175 ^ n10171;
  assign n10177 = n10176 ^ n10138;
  assign n10178 = n10140 & n10177;
  assign n10179 = n10178 ^ n10139;
  assign n10181 = n10180 ^ n10179;
  assign n10182 = n10115 ^ n10089;
  assign n10183 = n10182 ^ n10180;
  assign n10184 = ~n10181 & n10183;
  assign n10185 = n10184 ^ n10179;
  assign n10186 = n10185 ^ n10135;
  assign n10187 = n10137 & ~n10186;
  assign n10188 = n10187 ^ n10136;
  assign n10189 = n6674 & ~n10188;
  assign n10190 = n10133 ^ n10118;
  assign n10191 = ~n10134 & n10190;
  assign n10192 = n10191 ^ n10118;
  assign n10193 = n10189 & ~n10192;
  assign n10194 = n10137 & n10185;
  assign n10195 = ~n10179 & n10180;
  assign n10196 = ~n10182 & n10195;
  assign n10197 = ~n10170 & n10171;
  assign n10198 = ~n10173 & n10197;
  assign n10199 = n10176 & ~n10198;
  assign n10200 = n10140 & ~n10199;
  assign n10201 = n10168 & ~n10169;
  assign n10202 = n10142 ^ n10141;
  assign n10203 = n10144 & n10145;
  assign n10204 = ~n10164 & n10203;
  assign n10205 = n10160 ^ n10158;
  assign n10206 = n10160 ^ n10157;
  assign n10207 = ~n10205 & n10206;
  assign n10208 = ~x1000 & n10207;
  assign n10209 = ~n10204 & ~n10208;
  assign n10210 = n10167 & ~n10209;
  assign n10211 = n10202 & ~n10210;
  assign n10212 = ~n10144 & ~n10145;
  assign n10213 = n10164 & ~n10208;
  assign n10214 = n10212 & n10213;
  assign n10215 = ~n10211 & ~n10214;
  assign n10216 = ~n10201 & n10215;
  assign n10217 = ~n10200 & ~n10216;
  assign n10218 = n10170 & ~n10171;
  assign n10219 = n10173 & n10218;
  assign n10220 = ~n10140 & ~n10219;
  assign n10221 = n10217 & ~n10220;
  assign n10222 = ~n10196 & n10221;
  assign n10223 = ~n10194 & n10222;
  assign n10224 = n10179 & ~n10180;
  assign n10225 = n10182 & n10224;
  assign n10226 = ~n10137 & ~n10225;
  assign n10227 = n10223 & ~n10226;
  assign n10228 = ~n10193 & n10227;
  assign n10229 = ~n10189 & n10192;
  assign n10230 = n10188 ^ n6673;
  assign n10231 = n6673 ^ n4475;
  assign n10232 = ~n10230 & n10231;
  assign n10233 = n10232 ^ n10188;
  assign n10234 = ~n10229 & ~n10233;
  assign n10235 = ~n10228 & n10234;
  assign y0 = ~n10235;
endmodule
