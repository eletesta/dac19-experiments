module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700, x701, x702, x703, x704, x705, x706, x707, x708, x709, x710, x711, x712, x713, x714, x715, x716, x717, x718, x719, x720, x721, x722, x723, x724, x725, x726, x727, x728, x729, x730, x731, x732, x733, x734, x735, x736, x737, x738, x739, x740, x741, x742, x743, x744, x745, x746, x747, x748, x749, x750, x751, x752, x753, x754, x755, x756, x757, x758, x759, x760, x761, x762, x763, x764, x765, x766, x767, x768, x769, x770, x771, x772, x773, x774, x775, x776, x777, x778, x779, x780, x781, x782, x783, x784, x785, x786, x787, x788, x789, x790, x791, x792, x793, x794, x795, x796, x797, x798, x799, x800, x801, x802, x803, x804, x805, x806, x807, x808, x809, x810, x811, x812, x813, x814, x815, x816, x817, x818, x819, x820, x821, x822, x823, x824, x825, x826, x827, x828, x829, x830, x831, x832, x833, x834, x835, x836, x837, x838, x839, x840, x841, x842, x843, x844, x845, x846, x847, x848, x849, x850, x851, x852, x853, x854, x855, x856, x857, x858, x859, x860, x861, x862, x863, x864, x865, x866, x867, x868, x869, x870, x871, x872, x873, x874, x875, x876, x877, x878, x879, x880, x881, x882, x883, x884, x885, x886, x887, x888, x889, x890, x891, x892, x893, x894, x895, x896, x897, x898, x899, x900, x901, x902, x903, x904, x905, x906, x907, x908, x909, x910, x911, x912, x913, x914, x915, x916, x917, x918, x919, x920, x921, x922, x923, x924, x925, x926, x927, x928, x929, x930, x931, x932, x933, x934, x935, x936, x937, x938, x939, x940, x941, x942, x943, x944, x945, x946, x947, x948, x949, x950, x951, x952, x953, x954, x955, x956, x957, x958, x959, x960, x961, x962, x963, x964, x965, x966, x967, x968, x969, x970, x971, x972, x973, x974, x975, x976, x977, x978, x979, x980, x981, x982, x983, x984, x985, x986, x987, x988, x989, x990, x991, x992, x993, x994, x995, x996, x997, x998, x999, x1000, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700, x701, x702, x703, x704, x705, x706, x707, x708, x709, x710, x711, x712, x713, x714, x715, x716, x717, x718, x719, x720, x721, x722, x723, x724, x725, x726, x727, x728, x729, x730, x731, x732, x733, x734, x735, x736, x737, x738, x739, x740, x741, x742, x743, x744, x745, x746, x747, x748, x749, x750, x751, x752, x753, x754, x755, x756, x757, x758, x759, x760, x761, x762, x763, x764, x765, x766, x767, x768, x769, x770, x771, x772, x773, x774, x775, x776, x777, x778, x779, x780, x781, x782, x783, x784, x785, x786, x787, x788, x789, x790, x791, x792, x793, x794, x795, x796, x797, x798, x799, x800, x801, x802, x803, x804, x805, x806, x807, x808, x809, x810, x811, x812, x813, x814, x815, x816, x817, x818, x819, x820, x821, x822, x823, x824, x825, x826, x827, x828, x829, x830, x831, x832, x833, x834, x835, x836, x837, x838, x839, x840, x841, x842, x843, x844, x845, x846, x847, x848, x849, x850, x851, x852, x853, x854, x855, x856, x857, x858, x859, x860, x861, x862, x863, x864, x865, x866, x867, x868, x869, x870, x871, x872, x873, x874, x875, x876, x877, x878, x879, x880, x881, x882, x883, x884, x885, x886, x887, x888, x889, x890, x891, x892, x893, x894, x895, x896, x897, x898, x899, x900, x901, x902, x903, x904, x905, x906, x907, x908, x909, x910, x911, x912, x913, x914, x915, x916, x917, x918, x919, x920, x921, x922, x923, x924, x925, x926, x927, x928, x929, x930, x931, x932, x933, x934, x935, x936, x937, x938, x939, x940, x941, x942, x943, x944, x945, x946, x947, x948, x949, x950, x951, x952, x953, x954, x955, x956, x957, x958, x959, x960, x961, x962, x963, x964, x965, x966, x967, x968, x969, x970, x971, x972, x973, x974, x975, x976, x977, x978, x979, x980, x981, x982, x983, x984, x985, x986, x987, x988, x989, x990, x991, x992, x993, x994, x995, x996, x997, x998, x999, x1000;
  output y0;
  wire n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964;
  assign n4619 = x189 & x190;
  assign n4618 = x191 & x192;
  assign n4620 = n4619 ^ n4618;
  assign n4621 = ~x189 & ~x190;
  assign n4622 = ~x191 & ~x192;
  assign n4623 = ~n4621 & ~n4622;
  assign n4624 = n4623 ^ n4618;
  assign n4625 = n4624 ^ n4618;
  assign n4626 = n4618 ^ x188;
  assign n4627 = n4626 ^ n4618;
  assign n4628 = n4625 & n4627;
  assign n4629 = n4628 ^ n4618;
  assign n4630 = n4620 & ~n4629;
  assign n4631 = n4630 ^ n4619;
  assign n4633 = ~n4618 & ~n4619;
  assign n4646 = n4623 & ~n4633;
  assign n4645 = x192 & n4619;
  assign n4647 = n4646 ^ n4645;
  assign n4648 = n4647 ^ n4646;
  assign n4649 = ~n4623 & n4633;
  assign n4650 = n4649 ^ n4646;
  assign n4651 = n4650 ^ n4646;
  assign n4652 = ~n4648 & ~n4651;
  assign n4653 = n4652 ^ n4646;
  assign n4654 = x188 & n4653;
  assign n4655 = n4654 ^ n4646;
  assign n6582 = x187 & n4655;
  assign n6583 = ~n4631 & ~n6582;
  assign n4663 = x197 & x198;
  assign n4664 = x195 & x196;
  assign n4668 = n4663 & n4664;
  assign n4672 = x193 & x194;
  assign n4674 = ~n4668 & n4672;
  assign n4665 = ~n4663 & ~n4664;
  assign n4675 = n4674 ^ n4665;
  assign n3043 = x194 ^ x193;
  assign n4676 = n4674 ^ n3043;
  assign n4660 = ~x197 & ~x198;
  assign n4661 = ~x195 & ~x196;
  assign n4662 = ~n4660 & ~n4661;
  assign n4677 = n4665 ^ n4662;
  assign n4678 = n4677 ^ n4674;
  assign n4679 = ~n4674 & ~n4678;
  assign n4680 = n4679 ^ n4674;
  assign n4681 = n4676 & ~n4680;
  assign n4682 = n4681 ^ n4679;
  assign n4683 = n4682 ^ n4674;
  assign n4684 = n4683 ^ n4677;
  assign n4685 = ~n4675 & ~n4684;
  assign n4686 = n4685 ^ n4674;
  assign n6581 = ~n4668 & ~n4686;
  assign n6584 = n6583 ^ n6581;
  assign n4666 = ~n4662 & n4665;
  assign n4667 = ~n3043 & n4666;
  assign n4669 = n4660 & n4661;
  assign n4670 = ~n4668 & ~n4669;
  assign n4671 = ~n4667 & n4670;
  assign n4673 = ~n4671 & ~n4672;
  assign n4687 = ~n4673 & ~n4686;
  assign n3038 = x190 ^ x189;
  assign n4609 = x187 & x188;
  assign n4610 = n4609 ^ x190;
  assign n4611 = n4610 ^ n4609;
  assign n4612 = ~x188 & ~x192;
  assign n4613 = n4612 ^ n4609;
  assign n4614 = ~n4611 & n4613;
  assign n4615 = n4614 ^ n4609;
  assign n4616 = ~n3038 & n4615;
  assign n4617 = ~x191 & n4616;
  assign n4632 = n4622 ^ n4621;
  assign n4634 = n4633 ^ n4622;
  assign n4635 = n4634 ^ n4622;
  assign n4636 = n4622 ^ x188;
  assign n4637 = n4636 ^ n4622;
  assign n4638 = n4635 & ~n4637;
  assign n4639 = n4638 ^ n4622;
  assign n4640 = n4632 & ~n4639;
  assign n4641 = n4640 ^ n4621;
  assign n4642 = ~n4631 & ~n4641;
  assign n4643 = n4642 ^ x187;
  assign n4644 = n4643 ^ n4642;
  assign n4656 = n4655 ^ n4642;
  assign n4657 = n4644 & ~n4656;
  assign n4658 = n4657 ^ n4642;
  assign n4659 = ~n4617 & n4658;
  assign n4688 = n4687 ^ n4659;
  assign n3037 = x192 ^ x191;
  assign n3039 = n3038 ^ n3037;
  assign n3036 = x188 ^ x187;
  assign n3040 = n3039 ^ n3036;
  assign n3042 = x198 ^ x197;
  assign n3044 = n3043 ^ n3042;
  assign n3041 = x196 ^ x195;
  assign n3045 = n3044 ^ n3041;
  assign n4608 = n3040 & n3045;
  assign n6578 = n4687 ^ n4608;
  assign n6579 = n4688 & ~n6578;
  assign n6580 = n6579 ^ n4659;
  assign n6585 = n6584 ^ n6580;
  assign n4536 = x179 & x180;
  assign n4537 = x177 & x178;
  assign n4538 = ~n4536 & ~n4537;
  assign n4539 = ~x179 & ~x180;
  assign n4540 = ~x177 & ~x178;
  assign n4541 = ~n4539 & ~n4540;
  assign n4542 = ~n4538 & n4541;
  assign n4543 = x176 & n4542;
  assign n4544 = n4536 & n4537;
  assign n4545 = ~n4543 & ~n4544;
  assign n4552 = n4542 ^ x176;
  assign n4553 = n4552 ^ n4542;
  assign n4546 = n4538 & ~n4541;
  assign n4554 = ~n4544 & ~n4546;
  assign n4555 = n4554 ^ n4542;
  assign n4556 = n4553 & n4555;
  assign n4557 = n4556 ^ n4542;
  assign n4558 = x175 & n4557;
  assign n6575 = n4545 & ~n4558;
  assign n4562 = x185 & x186;
  assign n4561 = x183 & x184;
  assign n4563 = n4562 ^ n4561;
  assign n4564 = ~x185 & ~x186;
  assign n4565 = ~x183 & ~x184;
  assign n4566 = ~n4564 & ~n4565;
  assign n4567 = n4566 ^ n4561;
  assign n4568 = n4567 ^ n4561;
  assign n4569 = n4561 ^ x182;
  assign n4570 = n4569 ^ n4561;
  assign n4571 = n4568 & n4570;
  assign n4572 = n4571 ^ n4561;
  assign n4573 = n4563 & ~n4572;
  assign n4574 = n4573 ^ n4562;
  assign n3054 = x182 ^ x181;
  assign n4576 = ~n4561 & ~n4562;
  assign n4587 = n4566 & ~n4576;
  assign n4588 = n3054 & n4587;
  assign n4589 = ~n4566 & n4576;
  assign n4590 = x181 & x182;
  assign n4591 = n4561 & n4590;
  assign n4592 = x186 & n4591;
  assign n4593 = n4592 ^ n4590;
  assign n4594 = ~n4589 & n4593;
  assign n4595 = ~n4588 & ~n4594;
  assign n6574 = ~n4574 & n4595;
  assign n6576 = n6575 ^ n6574;
  assign n4575 = n4565 ^ n4564;
  assign n4577 = n4576 ^ n4565;
  assign n4578 = n4577 ^ n4565;
  assign n4579 = n4565 ^ x182;
  assign n4580 = n4579 ^ n4565;
  assign n4581 = n4578 & ~n4580;
  assign n4582 = n4581 ^ n4565;
  assign n4583 = n4575 & ~n4582;
  assign n4584 = n4583 ^ n4564;
  assign n4585 = ~n4574 & ~n4584;
  assign n4586 = ~x181 & ~n4585;
  assign n3053 = x184 ^ x183;
  assign n4596 = n4590 ^ x184;
  assign n4597 = n4596 ^ n4590;
  assign n4598 = ~x182 & ~x186;
  assign n4599 = n4598 ^ n4590;
  assign n4600 = ~n4597 & n4599;
  assign n4601 = n4600 ^ n4590;
  assign n4602 = ~n3053 & n4601;
  assign n4603 = ~x185 & n4602;
  assign n4604 = n4595 & ~n4603;
  assign n4605 = ~n4586 & n4604;
  assign n4547 = ~x176 & n4546;
  assign n4548 = n4545 & ~n4547;
  assign n4549 = ~x175 & ~n4548;
  assign n3049 = x176 ^ x175;
  assign n4550 = n4539 & n4540;
  assign n4551 = n3049 & n4550;
  assign n4559 = ~n4551 & ~n4558;
  assign n4560 = ~n4549 & n4559;
  assign n4606 = n4605 ^ n4560;
  assign n3048 = x178 ^ x177;
  assign n3050 = n3049 ^ n3048;
  assign n3047 = x180 ^ x179;
  assign n3051 = n3050 ^ n3047;
  assign n3055 = n3054 ^ n3053;
  assign n3052 = x186 ^ x185;
  assign n3056 = n3055 ^ n3052;
  assign n4535 = n3051 & n3056;
  assign n6571 = n4560 ^ n4535;
  assign n6572 = n4606 & ~n6571;
  assign n6573 = n6572 ^ n4605;
  assign n6577 = n6576 ^ n6573;
  assign n6586 = n6585 ^ n6577;
  assign n4689 = n4688 ^ n4608;
  assign n4607 = n4606 ^ n4535;
  assign n4690 = n4689 ^ n4607;
  assign n3046 = n3045 ^ n3040;
  assign n3057 = n3056 ^ n3051;
  assign n6540 = n3046 & n3057;
  assign n6568 = n6540 ^ n4607;
  assign n6569 = n4690 & ~n6568;
  assign n6570 = n6569 ^ n4689;
  assign n6587 = n6586 ^ n6570;
  assign n6947 = ~n6570 & n6574;
  assign n6948 = ~n6587 & ~n6947;
  assign n6949 = n6575 ^ n6573;
  assign n6950 = n6585 ^ n6573;
  assign n6951 = n6949 & n6950;
  assign n6952 = n6951 ^ n6585;
  assign n6953 = n6948 & n6952;
  assign n6954 = n6574 ^ n6570;
  assign n6955 = n6587 ^ n6574;
  assign n6956 = ~n6954 & n6955;
  assign n6957 = n6956 ^ n6574;
  assign n6958 = ~n6952 & n6957;
  assign n6959 = ~n6953 & ~n6958;
  assign n6944 = n6583 ^ n6580;
  assign n6945 = ~n6584 & ~n6944;
  assign n6946 = n6945 ^ n6580;
  assign n6960 = n6959 ^ n6946;
  assign n3061 = x206 ^ x205;
  assign n4778 = ~x209 & ~x210;
  assign n4783 = n3061 & ~n4778;
  assign n3060 = x208 ^ x207;
  assign n4771 = x209 & x210;
  assign n4785 = n4771 ^ x208;
  assign n4786 = n3060 & ~n4785;
  assign n4787 = n4786 ^ x207;
  assign n4788 = n4783 & n4787;
  assign n4773 = x207 & x208;
  assign n4772 = ~x207 & ~x208;
  assign n4774 = n4773 ^ n4772;
  assign n4775 = ~n4771 & n4774;
  assign n4776 = n4775 ^ n4773;
  assign n4779 = ~n4773 & n4778;
  assign n4789 = x205 & x206;
  assign n4790 = ~n4779 & n4789;
  assign n4791 = ~n4776 & n4790;
  assign n4792 = ~n4788 & ~n4791;
  assign n6545 = n4771 & n4773;
  assign n6546 = n4792 & ~n6545;
  assign n4794 = ~x203 & ~x204;
  assign n4795 = x200 & ~n4794;
  assign n4796 = x203 & x204;
  assign n4797 = ~x201 & ~x202;
  assign n4798 = ~n4796 & n4797;
  assign n4799 = ~n4795 & n4798;
  assign n4800 = x201 & x202;
  assign n4801 = n4800 ^ n4796;
  assign n4802 = n4800 ^ n4795;
  assign n4803 = n4801 & n4802;
  assign n4804 = n4803 ^ n4800;
  assign n4805 = ~n4797 & n4804;
  assign n4806 = ~n4799 & ~n4805;
  assign n4807 = ~x199 & ~n4806;
  assign n4808 = ~n4796 & ~n4800;
  assign n4809 = ~n4797 & ~n4808;
  assign n4810 = x199 & ~n4794;
  assign n4811 = n4809 & n4810;
  assign n4812 = x199 & x200;
  assign n4813 = ~n4811 & ~n4812;
  assign n4814 = ~n4794 & ~n4800;
  assign n4815 = ~n4798 & n4814;
  assign n4816 = ~x204 & n4800;
  assign n4817 = x200 & ~n4816;
  assign n4818 = ~n4815 & n4817;
  assign n4819 = ~n4813 & ~n4818;
  assign n4820 = ~n4807 & ~n4819;
  assign n4821 = ~x200 & ~x204;
  assign n4822 = n4821 ^ n4812;
  assign n4823 = n4822 ^ n4812;
  assign n4824 = x199 & ~n4797;
  assign n4825 = n4824 ^ n4812;
  assign n4826 = n4825 ^ n4812;
  assign n4827 = n4823 & ~n4826;
  assign n4828 = n4827 ^ n4812;
  assign n4829 = ~n4800 & n4828;
  assign n4830 = n4829 ^ n4812;
  assign n4831 = ~x203 & n4830;
  assign n4832 = n4820 & ~n4831;
  assign n4777 = ~x205 & n4776;
  assign n3062 = n3061 ^ n3060;
  assign n4780 = ~x206 & n4779;
  assign n4781 = n3062 & n4780;
  assign n4782 = ~n4777 & ~n4781;
  assign n4784 = ~n4782 & ~n4783;
  assign n4793 = ~n4784 & n4792;
  assign n4833 = n4832 ^ n4793;
  assign n3072 = x222 ^ x221;
  assign n3071 = x218 ^ x217;
  assign n3073 = n3072 ^ n3071;
  assign n3070 = x220 ^ x219;
  assign n3074 = n3073 ^ n3070;
  assign n3077 = x216 ^ x215;
  assign n3076 = x212 ^ x211;
  assign n3078 = n3077 ^ n3076;
  assign n3075 = x214 ^ x213;
  assign n3079 = n3078 ^ n3075;
  assign n4763 = n3074 & n3079;
  assign n3059 = x210 ^ x209;
  assign n3063 = n3062 ^ n3059;
  assign n3066 = x204 ^ x203;
  assign n3065 = x202 ^ x201;
  assign n3067 = n3066 ^ n3065;
  assign n3064 = x200 ^ x199;
  assign n3068 = n3067 ^ n3064;
  assign n4767 = n3063 & n3068;
  assign n3069 = n3068 ^ n3063;
  assign n3080 = n3079 ^ n3074;
  assign n4764 = n3080 ^ n3068;
  assign n4765 = ~n3069 & n4764;
  assign n4766 = n4765 ^ n3080;
  assign n4768 = n4767 ^ n4766;
  assign n4769 = ~n4763 & ~n4768;
  assign n4770 = n4769 ^ n4767;
  assign n4834 = n4833 ^ n4770;
  assign n4737 = x213 & x214;
  assign n4738 = x215 & x216;
  assign n4739 = ~n4737 & ~n4738;
  assign n4740 = ~x213 & ~x214;
  assign n4741 = ~x215 & ~x216;
  assign n4742 = ~n4740 & ~n4741;
  assign n4743 = ~n4739 & n4742;
  assign n4744 = x212 & n4743;
  assign n4745 = n4737 & n4738;
  assign n4746 = ~n4744 & ~n4745;
  assign n4747 = n4739 & ~n4742;
  assign n4748 = ~x212 & n4747;
  assign n4749 = n4746 & ~n4748;
  assign n4750 = ~x211 & ~n4749;
  assign n4751 = n4740 & n4741;
  assign n4752 = n3076 & n4751;
  assign n4753 = n4743 ^ x212;
  assign n4754 = n4753 ^ n4743;
  assign n4755 = ~n4745 & ~n4747;
  assign n4756 = n4755 ^ n4743;
  assign n4757 = n4754 & n4756;
  assign n4758 = n4757 ^ n4743;
  assign n4759 = x211 & n4758;
  assign n4760 = ~n4752 & ~n4759;
  assign n4761 = ~n4750 & n4760;
  assign n4693 = x221 & x222;
  assign n4692 = x219 & x220;
  assign n4694 = n4693 ^ n4692;
  assign n4695 = ~x221 & ~x222;
  assign n4696 = ~x219 & ~x220;
  assign n4697 = ~n4695 & ~n4696;
  assign n4698 = n4697 ^ n4692;
  assign n4699 = n4698 ^ n4692;
  assign n4700 = n4692 ^ x218;
  assign n4701 = n4700 ^ n4692;
  assign n4702 = n4699 & n4701;
  assign n4703 = n4702 ^ n4692;
  assign n4704 = n4694 & ~n4703;
  assign n4705 = n4704 ^ n4693;
  assign n4706 = n4696 ^ n4695;
  assign n4707 = ~n4692 & ~n4693;
  assign n4708 = n4707 ^ n4696;
  assign n4709 = n4708 ^ n4696;
  assign n4710 = n4696 ^ x218;
  assign n4711 = n4710 ^ n4696;
  assign n4712 = n4709 & ~n4711;
  assign n4713 = n4712 ^ n4696;
  assign n4714 = n4706 & ~n4713;
  assign n4715 = n4714 ^ n4695;
  assign n4716 = ~n4705 & ~n4715;
  assign n4717 = ~x217 & ~n4716;
  assign n4718 = n4697 & ~n4707;
  assign n4719 = n3071 & n4718;
  assign n4720 = ~n4697 & n4707;
  assign n4721 = x217 & x218;
  assign n4722 = n4692 & n4721;
  assign n4723 = x222 & n4722;
  assign n4724 = n4723 ^ n4721;
  assign n4725 = ~n4720 & n4724;
  assign n4726 = ~n4719 & ~n4725;
  assign n4727 = n4721 ^ x220;
  assign n4728 = n4727 ^ n4721;
  assign n4729 = ~x218 & ~x222;
  assign n4730 = n4729 ^ n4721;
  assign n4731 = ~n4728 & n4730;
  assign n4732 = n4731 ^ n4721;
  assign n4733 = ~n3070 & n4732;
  assign n4734 = ~x221 & n4733;
  assign n4735 = n4726 & ~n4734;
  assign n4736 = ~n4717 & n4735;
  assign n4762 = n4761 ^ n4736;
  assign n4835 = n4834 ^ n4762;
  assign n6560 = n4762 & ~n4763;
  assign n6561 = ~n4835 & ~n6560;
  assign n6562 = ~n4768 & ~n4833;
  assign n6563 = n6562 ^ n4767;
  assign n6564 = ~n6561 & ~n6563;
  assign n6556 = n4746 & ~n4759;
  assign n6555 = ~n4705 & n4726;
  assign n6557 = n6556 ^ n6555;
  assign n6552 = n4763 ^ n4761;
  assign n6553 = ~n4762 & n6552;
  assign n6554 = n6553 ^ n4763;
  assign n6558 = n6557 ^ n6554;
  assign n6548 = n4767 & n4833;
  assign n6549 = n4793 & n4832;
  assign n6550 = ~n6548 & ~n6549;
  assign n6547 = ~n4805 & ~n4819;
  assign n6551 = n6550 ^ n6547;
  assign n6559 = n6558 ^ n6551;
  assign n6565 = n6564 ^ n6559;
  assign n6931 = n6546 & n6565;
  assign n6932 = n6564 ^ n6550;
  assign n6933 = ~n6551 & ~n6932;
  assign n6934 = n6933 ^ n6564;
  assign n6935 = n6931 & ~n6934;
  assign n6936 = n6547 & n6550;
  assign n6937 = ~n6558 & n6936;
  assign n6938 = ~n6564 & n6937;
  assign n6939 = ~n6935 & ~n6938;
  assign n6566 = n6565 ^ n6546;
  assign n6940 = n6558 & n6934;
  assign n6941 = n6566 & n6940;
  assign n6942 = n6939 & ~n6941;
  assign n6928 = n6556 ^ n6554;
  assign n6929 = ~n6557 & ~n6928;
  assign n6930 = n6929 ^ n6554;
  assign n6943 = n6942 ^ n6930;
  assign n6961 = n6960 ^ n6943;
  assign n3058 = n3057 ^ n3046;
  assign n3081 = n3080 ^ n3069;
  assign n4532 = n3081 ^ n3046;
  assign n4533 = n3058 & ~n4532;
  assign n4534 = n4533 ^ n3057;
  assign n4691 = n4690 ^ n4534;
  assign n6539 = n4691 & n4835;
  assign n6541 = n4690 & n6540;
  assign n6542 = ~n4534 & ~n4690;
  assign n6543 = ~n6541 & ~n6542;
  assign n6544 = ~n6539 & n6543;
  assign n6567 = n6566 ^ n6544;
  assign n6925 = n6587 ^ n6566;
  assign n6926 = n6567 & ~n6925;
  assign n6927 = n6926 ^ n6587;
  assign n7341 = n6943 ^ n6927;
  assign n7342 = n6961 & ~n7341;
  assign n7343 = n7342 ^ n6960;
  assign n7344 = ~n6946 & ~n6953;
  assign n7345 = ~n6958 & ~n7344;
  assign n7346 = ~n6930 & ~n6941;
  assign n7347 = n6939 & ~n7346;
  assign n7568 = ~n7345 & ~n7347;
  assign n7591 = ~n7343 & n7568;
  assign n4972 = x243 & x244;
  assign n4973 = x245 & x246;
  assign n4985 = n4972 & n4973;
  assign n4992 = x241 & x242;
  assign n4993 = ~n4985 & n4992;
  assign n4975 = ~x243 & ~x244;
  assign n4976 = ~x245 & ~x246;
  assign n4977 = ~n4975 & ~n4976;
  assign n4994 = n4993 ^ n4977;
  assign n3025 = x242 ^ x241;
  assign n4995 = n4993 ^ n3025;
  assign n4974 = ~n4972 & ~n4973;
  assign n4996 = n4977 ^ n4974;
  assign n4997 = n4996 ^ n4993;
  assign n4998 = ~n4993 & ~n4997;
  assign n4999 = n4998 ^ n4993;
  assign n5000 = n4995 & ~n4999;
  assign n5001 = n5000 ^ n4998;
  assign n5002 = n5001 ^ n4993;
  assign n5003 = n5002 ^ n4996;
  assign n5004 = n4994 & ~n5003;
  assign n5005 = n5004 ^ n4993;
  assign n6520 = ~n4985 & ~n5005;
  assign n5007 = x239 & x240;
  assign n5008 = x237 & x238;
  assign n5015 = n5007 & n5008;
  assign n5019 = x235 & x236;
  assign n5021 = ~n5015 & n5019;
  assign n5010 = ~x239 & ~x240;
  assign n5011 = ~x237 & ~x238;
  assign n5012 = ~n5010 & ~n5011;
  assign n5022 = n5021 ^ n5012;
  assign n3030 = x236 ^ x235;
  assign n5023 = n5021 ^ n3030;
  assign n5009 = ~n5007 & ~n5008;
  assign n5024 = n5012 ^ n5009;
  assign n5025 = n5024 ^ n5021;
  assign n5026 = ~n5021 & ~n5025;
  assign n5027 = n5026 ^ n5021;
  assign n5028 = n5023 & ~n5027;
  assign n5029 = n5028 ^ n5026;
  assign n5030 = n5029 ^ n5021;
  assign n5031 = n5030 ^ n5024;
  assign n5032 = n5022 & ~n5031;
  assign n5033 = n5032 ^ n5021;
  assign n6521 = ~n5015 & ~n5033;
  assign n6915 = ~n6520 & ~n6521;
  assign n5063 = x225 & x226;
  assign n5064 = x227 & x228;
  assign n5065 = ~n5063 & ~n5064;
  assign n5066 = ~x225 & ~x226;
  assign n5067 = ~x227 & ~x228;
  assign n5068 = ~n5066 & ~n5067;
  assign n5069 = ~n5065 & n5068;
  assign n5070 = x224 & n5069;
  assign n5071 = n5063 & n5064;
  assign n5072 = ~n5070 & ~n5071;
  assign n5073 = n5065 & ~n5068;
  assign n5074 = ~x224 & n5073;
  assign n5075 = n5072 & ~n5074;
  assign n5076 = ~x223 & ~n5075;
  assign n3019 = x224 ^ x223;
  assign n5077 = n5066 & n5067;
  assign n5078 = n3019 & n5077;
  assign n5079 = n5069 ^ x224;
  assign n5080 = n5079 ^ n5069;
  assign n5081 = ~n5071 & ~n5073;
  assign n5082 = n5081 ^ n5069;
  assign n5083 = n5080 & n5082;
  assign n5084 = n5083 ^ n5069;
  assign n5085 = x223 & n5084;
  assign n5086 = ~n5078 & ~n5085;
  assign n5087 = ~n5076 & n5086;
  assign n5038 = x231 & x232;
  assign n5039 = x233 & x234;
  assign n5040 = ~n5038 & ~n5039;
  assign n5041 = ~x231 & ~x232;
  assign n5042 = ~x233 & ~x234;
  assign n5043 = ~n5041 & ~n5042;
  assign n5044 = ~n5040 & n5043;
  assign n5045 = x230 & n5044;
  assign n5046 = n5038 & n5039;
  assign n5047 = ~n5045 & ~n5046;
  assign n5048 = n5040 & ~n5043;
  assign n5049 = ~x230 & n5048;
  assign n5050 = n5047 & ~n5049;
  assign n5051 = ~x229 & ~n5050;
  assign n3014 = x230 ^ x229;
  assign n5052 = n5041 & n5042;
  assign n5053 = n3014 & n5052;
  assign n5054 = n5044 ^ x230;
  assign n5055 = n5054 ^ n5044;
  assign n5056 = ~n5046 & ~n5048;
  assign n5057 = n5056 ^ n5044;
  assign n5058 = n5055 & n5057;
  assign n5059 = n5058 ^ n5044;
  assign n5060 = x229 & n5059;
  assign n5061 = ~n5053 & ~n5060;
  assign n5062 = ~n5051 & n5061;
  assign n5088 = n5087 ^ n5062;
  assign n3013 = x234 ^ x233;
  assign n3015 = n3014 ^ n3013;
  assign n3012 = x232 ^ x231;
  assign n3016 = n3015 ^ n3012;
  assign n3018 = x228 ^ x227;
  assign n3020 = n3019 ^ n3018;
  assign n3017 = x226 ^ x225;
  assign n3021 = n3020 ^ n3017;
  assign n5037 = n3016 & n3021;
  assign n5089 = n5088 ^ n5037;
  assign n5013 = n5009 & ~n5012;
  assign n5014 = ~n3030 & n5013;
  assign n5016 = n5010 & n5011;
  assign n5017 = ~n5015 & ~n5016;
  assign n5018 = ~n5014 & n5017;
  assign n5020 = ~n5018 & ~n5019;
  assign n5034 = ~n5020 & ~n5033;
  assign n4978 = n4974 & ~n4977;
  assign n4979 = ~x241 & ~x242;
  assign n4980 = n4978 & n4979;
  assign n4981 = n4975 & n4976;
  assign n4982 = n4981 ^ x241;
  assign n4983 = n4981 ^ x242;
  assign n4984 = n4983 ^ x242;
  assign n4986 = n4985 ^ x242;
  assign n4987 = ~n4984 & n4986;
  assign n4988 = n4987 ^ x242;
  assign n4989 = ~n4982 & ~n4988;
  assign n4990 = n4989 ^ x241;
  assign n4991 = ~n4980 & n4990;
  assign n5006 = n4991 & ~n5005;
  assign n5035 = n5034 ^ n5006;
  assign n3024 = x246 ^ x245;
  assign n3026 = n3025 ^ n3024;
  assign n3023 = x244 ^ x243;
  assign n3027 = n3026 ^ n3023;
  assign n3029 = x240 ^ x239;
  assign n3031 = n3030 ^ n3029;
  assign n3028 = x238 ^ x237;
  assign n3032 = n3031 ^ n3028;
  assign n4971 = n3027 & n3032;
  assign n5036 = n5035 ^ n4971;
  assign n5090 = n5089 ^ n5036;
  assign n3022 = n3021 ^ n3016;
  assign n3033 = n3032 ^ n3027;
  assign n4837 = n3022 & n3033;
  assign n6514 = n5036 ^ n4837;
  assign n6515 = n5090 & ~n6514;
  assign n6516 = n6515 ^ n5089;
  assign n6517 = n5006 ^ n4971;
  assign n6518 = n5035 & ~n6517;
  assign n6519 = n6518 ^ n5034;
  assign n6911 = ~n6516 & ~n6519;
  assign n6528 = n5047 & ~n5060;
  assign n6527 = n5072 & ~n5085;
  assign n6529 = n6528 ^ n6527;
  assign n6524 = n5062 ^ n5037;
  assign n6525 = n5088 & ~n6524;
  assign n6526 = n6525 ^ n5087;
  assign n6530 = n6529 ^ n6526;
  assign n6522 = n6521 ^ n6520;
  assign n6523 = n6522 ^ n6519;
  assign n6531 = n6530 ^ n6523;
  assign n6532 = n6531 ^ n6516;
  assign n6913 = ~n6519 & ~n6530;
  assign n6914 = ~n6532 & ~n6913;
  assign n6916 = ~n6914 & ~n6915;
  assign n6912 = n6520 & n6521;
  assign n6917 = n6916 ^ n6912;
  assign n6918 = n6916 ^ n6530;
  assign n6919 = ~n6917 & n6918;
  assign n6920 = n6919 ^ n6916;
  assign n6921 = ~n6911 & n6920;
  assign n6922 = n6921 ^ n6916;
  assign n6908 = n6528 ^ n6526;
  assign n6909 = ~n6529 & ~n6908;
  assign n6910 = n6909 ^ n6526;
  assign n6923 = n6922 ^ n6910;
  assign n7356 = ~n6915 & ~n6923;
  assign n7357 = ~n6910 & ~n6914;
  assign n7358 = ~n7356 & ~n7357;
  assign n4943 = x251 & x252;
  assign n4944 = x249 & x250;
  assign n4945 = ~n4943 & ~n4944;
  assign n4946 = ~x251 & ~x252;
  assign n4947 = ~x249 & ~x250;
  assign n4948 = ~n4946 & ~n4947;
  assign n4949 = ~n4945 & n4948;
  assign n4950 = x248 & n4949;
  assign n4951 = n4943 & n4944;
  assign n4952 = ~n4950 & ~n4951;
  assign n4959 = n4949 ^ x248;
  assign n4960 = n4959 ^ n4949;
  assign n4953 = n4945 & ~n4948;
  assign n4961 = ~n4951 & ~n4953;
  assign n4962 = n4961 ^ n4949;
  assign n4963 = n4960 & n4962;
  assign n4964 = n4963 ^ n4949;
  assign n4965 = x247 & n4964;
  assign n6500 = n4952 & ~n4965;
  assign n4918 = x257 & x258;
  assign n4919 = x255 & x256;
  assign n4920 = ~n4918 & ~n4919;
  assign n4921 = ~x257 & ~x258;
  assign n4922 = ~x255 & ~x256;
  assign n4923 = ~n4921 & ~n4922;
  assign n4924 = ~n4920 & n4923;
  assign n4925 = x254 & n4924;
  assign n4926 = n4918 & n4919;
  assign n4927 = ~n4925 & ~n4926;
  assign n4934 = n4924 ^ x254;
  assign n4935 = n4934 ^ n4924;
  assign n4928 = n4920 & ~n4923;
  assign n4936 = ~n4926 & ~n4928;
  assign n4937 = n4936 ^ n4924;
  assign n4938 = n4935 & n4937;
  assign n4939 = n4938 ^ n4924;
  assign n4940 = x253 & n4939;
  assign n6499 = n4927 & ~n4940;
  assign n6501 = n6500 ^ n6499;
  assign n4954 = ~x248 & n4953;
  assign n4955 = n4952 & ~n4954;
  assign n4956 = ~x247 & ~n4955;
  assign n3007 = x248 ^ x247;
  assign n4957 = n4946 & n4947;
  assign n4958 = n3007 & n4957;
  assign n4966 = ~n4958 & ~n4965;
  assign n4967 = ~n4956 & n4966;
  assign n4929 = ~x254 & n4928;
  assign n4930 = n4927 & ~n4929;
  assign n4931 = ~x253 & ~n4930;
  assign n3002 = x254 ^ x253;
  assign n4932 = n4921 & n4922;
  assign n4933 = n3002 & n4932;
  assign n4941 = ~n4933 & ~n4940;
  assign n4942 = ~n4931 & n4941;
  assign n4968 = n4967 ^ n4942;
  assign n3001 = x256 ^ x255;
  assign n3003 = n3002 ^ n3001;
  assign n3000 = x258 ^ x257;
  assign n3004 = n3003 ^ n3000;
  assign n3006 = x250 ^ x249;
  assign n3008 = n3007 ^ n3006;
  assign n3005 = x252 ^ x251;
  assign n3009 = n3008 ^ n3005;
  assign n6495 = n3004 & n3009;
  assign n6496 = n6495 ^ n4942;
  assign n6497 = n4968 & ~n6496;
  assign n6498 = n6497 ^ n4967;
  assign n6502 = n6501 ^ n6498;
  assign n4868 = x269 & x270;
  assign n4867 = x267 & x268;
  assign n4869 = n4868 ^ n4867;
  assign n4870 = ~x269 & ~x270;
  assign n4871 = ~x267 & ~x268;
  assign n4872 = ~n4870 & ~n4871;
  assign n4873 = n4872 ^ n4867;
  assign n4874 = n4873 ^ n4867;
  assign n4875 = n4867 ^ x266;
  assign n4876 = n4875 ^ n4867;
  assign n4877 = n4874 & n4876;
  assign n4878 = n4877 ^ n4867;
  assign n4879 = n4869 & ~n4878;
  assign n4880 = n4879 ^ n4868;
  assign n4881 = n4871 ^ n4870;
  assign n4882 = ~n4867 & ~n4868;
  assign n4883 = n4882 ^ n4871;
  assign n4884 = n4883 ^ n4871;
  assign n4885 = n4871 ^ x266;
  assign n4886 = n4885 ^ n4871;
  assign n4887 = n4884 & ~n4886;
  assign n4888 = n4887 ^ n4871;
  assign n4889 = n4881 & ~n4888;
  assign n4890 = n4889 ^ n4870;
  assign n4891 = ~n4880 & ~n4890;
  assign n4892 = ~x265 & ~n4891;
  assign n2996 = x266 ^ x265;
  assign n4893 = n4872 & ~n4882;
  assign n4894 = n2996 & n4893;
  assign n4895 = ~n4872 & n4882;
  assign n4896 = x265 & x266;
  assign n4897 = n4867 & n4896;
  assign n4898 = x270 & n4897;
  assign n4899 = n4898 ^ n4896;
  assign n4900 = ~n4895 & n4899;
  assign n4901 = ~n4894 & ~n4900;
  assign n2995 = x268 ^ x267;
  assign n4902 = n4896 ^ x268;
  assign n4903 = n4902 ^ n4896;
  assign n4904 = ~x266 & ~x270;
  assign n4905 = n4904 ^ n4896;
  assign n4906 = ~n4903 & n4905;
  assign n4907 = n4906 ^ n4896;
  assign n4908 = ~n2995 & n4907;
  assign n4909 = ~x269 & n4908;
  assign n4910 = n4901 & ~n4909;
  assign n4911 = ~n4892 & n4910;
  assign n4840 = x263 & x264;
  assign n4841 = ~x261 & ~x262;
  assign n4842 = ~n4840 & n4841;
  assign n4843 = ~x263 & ~x264;
  assign n4844 = x260 & ~n4843;
  assign n4845 = n4842 & ~n4844;
  assign n4846 = x261 & x262;
  assign n4847 = n4840 & n4846;
  assign n4848 = ~n4845 & ~n4847;
  assign n4849 = ~x259 & ~n4848;
  assign n2991 = x260 ^ x259;
  assign n2990 = x262 ^ x261;
  assign n2992 = n2991 ^ n2990;
  assign n4850 = ~x260 & n4843;
  assign n4851 = ~n4846 & n4850;
  assign n4852 = n2992 & n4851;
  assign n4853 = x259 & x260;
  assign n4854 = n4846 & n4853;
  assign n4855 = ~n4840 & n4854;
  assign n4856 = ~n4852 & ~n4855;
  assign n4857 = ~n4849 & n4856;
  assign n4858 = ~n4846 & n4853;
  assign n4859 = ~n4842 & n4858;
  assign n4860 = n4840 ^ x262;
  assign n4861 = n2990 & n4860;
  assign n4862 = n4861 ^ x262;
  assign n4863 = n2991 & n4862;
  assign n4864 = ~n4859 & ~n4863;
  assign n4865 = ~n4843 & ~n4864;
  assign n4866 = n4857 & ~n4865;
  assign n4912 = n4911 ^ n4866;
  assign n2989 = x264 ^ x263;
  assign n2993 = n2992 ^ n2989;
  assign n2997 = n2996 ^ n2995;
  assign n2994 = x270 ^ x269;
  assign n2998 = n2997 ^ n2994;
  assign n6490 = n2993 & n2998;
  assign n6491 = n4912 & n6490;
  assign n6492 = n4866 & n4911;
  assign n6493 = ~n6491 & ~n6492;
  assign n6901 = n6502 ^ n6493;
  assign n4913 = n3004 ^ n2998;
  assign n4915 = n4913 ^ n2993;
  assign n4916 = ~n3009 & n4915;
  assign n2999 = n2998 ^ n2993;
  assign n4914 = ~n2999 & ~n4913;
  assign n4917 = n4916 ^ n4914;
  assign n4969 = n4968 ^ n4917;
  assign n4970 = n4969 ^ n4912;
  assign n6504 = n4968 & ~n6495;
  assign n6505 = ~n4970 & ~n6504;
  assign n3010 = n3009 ^ n3004;
  assign n6506 = ~n2993 & ~n2998;
  assign n6507 = n3010 & ~n6506;
  assign n6508 = ~n6490 & ~n6507;
  assign n6509 = n6508 ^ n6490;
  assign n6510 = ~n4912 & n6509;
  assign n6511 = n6510 ^ n6490;
  assign n6512 = ~n6505 & ~n6511;
  assign n6902 = n6512 ^ n6502;
  assign n6903 = n6901 & n6902;
  assign n6904 = n6903 ^ n6512;
  assign n6898 = n6500 ^ n6498;
  assign n6899 = ~n6501 & ~n6898;
  assign n6900 = n6899 ^ n6498;
  assign n6905 = n6904 ^ n6900;
  assign n6487 = ~n4847 & ~n4854;
  assign n6488 = ~n4865 & n6487;
  assign n6486 = ~n4880 & n4901;
  assign n6489 = n6488 ^ n6486;
  assign n6494 = n6493 ^ n6489;
  assign n6503 = n6502 ^ n6494;
  assign n6513 = n6512 ^ n6503;
  assign n6895 = n6513 ^ n6486;
  assign n6896 = n6489 & n6895;
  assign n6897 = n6896 ^ n6488;
  assign n7353 = n6900 ^ n6897;
  assign n7354 = n6905 & n7353;
  assign n7355 = n7354 ^ n6904;
  assign n7359 = n7358 ^ n7355;
  assign n6906 = n6905 ^ n6897;
  assign n3011 = n3010 ^ n2999;
  assign n3034 = n3033 ^ n3022;
  assign n4838 = n3011 & n3034;
  assign n5091 = n5090 ^ n4970;
  assign n4839 = ~n4837 & ~n4838;
  assign n5092 = n5091 ^ n4839;
  assign n6534 = ~n4838 & n5092;
  assign n6535 = ~n4837 & n5090;
  assign n6536 = n4970 & ~n6535;
  assign n6537 = ~n6534 & ~n6536;
  assign n6891 = n6537 ^ n6532;
  assign n6892 = n6537 ^ n6513;
  assign n6893 = n6891 & n6892;
  assign n6894 = n6893 ^ n6532;
  assign n6907 = n6906 ^ n6894;
  assign n7350 = n6923 ^ n6894;
  assign n7351 = n6907 & ~n7350;
  assign n7352 = n7351 ^ n6923;
  assign n7360 = n7359 ^ n7352;
  assign n7592 = n7591 ^ n7360;
  assign n7572 = n7345 & n7347;
  assign n7573 = ~n7343 & ~n7572;
  assign n7593 = ~n7568 & ~n7573;
  assign n7594 = n7593 ^ n7591;
  assign n6962 = n6961 ^ n6927;
  assign n6924 = n6923 ^ n6907;
  assign n6963 = n6962 ^ n6924;
  assign n6588 = n6587 ^ n6567;
  assign n6533 = n6532 ^ n6513;
  assign n6538 = n6537 ^ n6533;
  assign n6589 = n6588 ^ n6538;
  assign n3035 = n3034 ^ n3011;
  assign n3082 = n3081 ^ n3058;
  assign n4528 = n3035 & n3082;
  assign n4836 = n4835 ^ n4691;
  assign n5093 = n5092 ^ n4836;
  assign n6590 = ~n4528 & ~n5093;
  assign n6591 = n3011 & n3082;
  assign n6592 = n6590 & ~n6591;
  assign n6593 = n4836 & ~n4837;
  assign n6594 = ~n6592 & ~n6593;
  assign n6595 = n5091 & ~n6594;
  assign n6596 = n4836 ^ n4528;
  assign n6597 = ~n4839 & ~n5091;
  assign n6598 = n6597 ^ n4528;
  assign n6599 = ~n6596 & n6598;
  assign n6600 = n6599 ^ n4836;
  assign n6601 = ~n6595 & ~n6600;
  assign n6888 = n6601 ^ n6588;
  assign n6889 = ~n6589 & ~n6888;
  assign n6890 = n6889 ^ n6601;
  assign n7338 = n6924 ^ n6890;
  assign n7339 = n6963 & ~n7338;
  assign n7340 = n7339 ^ n6962;
  assign n7595 = n7360 ^ n7340;
  assign n7596 = n7595 ^ n7593;
  assign n7597 = n7593 & n7596;
  assign n7598 = n7597 ^ n7593;
  assign n7599 = ~n7594 & n7598;
  assign n7600 = n7599 ^ n7597;
  assign n7601 = n7600 ^ n7593;
  assign n7602 = n7601 ^ n7595;
  assign n7603 = n7592 & n7602;
  assign n7604 = n7603 ^ n7591;
  assign n7564 = n7355 ^ n7352;
  assign n7565 = n7359 & n7564;
  assign n7566 = n7565 ^ n7358;
  assign n7563 = n7340 & ~n7360;
  assign n7567 = ~n7563 & ~n7566;
  assign n7348 = n7347 ^ n7345;
  assign n7569 = n7343 & ~n7348;
  assign n7570 = ~n7568 & ~n7569;
  assign n7571 = ~n7567 & n7570;
  assign n7349 = n7348 ^ n7343;
  assign n7361 = n7360 ^ n7349;
  assign n7362 = n7361 ^ n7340;
  assign n7574 = ~n7362 & n7573;
  assign n7575 = n7571 & ~n7574;
  assign n7576 = n7347 & n7358;
  assign n7577 = n6941 & n7355;
  assign n7578 = ~n7576 & ~n7577;
  assign n7579 = n7345 & ~n7578;
  assign n7580 = n7352 & n7579;
  assign n7581 = n7355 & n7358;
  assign n7582 = n7581 ^ n7345;
  assign n7583 = n7582 ^ n7345;
  assign n7584 = n7572 ^ n7345;
  assign n7585 = ~n7583 & ~n7584;
  assign n7586 = n7585 ^ n7345;
  assign n7587 = ~n7352 & ~n7586;
  assign n7588 = ~n7580 & ~n7587;
  assign n7589 = n7343 & ~n7588;
  assign n7590 = ~n7575 & ~n7589;
  assign n7699 = ~n7566 & n7590;
  assign n7700 = ~n7604 & ~n7699;
  assign n3250 = x281 & x282;
  assign n3251 = ~x279 & ~x280;
  assign n3252 = ~n3250 & n3251;
  assign n3253 = x279 & x280;
  assign n3254 = x277 & x278;
  assign n3255 = ~n3253 & n3254;
  assign n3256 = ~n3252 & n3255;
  assign n2900 = x278 ^ x277;
  assign n2898 = x280 ^ x279;
  assign n3257 = n3250 ^ x280;
  assign n3258 = n2898 & n3257;
  assign n3259 = n3258 ^ x280;
  assign n3260 = n2900 & n3259;
  assign n3261 = ~n3256 & ~n3260;
  assign n3262 = ~x281 & ~x282;
  assign n3263 = ~n3261 & ~n3262;
  assign n3267 = n3253 & n3254;
  assign n3273 = n3250 & n3253;
  assign n6302 = ~n3267 & ~n3273;
  assign n6303 = ~n3263 & n6302;
  assign n2895 = x290 ^ x289;
  assign n3220 = x291 & x292;
  assign n3221 = x293 & x294;
  assign n3222 = ~n3220 & ~n3221;
  assign n3223 = ~x291 & ~x292;
  assign n3224 = ~x293 & ~x294;
  assign n3225 = ~n3223 & ~n3224;
  assign n3226 = n3222 & ~n3225;
  assign n3227 = ~n2895 & n3226;
  assign n3228 = n3220 & n3221;
  assign n3229 = n3223 & n3224;
  assign n3230 = ~n3228 & ~n3229;
  assign n3231 = ~n3227 & n3230;
  assign n3232 = x289 & x290;
  assign n3233 = ~n3231 & ~n3232;
  assign n3234 = ~n3228 & n3232;
  assign n3235 = n3234 ^ n3225;
  assign n3236 = n3234 ^ n2895;
  assign n3237 = n3225 ^ n3222;
  assign n3238 = n3237 ^ n3234;
  assign n3239 = ~n3234 & ~n3238;
  assign n3240 = n3239 ^ n3234;
  assign n3241 = n3236 & ~n3240;
  assign n3242 = n3241 ^ n3239;
  assign n3243 = n3242 ^ n3234;
  assign n3244 = n3243 ^ n3237;
  assign n3245 = n3235 & ~n3244;
  assign n3246 = n3245 ^ n3234;
  assign n3247 = ~n3233 & ~n3246;
  assign n2911 = x284 ^ x283;
  assign n3192 = ~x285 & ~x286;
  assign n3193 = ~x287 & ~x288;
  assign n3194 = ~n3192 & ~n3193;
  assign n3195 = x285 & x286;
  assign n3196 = x287 & x288;
  assign n3197 = ~n3195 & ~n3196;
  assign n3198 = ~n3194 & n3197;
  assign n3199 = ~n2911 & n3198;
  assign n3200 = n3195 & n3196;
  assign n3201 = n3192 & n3193;
  assign n3202 = ~n3200 & ~n3201;
  assign n3203 = ~n3199 & n3202;
  assign n3204 = x283 & x284;
  assign n3205 = ~n3203 & ~n3204;
  assign n3206 = ~n3200 & n3204;
  assign n3207 = n3206 ^ n3197;
  assign n3208 = n3206 ^ n2911;
  assign n3209 = n3197 ^ n3194;
  assign n3210 = n3209 ^ n3206;
  assign n3211 = ~n3206 & ~n3210;
  assign n3212 = n3211 ^ n3206;
  assign n3213 = n3208 & ~n3212;
  assign n3214 = n3213 ^ n3211;
  assign n3215 = n3214 ^ n3206;
  assign n3216 = n3215 ^ n3209;
  assign n3217 = ~n3207 & ~n3216;
  assign n3218 = n3217 ^ n3206;
  assign n3219 = ~n3205 & ~n3218;
  assign n3248 = n3247 ^ n3219;
  assign n2894 = x292 ^ x291;
  assign n2896 = n2895 ^ n2894;
  assign n2893 = x294 ^ x293;
  assign n2897 = n2896 ^ n2893;
  assign n2910 = x286 ^ x285;
  assign n2912 = n2911 ^ n2910;
  assign n2909 = x288 ^ x287;
  assign n2913 = n2912 ^ n2909;
  assign n6304 = n2897 & n2913;
  assign n6319 = n3248 & n6304;
  assign n3277 = ~x275 & ~x276;
  assign n3278 = x272 & ~n3277;
  assign n3279 = x275 & x276;
  assign n3280 = ~x273 & ~x274;
  assign n3281 = ~n3279 & n3280;
  assign n3282 = ~n3278 & n3281;
  assign n3283 = x273 & x274;
  assign n3284 = n3283 ^ n3279;
  assign n3285 = n3283 ^ n3278;
  assign n3286 = n3284 & n3285;
  assign n3287 = n3286 ^ n3283;
  assign n3288 = ~n3280 & n3287;
  assign n3289 = ~n3282 & ~n3288;
  assign n3290 = ~x271 & ~n3289;
  assign n3291 = ~n3279 & ~n3283;
  assign n3292 = ~n3280 & ~n3291;
  assign n3293 = x271 & ~n3277;
  assign n3294 = n3292 & n3293;
  assign n3295 = x271 & x272;
  assign n3296 = ~n3294 & ~n3295;
  assign n3297 = ~n3277 & ~n3283;
  assign n3298 = ~n3281 & n3297;
  assign n3299 = ~x276 & n3283;
  assign n3300 = x272 & ~n3299;
  assign n3301 = ~n3298 & n3300;
  assign n3302 = ~n3296 & ~n3301;
  assign n3303 = ~n3290 & ~n3302;
  assign n3304 = n3295 ^ n3283;
  assign n3305 = n3304 ^ n3295;
  assign n3306 = x271 & ~n3280;
  assign n3307 = ~x272 & ~x276;
  assign n3308 = ~n3306 & n3307;
  assign n3309 = n3308 ^ n3295;
  assign n3310 = ~n3305 & n3309;
  assign n3311 = n3310 ^ n3295;
  assign n3312 = ~x275 & n3311;
  assign n3313 = n3303 & ~n3312;
  assign n2899 = x282 ^ x281;
  assign n2901 = n2900 ^ n2899;
  assign n2902 = n2901 ^ n2898;
  assign n3264 = ~x278 & ~n3253;
  assign n3265 = n3262 & n3264;
  assign n3266 = n2902 & n3265;
  assign n3268 = ~n3250 & n3267;
  assign n3269 = ~n3266 & ~n3268;
  assign n3270 = ~n3263 & n3269;
  assign n3271 = x278 & ~n3262;
  assign n3272 = n3252 & ~n3271;
  assign n3274 = ~n3272 & ~n3273;
  assign n3275 = ~x277 & ~n3274;
  assign n3276 = n3270 & ~n3275;
  assign n3314 = n3313 ^ n3276;
  assign n2903 = n2902 ^ n2897;
  assign n2906 = x276 ^ x275;
  assign n2905 = x274 ^ x273;
  assign n2907 = n2906 ^ n2905;
  assign n2904 = x272 ^ x271;
  assign n2908 = n2907 ^ n2904;
  assign n2914 = n2913 ^ n2908;
  assign n3187 = n2903 & n2914;
  assign n3189 = n2908 & n2913;
  assign n3188 = n2897 & n2902;
  assign n3190 = n3189 ^ n3188;
  assign n3191 = ~n3187 & ~n3190;
  assign n6320 = ~n3191 & n3248;
  assign n6321 = n3188 & n3189;
  assign n6322 = ~n6320 & ~n6321;
  assign n6312 = n2902 & n2908;
  assign n6323 = n6322 ^ n6312;
  assign n6324 = n6323 ^ n6322;
  assign n6325 = n3191 & ~n3248;
  assign n6326 = n6325 ^ n6322;
  assign n6327 = n6326 ^ n6322;
  assign n6328 = ~n6324 & ~n6327;
  assign n6329 = n6328 ^ n6322;
  assign n6330 = n3314 & ~n6329;
  assign n6331 = n6330 ^ n6322;
  assign n6332 = ~n6319 & ~n6331;
  assign n6316 = ~n3288 & ~n3302;
  assign n6313 = n6312 ^ n3276;
  assign n6314 = n3314 & ~n6313;
  assign n6315 = n6314 ^ n3313;
  assign n6317 = n6316 ^ n6315;
  assign n6309 = ~n3200 & ~n3218;
  assign n6308 = ~n3228 & ~n3246;
  assign n6310 = n6309 ^ n6308;
  assign n6305 = n6304 ^ n3219;
  assign n6306 = n3248 & ~n6305;
  assign n6307 = n6306 ^ n3247;
  assign n6311 = n6310 ^ n6307;
  assign n6318 = n6317 ^ n6311;
  assign n6333 = n6332 ^ n6318;
  assign n7168 = n6303 & ~n6333;
  assign n7169 = n6332 ^ n6315;
  assign n7170 = n6317 & n7169;
  assign n7171 = n7170 ^ n6332;
  assign n7172 = n7168 & ~n7171;
  assign n7173 = ~n6315 & n6316;
  assign n7174 = ~n6311 & n7173;
  assign n7175 = ~n6332 & n7174;
  assign n7176 = ~n7172 & ~n7175;
  assign n7165 = n6309 ^ n6307;
  assign n7166 = ~n6310 & ~n7165;
  assign n7167 = n7166 ^ n6307;
  assign n6334 = n6333 ^ n6303;
  assign n7177 = n6311 & n7171;
  assign n7178 = ~n6334 & n7177;
  assign n7493 = ~n7167 & ~n7178;
  assign n7494 = n7176 & ~n7493;
  assign n3706 = x339 & x340;
  assign n3707 = x341 & x342;
  assign n3708 = ~n3706 & ~n3707;
  assign n3709 = ~x339 & ~x340;
  assign n3710 = ~x341 & ~x342;
  assign n3711 = ~n3709 & ~n3710;
  assign n3712 = ~n3708 & n3711;
  assign n3713 = x338 & n3712;
  assign n3714 = n3706 & n3707;
  assign n3715 = ~n3713 & ~n3714;
  assign n3722 = n3712 ^ x338;
  assign n3723 = n3722 ^ n3712;
  assign n3716 = n3708 & ~n3711;
  assign n3724 = ~n3714 & ~n3716;
  assign n3725 = n3724 ^ n3712;
  assign n3726 = n3723 & n3725;
  assign n3727 = n3726 ^ n3712;
  assign n3728 = x337 & n3727;
  assign n6247 = n3715 & ~n3728;
  assign n3680 = x335 & x336;
  assign n3681 = x333 & x334;
  assign n3682 = ~n3680 & ~n3681;
  assign n3683 = ~x335 & ~x336;
  assign n3684 = ~x333 & ~x334;
  assign n3685 = ~n3683 & ~n3684;
  assign n3686 = ~n3682 & n3685;
  assign n3687 = x332 & n3686;
  assign n3688 = n3680 & n3681;
  assign n3689 = ~n3687 & ~n3688;
  assign n3696 = n3686 ^ x332;
  assign n3697 = n3696 ^ n3686;
  assign n3690 = n3682 & ~n3685;
  assign n3698 = ~n3688 & ~n3690;
  assign n3699 = n3698 ^ n3686;
  assign n3700 = n3697 & n3699;
  assign n3701 = n3700 ^ n3686;
  assign n3702 = x331 & n3701;
  assign n6246 = n3689 & ~n3702;
  assign n6248 = n6247 ^ n6246;
  assign n3717 = ~x338 & n3716;
  assign n3718 = n3715 & ~n3717;
  assign n3719 = ~x337 & ~n3718;
  assign n2976 = x338 ^ x337;
  assign n3720 = n3709 & n3710;
  assign n3721 = n2976 & n3720;
  assign n3729 = ~n3721 & ~n3728;
  assign n3730 = ~n3719 & n3729;
  assign n2975 = x342 ^ x341;
  assign n2977 = n2976 ^ n2975;
  assign n2974 = x340 ^ x339;
  assign n2978 = n2977 ^ n2974;
  assign n2981 = x332 ^ x331;
  assign n2980 = x334 ^ x333;
  assign n2982 = n2981 ^ n2980;
  assign n2979 = x336 ^ x335;
  assign n2983 = n2982 ^ n2979;
  assign n3705 = n2978 & n2983;
  assign n3731 = n3730 ^ n3705;
  assign n3691 = ~x332 & n3690;
  assign n3692 = n3689 & ~n3691;
  assign n3693 = ~x331 & ~n3692;
  assign n3694 = n3683 & n3684;
  assign n3695 = n2981 & n3694;
  assign n3703 = ~n3695 & ~n3702;
  assign n3704 = ~n3693 & n3703;
  assign n6243 = n3705 ^ n3704;
  assign n6244 = n3731 & ~n6243;
  assign n6245 = n6244 ^ n3730;
  assign n7154 = n6247 ^ n6245;
  assign n7155 = ~n6248 & ~n7154;
  assign n7156 = n7155 ^ n6245;
  assign n3734 = x323 & x324;
  assign n3733 = x321 & x322;
  assign n3735 = n3734 ^ n3733;
  assign n3736 = ~x323 & ~x324;
  assign n3737 = ~x321 & ~x322;
  assign n3738 = ~n3736 & ~n3737;
  assign n3739 = n3738 ^ n3733;
  assign n3740 = n3739 ^ n3733;
  assign n3741 = n3733 ^ x320;
  assign n3742 = n3741 ^ n3733;
  assign n3743 = n3740 & n3742;
  assign n3744 = n3743 ^ n3733;
  assign n3745 = n3735 & ~n3744;
  assign n3746 = n3745 ^ n3734;
  assign n2970 = x320 ^ x319;
  assign n3748 = ~n3733 & ~n3734;
  assign n3759 = n3738 & ~n3748;
  assign n3760 = n2970 & n3759;
  assign n3761 = ~n3738 & n3748;
  assign n3762 = x319 & x320;
  assign n3763 = n3733 & n3762;
  assign n3764 = x324 & n3763;
  assign n3765 = n3764 ^ n3762;
  assign n3766 = ~n3761 & n3765;
  assign n3767 = ~n3760 & ~n3766;
  assign n6240 = ~n3746 & n3767;
  assign n3780 = x329 & x330;
  assign n3779 = x327 & x328;
  assign n3781 = n3780 ^ n3779;
  assign n3782 = ~x329 & ~x330;
  assign n3783 = ~x327 & ~x328;
  assign n3784 = ~n3782 & ~n3783;
  assign n3785 = n3784 ^ n3779;
  assign n3786 = n3785 ^ n3779;
  assign n3787 = n3779 ^ x326;
  assign n3788 = n3787 ^ n3779;
  assign n3789 = n3786 & n3788;
  assign n3790 = n3789 ^ n3779;
  assign n3791 = n3781 & ~n3790;
  assign n3792 = n3791 ^ n3780;
  assign n2965 = x326 ^ x325;
  assign n3794 = ~n3779 & ~n3780;
  assign n3805 = n3784 & ~n3794;
  assign n3806 = n2965 & n3805;
  assign n3807 = ~n3784 & n3794;
  assign n3808 = x325 & x326;
  assign n3809 = n3779 & n3808;
  assign n3810 = x330 & n3809;
  assign n3811 = n3810 ^ n3808;
  assign n3812 = ~n3807 & n3811;
  assign n3813 = ~n3806 & ~n3812;
  assign n6239 = ~n3792 & n3813;
  assign n6241 = n6240 ^ n6239;
  assign n3793 = n3783 ^ n3782;
  assign n3795 = n3794 ^ n3783;
  assign n3796 = n3795 ^ n3783;
  assign n3797 = n3783 ^ x326;
  assign n3798 = n3797 ^ n3783;
  assign n3799 = n3796 & ~n3798;
  assign n3800 = n3799 ^ n3783;
  assign n3801 = n3793 & ~n3800;
  assign n3802 = n3801 ^ n3782;
  assign n3803 = ~n3792 & ~n3802;
  assign n3804 = ~x325 & ~n3803;
  assign n2964 = x328 ^ x327;
  assign n3814 = n3808 ^ x328;
  assign n3815 = n3814 ^ n3808;
  assign n3816 = ~x326 & ~x330;
  assign n3817 = n3816 ^ n3808;
  assign n3818 = ~n3815 & n3817;
  assign n3819 = n3818 ^ n3808;
  assign n3820 = ~n2964 & n3819;
  assign n3821 = ~x329 & n3820;
  assign n3822 = n3813 & ~n3821;
  assign n3823 = ~n3804 & n3822;
  assign n2966 = n2965 ^ n2964;
  assign n2963 = x330 ^ x329;
  assign n2967 = n2966 ^ n2963;
  assign n2969 = x322 ^ x321;
  assign n2971 = n2970 ^ n2969;
  assign n2968 = x324 ^ x323;
  assign n2972 = n2971 ^ n2968;
  assign n3778 = n2967 & n2972;
  assign n3824 = n3823 ^ n3778;
  assign n3747 = n3737 ^ n3736;
  assign n3749 = n3748 ^ n3737;
  assign n3750 = n3749 ^ n3737;
  assign n3751 = n3737 ^ x320;
  assign n3752 = n3751 ^ n3737;
  assign n3753 = n3750 & ~n3752;
  assign n3754 = n3753 ^ n3737;
  assign n3755 = n3747 & ~n3754;
  assign n3756 = n3755 ^ n3736;
  assign n3757 = ~n3746 & ~n3756;
  assign n3758 = ~x319 & ~n3757;
  assign n3768 = n3762 ^ x322;
  assign n3769 = n3768 ^ n3762;
  assign n3770 = ~x320 & ~x324;
  assign n3771 = n3770 ^ n3762;
  assign n3772 = ~n3769 & n3771;
  assign n3773 = n3772 ^ n3762;
  assign n3774 = ~n2969 & n3773;
  assign n3775 = ~x323 & n3774;
  assign n3776 = n3767 & ~n3775;
  assign n3777 = ~n3758 & n3776;
  assign n6236 = n3778 ^ n3777;
  assign n6237 = n3824 & ~n6236;
  assign n6238 = n6237 ^ n3823;
  assign n7151 = n6240 ^ n6238;
  assign n7152 = ~n6241 & ~n7151;
  assign n7153 = n7152 ^ n6238;
  assign n7157 = n7156 ^ n7153;
  assign n6249 = n6248 ^ n6245;
  assign n6242 = n6241 ^ n6238;
  assign n6250 = n6249 ^ n6242;
  assign n3825 = n3824 ^ n3777;
  assign n3732 = n3731 ^ n3704;
  assign n3826 = n3825 ^ n3732;
  assign n2973 = n2972 ^ n2967;
  assign n2984 = n2983 ^ n2978;
  assign n3501 = n2973 & n2984;
  assign n6233 = n3732 ^ n3501;
  assign n6234 = n3826 & ~n6233;
  assign n6235 = n6234 ^ n3825;
  assign n7148 = n6242 ^ n6235;
  assign n7149 = n6250 & ~n7148;
  assign n7150 = n7149 ^ n6249;
  assign n7158 = n7157 ^ n7150;
  assign n2953 = x344 ^ x343;
  assign n2952 = x346 ^ x345;
  assign n3641 = x347 & x348;
  assign n3642 = n3641 ^ x346;
  assign n3643 = n2952 & ~n3642;
  assign n3644 = n3643 ^ x345;
  assign n3645 = n2953 & n3644;
  assign n3646 = ~x345 & ~x346;
  assign n3647 = ~n3641 & n3646;
  assign n3648 = x345 & x346;
  assign n3649 = x343 & x344;
  assign n3650 = ~n3648 & n3649;
  assign n3651 = ~n3647 & n3650;
  assign n3652 = ~n3645 & ~n3651;
  assign n3653 = ~x347 & ~x348;
  assign n3654 = ~n3652 & ~n3653;
  assign n3655 = n3648 & n3649;
  assign n3656 = ~x348 & n3655;
  assign n3657 = ~n3654 & ~n3656;
  assign n3658 = x344 & ~n3653;
  assign n3659 = n3641 & n3648;
  assign n3660 = ~n3658 & ~n3659;
  assign n3661 = n3644 & ~n3660;
  assign n6257 = n3657 & ~n3661;
  assign n3615 = ~x353 & ~x354;
  assign n3616 = ~x351 & ~x352;
  assign n3617 = ~n3615 & ~n3616;
  assign n3600 = x351 & x352;
  assign n3601 = x349 & x350;
  assign n3612 = n3600 & n3601;
  assign n3613 = x354 & n3612;
  assign n3614 = n3613 ^ n3601;
  assign n3618 = n3617 ^ n3614;
  assign n2958 = x350 ^ x349;
  assign n3619 = n3614 ^ n2958;
  assign n3620 = x353 & x354;
  assign n3621 = ~n3600 & ~n3620;
  assign n3622 = n3621 ^ n3617;
  assign n3623 = n3622 ^ n3614;
  assign n3624 = ~n3614 & ~n3623;
  assign n3625 = n3624 ^ n3614;
  assign n3626 = n3619 & ~n3625;
  assign n3627 = n3626 ^ n3624;
  assign n3628 = n3627 ^ n3614;
  assign n3629 = n3628 ^ n3622;
  assign n3630 = n3618 & ~n3629;
  assign n3631 = n3630 ^ n3614;
  assign n2956 = x354 ^ x353;
  assign n3633 = x353 ^ x350;
  assign n3634 = ~n2956 & n3633;
  assign n3635 = n3634 ^ x350;
  assign n6255 = n3600 & n3635;
  assign n6256 = ~n3631 & ~n6255;
  assign n6258 = n6257 ^ n6256;
  assign n2957 = x352 ^ x351;
  assign n2959 = n2958 ^ n2957;
  assign n3602 = n3601 ^ n2959;
  assign n3603 = n3602 ^ n3601;
  assign n3604 = ~x350 & ~x354;
  assign n3605 = n3604 ^ n3601;
  assign n3606 = n3605 ^ n3601;
  assign n3607 = n3603 & n3606;
  assign n3608 = n3607 ^ n3601;
  assign n3609 = ~n3600 & n3608;
  assign n3610 = n3609 ^ n3601;
  assign n3611 = ~x353 & n3610;
  assign n3632 = ~n3611 & ~n3631;
  assign n3636 = n3635 ^ x352;
  assign n3637 = ~n2957 & ~n3636;
  assign n3638 = ~x349 & n3637;
  assign n3639 = n3632 & ~n3638;
  assign n2954 = n2953 ^ n2952;
  assign n2951 = x348 ^ x347;
  assign n2955 = n2954 ^ n2951;
  assign n2960 = n2959 ^ n2956;
  assign n3599 = n2955 & n2960;
  assign n3640 = n3639 ^ n3599;
  assign n3662 = n3647 & ~n3658;
  assign n3663 = ~n3661 & ~n3662;
  assign n3664 = ~x343 & ~n3663;
  assign n3665 = n3657 & ~n3664;
  assign n3666 = ~x344 & ~x348;
  assign n3667 = n3666 ^ n3649;
  assign n3668 = n3667 ^ n3649;
  assign n3669 = n3649 ^ n2954;
  assign n3670 = n3669 ^ n3649;
  assign n3671 = n3668 & n3670;
  assign n3672 = n3671 ^ n3649;
  assign n3673 = ~n3648 & n3672;
  assign n3674 = n3673 ^ n3649;
  assign n3675 = ~x347 & n3674;
  assign n3676 = n3665 & ~n3675;
  assign n6252 = n3676 ^ n3639;
  assign n6253 = ~n3640 & n6252;
  assign n6254 = n6253 ^ n3676;
  assign n7143 = n6257 ^ n6254;
  assign n7144 = ~n6258 & ~n7143;
  assign n7145 = n7144 ^ n6254;
  assign n3508 = x365 & x366;
  assign n3507 = x363 & x364;
  assign n3509 = n3508 ^ n3507;
  assign n3510 = ~x365 & ~x366;
  assign n3511 = ~x363 & ~x364;
  assign n3512 = ~n3510 & ~n3511;
  assign n3513 = n3512 ^ n3507;
  assign n3514 = n3513 ^ n3507;
  assign n3515 = n3507 ^ x362;
  assign n3516 = n3515 ^ n3507;
  assign n3517 = n3514 & n3516;
  assign n3518 = n3517 ^ n3507;
  assign n3519 = n3509 & ~n3518;
  assign n3520 = n3519 ^ n3508;
  assign n2942 = x362 ^ x361;
  assign n3522 = ~n3507 & ~n3508;
  assign n3533 = n3512 & ~n3522;
  assign n3534 = n2942 & n3533;
  assign n3535 = ~n3512 & n3522;
  assign n3536 = x361 & x362;
  assign n3537 = n3507 & n3536;
  assign n3538 = x366 & n3537;
  assign n3539 = n3538 ^ n3536;
  assign n3540 = ~n3535 & n3539;
  assign n3541 = ~n3534 & ~n3540;
  assign n6267 = ~n3520 & n3541;
  assign n3553 = x359 & x360;
  assign n3552 = x357 & x358;
  assign n3554 = n3553 ^ n3552;
  assign n3555 = ~x359 & ~x360;
  assign n3556 = ~x357 & ~x358;
  assign n3557 = ~n3555 & ~n3556;
  assign n3558 = n3557 ^ n3552;
  assign n3559 = n3558 ^ n3552;
  assign n3560 = n3552 ^ x356;
  assign n3561 = n3560 ^ n3552;
  assign n3562 = n3559 & n3561;
  assign n3563 = n3562 ^ n3552;
  assign n3564 = n3554 & ~n3563;
  assign n3565 = n3564 ^ n3553;
  assign n2947 = x356 ^ x355;
  assign n3567 = ~n3552 & ~n3553;
  assign n3578 = n3557 & ~n3567;
  assign n3579 = n2947 & n3578;
  assign n3580 = ~n3557 & n3567;
  assign n3581 = x355 & x356;
  assign n3582 = n3552 & n3581;
  assign n3583 = x360 & n3582;
  assign n3584 = n3583 ^ n3581;
  assign n3585 = ~n3580 & n3584;
  assign n3586 = ~n3579 & ~n3585;
  assign n6266 = ~n3565 & n3586;
  assign n6268 = n6267 ^ n6266;
  assign n3566 = n3556 ^ n3555;
  assign n3568 = n3567 ^ n3556;
  assign n3569 = n3568 ^ n3556;
  assign n3570 = n3556 ^ x356;
  assign n3571 = n3570 ^ n3556;
  assign n3572 = n3569 & ~n3571;
  assign n3573 = n3572 ^ n3556;
  assign n3574 = n3566 & ~n3573;
  assign n3575 = n3574 ^ n3555;
  assign n3576 = ~n3565 & ~n3575;
  assign n3577 = ~x355 & ~n3576;
  assign n2946 = x358 ^ x357;
  assign n3587 = n3581 ^ x358;
  assign n3588 = n3587 ^ n3581;
  assign n3589 = ~x356 & ~x360;
  assign n3590 = n3589 ^ n3581;
  assign n3591 = ~n3588 & n3590;
  assign n3592 = n3591 ^ n3581;
  assign n3593 = ~n2946 & n3592;
  assign n3594 = ~x359 & n3593;
  assign n3595 = n3586 & ~n3594;
  assign n3596 = ~n3577 & n3595;
  assign n3521 = n3511 ^ n3510;
  assign n3523 = n3522 ^ n3511;
  assign n3524 = n3523 ^ n3511;
  assign n3525 = n3511 ^ x362;
  assign n3526 = n3525 ^ n3511;
  assign n3527 = n3524 & ~n3526;
  assign n3528 = n3527 ^ n3511;
  assign n3529 = n3521 & ~n3528;
  assign n3530 = n3529 ^ n3510;
  assign n3531 = ~n3520 & ~n3530;
  assign n3532 = ~x361 & ~n3531;
  assign n2941 = x364 ^ x363;
  assign n3542 = n3536 ^ x364;
  assign n3543 = n3542 ^ n3536;
  assign n3544 = ~x362 & ~x366;
  assign n3545 = n3544 ^ n3536;
  assign n3546 = ~n3543 & n3545;
  assign n3547 = n3546 ^ n3536;
  assign n3548 = ~n2941 & n3547;
  assign n3549 = ~x365 & n3548;
  assign n3550 = n3541 & ~n3549;
  assign n3551 = ~n3532 & n3550;
  assign n3597 = n3596 ^ n3551;
  assign n2943 = n2942 ^ n2941;
  assign n2940 = x366 ^ x365;
  assign n2944 = n2943 ^ n2940;
  assign n2948 = n2947 ^ n2946;
  assign n2945 = x360 ^ x359;
  assign n2949 = n2948 ^ n2945;
  assign n3504 = n2944 & n2949;
  assign n6263 = n3551 ^ n3504;
  assign n6264 = n3597 & ~n6263;
  assign n6265 = n6264 ^ n3596;
  assign n7140 = n6267 ^ n6265;
  assign n7141 = ~n6268 & ~n7140;
  assign n7142 = n7141 ^ n6265;
  assign n7146 = n7145 ^ n7142;
  assign n6269 = n6268 ^ n6265;
  assign n2950 = n2949 ^ n2944;
  assign n2961 = n2960 ^ n2955;
  assign n3505 = n2950 & n2961;
  assign n3506 = ~n3504 & ~n3505;
  assign n3598 = n3597 ^ n3506;
  assign n3677 = n3676 ^ n3640;
  assign n6260 = n3677 ^ n3505;
  assign n6261 = n3598 & n6260;
  assign n6262 = n6261 ^ n3677;
  assign n6270 = n6269 ^ n6262;
  assign n6259 = n6258 ^ n6254;
  assign n7137 = n6262 ^ n6259;
  assign n7138 = n6270 & ~n7137;
  assign n7139 = n7138 ^ n6269;
  assign n7147 = n7146 ^ n7139;
  assign n7159 = n7158 ^ n7147;
  assign n6271 = n6270 ^ n6259;
  assign n6251 = n6250 ^ n6235;
  assign n6272 = n6271 ^ n6251;
  assign n6228 = n3826 ^ n3501;
  assign n2962 = n2961 ^ n2950;
  assign n2985 = n2984 ^ n2973;
  assign n3502 = n2962 & n2985;
  assign n6229 = n6228 ^ n3502;
  assign n3678 = n3677 ^ n3598;
  assign n6230 = n3678 ^ n3502;
  assign n6231 = n6229 & n6230;
  assign n6232 = n6231 ^ n6228;
  assign n7134 = n6251 ^ n6232;
  assign n7135 = n6272 & ~n7134;
  assign n7136 = n7135 ^ n6271;
  assign n7160 = n7159 ^ n7136;
  assign n6273 = n6272 ^ n6232;
  assign n2929 = x314 ^ x313;
  assign n2928 = x316 ^ x315;
  assign n3461 = x317 & x318;
  assign n3462 = n3461 ^ x316;
  assign n3463 = n2928 & ~n3462;
  assign n3464 = n3463 ^ x315;
  assign n3465 = n2929 & n3464;
  assign n3466 = ~x315 & ~x316;
  assign n3467 = ~n3461 & n3466;
  assign n3468 = x315 & x316;
  assign n3469 = x313 & x314;
  assign n3470 = ~n3468 & n3469;
  assign n3471 = ~n3467 & n3470;
  assign n3472 = ~n3465 & ~n3471;
  assign n3473 = ~x317 & ~x318;
  assign n3474 = ~n3472 & ~n3473;
  assign n3475 = n3468 & n3469;
  assign n3476 = ~x318 & n3475;
  assign n3477 = ~n3474 & ~n3476;
  assign n3478 = x314 & ~n3473;
  assign n3479 = n3461 & n3468;
  assign n3480 = ~n3478 & ~n3479;
  assign n3481 = n3464 & ~n3480;
  assign n3482 = n3467 & ~n3478;
  assign n3483 = ~n3481 & ~n3482;
  assign n3484 = ~x313 & ~n3483;
  assign n3485 = n3477 & ~n3484;
  assign n3486 = ~x314 & ~x318;
  assign n3487 = n3486 ^ n3469;
  assign n3488 = n3487 ^ n3469;
  assign n2930 = n2929 ^ n2928;
  assign n3489 = n3469 ^ n2930;
  assign n3490 = n3489 ^ n3469;
  assign n3491 = n3488 & n3490;
  assign n3492 = n3491 ^ n3469;
  assign n3493 = ~n3468 & n3492;
  assign n3494 = n3493 ^ n3469;
  assign n3495 = ~x317 & n3494;
  assign n3496 = n3485 & ~n3495;
  assign n3422 = ~x311 & ~x312;
  assign n3423 = x308 & ~n3422;
  assign n3424 = x311 & x312;
  assign n3425 = ~x309 & ~x310;
  assign n3426 = ~n3424 & n3425;
  assign n3427 = ~n3423 & n3426;
  assign n3428 = x309 & x310;
  assign n3429 = n3428 ^ n3424;
  assign n3430 = n3428 ^ n3423;
  assign n3431 = n3429 & n3430;
  assign n3432 = n3431 ^ n3428;
  assign n3433 = ~n3425 & n3432;
  assign n3434 = ~n3427 & ~n3433;
  assign n3435 = ~x307 & ~n3434;
  assign n3436 = ~n3424 & ~n3428;
  assign n3437 = ~n3425 & ~n3436;
  assign n3438 = x307 & ~n3422;
  assign n3439 = n3437 & n3438;
  assign n3440 = x307 & x308;
  assign n3441 = ~n3439 & ~n3440;
  assign n3442 = ~n3422 & ~n3428;
  assign n3443 = ~n3426 & n3442;
  assign n3444 = ~x312 & n3428;
  assign n3445 = x308 & ~n3444;
  assign n3446 = ~n3443 & n3445;
  assign n3447 = ~n3441 & ~n3446;
  assign n3448 = ~n3435 & ~n3447;
  assign n3449 = ~x308 & ~x312;
  assign n3450 = n3449 ^ n3440;
  assign n3451 = n3450 ^ n3440;
  assign n3452 = x307 & ~n3425;
  assign n3453 = n3452 ^ n3440;
  assign n3454 = n3453 ^ n3440;
  assign n3455 = n3451 & ~n3454;
  assign n3456 = n3455 ^ n3440;
  assign n3457 = ~n3428 & n3456;
  assign n3458 = n3457 ^ n3440;
  assign n3459 = ~x311 & n3458;
  assign n3460 = n3448 & ~n3459;
  assign n3497 = n3496 ^ n3460;
  assign n3376 = x305 & x306;
  assign n3375 = x303 & x304;
  assign n3377 = n3376 ^ n3375;
  assign n3378 = ~x305 & ~x306;
  assign n3379 = ~x303 & ~x304;
  assign n3380 = ~n3378 & ~n3379;
  assign n3381 = n3380 ^ n3375;
  assign n3382 = n3381 ^ n3375;
  assign n3383 = n3375 ^ x302;
  assign n3384 = n3383 ^ n3375;
  assign n3385 = n3382 & n3384;
  assign n3386 = n3385 ^ n3375;
  assign n3387 = n3377 & ~n3386;
  assign n3388 = n3387 ^ n3376;
  assign n3389 = n3379 ^ n3378;
  assign n3390 = ~n3375 & ~n3376;
  assign n3391 = n3390 ^ n3379;
  assign n3392 = n3391 ^ n3379;
  assign n3393 = n3379 ^ x302;
  assign n3394 = n3393 ^ n3379;
  assign n3395 = n3392 & ~n3394;
  assign n3396 = n3395 ^ n3379;
  assign n3397 = n3389 & ~n3396;
  assign n3398 = n3397 ^ n3378;
  assign n3399 = ~n3388 & ~n3398;
  assign n3400 = ~x301 & ~n3399;
  assign n2923 = x302 ^ x301;
  assign n3401 = n3380 & ~n3390;
  assign n3402 = n2923 & n3401;
  assign n3403 = ~n3380 & n3390;
  assign n3404 = x301 & x302;
  assign n3405 = n3375 & n3404;
  assign n3406 = x306 & n3405;
  assign n3407 = n3406 ^ n3404;
  assign n3408 = ~n3403 & n3407;
  assign n3409 = ~n3402 & ~n3408;
  assign n2922 = x304 ^ x303;
  assign n3410 = n3404 ^ x304;
  assign n3411 = n3410 ^ n3404;
  assign n3412 = ~x302 & ~x306;
  assign n3413 = n3412 ^ n3404;
  assign n3414 = ~n3411 & n3413;
  assign n3415 = n3414 ^ n3404;
  assign n3416 = ~n2922 & n3415;
  assign n3417 = ~x305 & n3416;
  assign n3418 = n3409 & ~n3417;
  assign n3419 = ~n3400 & n3418;
  assign n2918 = x298 ^ x297;
  assign n3324 = x295 & x296;
  assign n3325 = n3324 ^ x298;
  assign n3326 = n3325 ^ n3324;
  assign n3327 = ~x296 & ~x300;
  assign n3328 = n3327 ^ n3324;
  assign n3329 = ~n3326 & n3328;
  assign n3330 = n3329 ^ n3324;
  assign n3331 = ~n2918 & n3330;
  assign n3332 = ~x299 & n3331;
  assign n3334 = x297 & x298;
  assign n3333 = x299 & x300;
  assign n3335 = n3334 ^ n3333;
  assign n3336 = ~x297 & ~x298;
  assign n3337 = ~x299 & ~x300;
  assign n3338 = ~n3336 & ~n3337;
  assign n3339 = n3338 ^ n3333;
  assign n3340 = n3339 ^ n3333;
  assign n3341 = n3333 ^ x296;
  assign n3342 = n3341 ^ n3333;
  assign n3343 = n3340 & n3342;
  assign n3344 = n3343 ^ n3333;
  assign n3345 = n3335 & ~n3344;
  assign n3346 = n3345 ^ n3334;
  assign n3347 = n3337 ^ n3336;
  assign n3348 = ~n3333 & ~n3334;
  assign n3349 = n3348 ^ n3337;
  assign n3350 = n3349 ^ n3337;
  assign n3351 = n3337 ^ x296;
  assign n3352 = n3351 ^ n3337;
  assign n3353 = n3350 & ~n3352;
  assign n3354 = n3353 ^ n3337;
  assign n3355 = n3347 & ~n3354;
  assign n3356 = n3355 ^ n3336;
  assign n3357 = ~n3346 & ~n3356;
  assign n3358 = n3357 ^ x295;
  assign n3359 = n3358 ^ n3357;
  assign n3361 = n3338 & ~n3348;
  assign n3360 = x300 & n3334;
  assign n3362 = n3361 ^ n3360;
  assign n3363 = n3362 ^ n3361;
  assign n3364 = ~n3338 & n3348;
  assign n3365 = n3364 ^ n3361;
  assign n3366 = n3365 ^ n3361;
  assign n3367 = ~n3363 & ~n3366;
  assign n3368 = n3367 ^ n3361;
  assign n3369 = x296 & n3368;
  assign n3370 = n3369 ^ n3361;
  assign n3371 = n3370 ^ n3357;
  assign n3372 = n3359 & ~n3371;
  assign n3373 = n3372 ^ n3357;
  assign n3374 = ~n3332 & n3373;
  assign n3420 = n3419 ^ n3374;
  assign n2927 = x318 ^ x317;
  assign n2931 = n2930 ^ n2927;
  assign n2934 = x312 ^ x311;
  assign n2933 = x310 ^ x309;
  assign n2935 = n2934 ^ n2933;
  assign n2932 = x308 ^ x307;
  assign n2936 = n2935 ^ n2932;
  assign n3316 = n2931 & n2936;
  assign n2917 = x300 ^ x299;
  assign n2919 = n2918 ^ n2917;
  assign n2916 = x296 ^ x295;
  assign n2920 = n2919 ^ n2916;
  assign n2924 = n2923 ^ n2922;
  assign n2921 = x306 ^ x305;
  assign n2925 = n2924 ^ n2921;
  assign n3320 = n2920 & n2925;
  assign n2926 = n2925 ^ n2920;
  assign n2937 = n2936 ^ n2931;
  assign n3317 = n2937 ^ n2925;
  assign n3318 = ~n2926 & n3317;
  assign n3319 = n3318 ^ n2937;
  assign n3321 = n3320 ^ n3319;
  assign n3322 = ~n3316 & ~n3321;
  assign n3323 = n3322 ^ n3320;
  assign n3421 = n3420 ^ n3323;
  assign n3498 = n3497 ^ n3421;
  assign n3249 = n3248 ^ n3191;
  assign n3315 = n3314 ^ n3249;
  assign n3499 = n3498 ^ n3315;
  assign n2915 = n2914 ^ n2903;
  assign n2938 = n2937 ^ n2926;
  assign n3184 = n2915 & n2938;
  assign n6218 = n3499 ^ n3184;
  assign n3503 = ~n3501 & ~n3502;
  assign n3679 = n3678 ^ n3503;
  assign n3827 = n3826 ^ n3679;
  assign n6219 = n6218 ^ n3827;
  assign n6220 = n3827 ^ n3184;
  assign n6221 = n6220 ^ n3827;
  assign n2939 = n2938 ^ n2915;
  assign n2986 = n2985 ^ n2962;
  assign n3185 = n2939 & n2986;
  assign n6222 = n3827 ^ n3185;
  assign n6223 = n6222 ^ n3827;
  assign n6224 = ~n6221 & n6223;
  assign n6225 = n6224 ^ n3827;
  assign n6226 = n6219 & n6225;
  assign n6227 = n6226 ^ n3827;
  assign n6274 = n6273 ^ n6227;
  assign n6299 = n3184 & n3499;
  assign n6300 = ~n3315 & ~n3498;
  assign n6301 = ~n6299 & ~n6300;
  assign n6335 = n6334 ^ n6301;
  assign n6290 = n3316 & n3497;
  assign n6291 = ~n3319 & ~n3420;
  assign n6292 = ~n6290 & ~n6291;
  assign n6293 = ~n3421 & ~n3497;
  assign n6294 = n3320 & n3420;
  assign n6295 = ~n6293 & ~n6294;
  assign n6296 = n6292 & n6295;
  assign n6285 = x295 & n3370;
  assign n6286 = ~n3346 & ~n6285;
  assign n6284 = ~n3388 & n3409;
  assign n6287 = n6286 ^ n6284;
  assign n6281 = n3374 ^ n3320;
  assign n6282 = n3420 & ~n6281;
  assign n6283 = n6282 ^ n3419;
  assign n6288 = n6287 ^ n6283;
  assign n6280 = n3477 & ~n3481;
  assign n6289 = n6288 ^ n6280;
  assign n6297 = n6296 ^ n6289;
  assign n6278 = ~n3433 & ~n3447;
  assign n6275 = n3460 ^ n3316;
  assign n6276 = n3497 & ~n6275;
  assign n6277 = n6276 ^ n3496;
  assign n6279 = n6278 ^ n6277;
  assign n6298 = n6297 ^ n6279;
  assign n6336 = n6335 ^ n6298;
  assign n7131 = n6336 ^ n6273;
  assign n7132 = ~n6274 & ~n7131;
  assign n7133 = n7132 ^ n6336;
  assign n7161 = n7160 ^ n7133;
  assign n7182 = n6286 ^ n6283;
  assign n7183 = ~n6287 & ~n7182;
  assign n7184 = n7183 ^ n6283;
  assign n7185 = n6280 & ~n6288;
  assign n7186 = ~n6296 & n7185;
  assign n7187 = n6277 & ~n6278;
  assign n7188 = n7186 & ~n7187;
  assign n7189 = n7184 & ~n7188;
  assign n7190 = ~n6280 & n6288;
  assign n7191 = n6296 & n7190;
  assign n7192 = ~n7189 & ~n7191;
  assign n7193 = n6296 ^ n6288;
  assign n7194 = n6289 & n7193;
  assign n7195 = n7194 ^ n6296;
  assign n7196 = n7187 & n7195;
  assign n7197 = n7192 & ~n7196;
  assign n7198 = ~n6277 & n6278;
  assign n7199 = ~n6297 & n7198;
  assign n7200 = ~n7197 & ~n7199;
  assign n7201 = n6288 & n6296;
  assign n7202 = n7200 & n7201;
  assign n7203 = n7195 ^ n6277;
  assign n7204 = n6279 & ~n7203;
  assign n7205 = ~n7188 & n7204;
  assign n7206 = n7205 ^ n7188;
  assign n7207 = ~n7202 & ~n7206;
  assign n7208 = n7207 ^ n7184;
  assign n7179 = n7176 & ~n7178;
  assign n7180 = n7179 ^ n7167;
  assign n7162 = n6301 ^ n6298;
  assign n7163 = ~n6335 & n7162;
  assign n7164 = n7163 ^ n6334;
  assign n7181 = n7180 ^ n7164;
  assign n7209 = n7208 ^ n7181;
  assign n7490 = n7209 ^ n7133;
  assign n7491 = n7161 & ~n7490;
  assign n7492 = n7491 ^ n7209;
  assign n7479 = n7153 & n7156;
  assign n7480 = n7150 & n7479;
  assign n7481 = n7139 & n7480;
  assign n7486 = n7208 ^ n7180;
  assign n7487 = ~n7181 & n7486;
  assign n7488 = n7487 ^ n7208;
  assign n7627 = ~n7200 & ~n7488;
  assign n7628 = ~n7481 & n7627;
  assign n7629 = ~n7492 & n7628;
  assign n7630 = ~n7494 & ~n7629;
  assign n7456 = n7156 ^ n7150;
  assign n7457 = ~n7157 & n7456;
  assign n7458 = n7457 ^ n7150;
  assign n7464 = ~n7142 & ~n7145;
  assign n7465 = ~n7136 & n7464;
  assign n7466 = n7465 ^ n7139;
  assign n7450 = n7145 ^ n7136;
  assign n7451 = ~n7146 & n7450;
  assign n7452 = n7451 ^ n7136;
  assign n7467 = n7465 ^ n7452;
  assign n7468 = n7158 ^ n7139;
  assign n7469 = n7468 ^ n7465;
  assign n7470 = ~n7465 & n7469;
  assign n7471 = n7470 ^ n7465;
  assign n7472 = ~n7467 & ~n7471;
  assign n7473 = n7472 ^ n7470;
  assign n7474 = n7473 ^ n7465;
  assign n7475 = n7474 ^ n7468;
  assign n7476 = ~n7466 & n7475;
  assign n7477 = n7476 ^ n7465;
  assign n7484 = ~n7458 & n7477;
  assign n7631 = n7200 & n7488;
  assign n7632 = n7484 & ~n7631;
  assign n7633 = n7492 & ~n7627;
  assign n7634 = n7632 & ~n7633;
  assign n7635 = n7630 & ~n7634;
  assign n7449 = n7139 & n7158;
  assign n7453 = n7449 & n7452;
  assign n7454 = n7142 & n7145;
  assign n7455 = n7136 & n7454;
  assign n7459 = ~n7455 & ~n7458;
  assign n7460 = ~n7153 & ~n7156;
  assign n7461 = ~n7150 & n7460;
  assign n7462 = ~n7459 & ~n7461;
  assign n7463 = ~n7453 & ~n7462;
  assign n7478 = ~n7463 & ~n7477;
  assign n7636 = n7492 & n7631;
  assign n7637 = ~n7478 & ~n7636;
  assign n7638 = ~n7627 & ~n7637;
  assign n7482 = n7452 & n7481;
  assign n7483 = n7478 & ~n7482;
  assign n7639 = n7483 & ~n7492;
  assign n7640 = ~n7631 & n7639;
  assign n7641 = n7638 & ~n7640;
  assign n7642 = n7635 & ~n7641;
  assign n7643 = ~n7478 & n7494;
  assign n7647 = ~n7492 & n7643;
  assign n7644 = n7643 ^ n7483;
  assign n7645 = n7492 & n7644;
  assign n7646 = n7645 ^ n7483;
  assign n7648 = n7647 ^ n7646;
  assign n7649 = n7647 ^ n7484;
  assign n7650 = n7488 ^ n7484;
  assign n7651 = ~n7484 & n7650;
  assign n7652 = n7651 ^ n7484;
  assign n7653 = ~n7649 & ~n7652;
  assign n7654 = n7653 ^ n7651;
  assign n7655 = n7654 ^ n7484;
  assign n7656 = n7655 ^ n7488;
  assign n7657 = n7648 & n7656;
  assign n7658 = n7657 ^ n7647;
  assign n7659 = ~n7200 & n7658;
  assign n7495 = n7494 ^ n7492;
  assign n7489 = n7488 ^ n7200;
  assign n7496 = n7495 ^ n7489;
  assign n7714 = ~n7484 & n7496;
  assign n7715 = ~n7478 & ~n7714;
  assign n7716 = ~n7659 & ~n7715;
  assign n7717 = ~n7642 & n7716;
  assign n7660 = n7200 & n7492;
  assign n7661 = n7488 & n7643;
  assign n7662 = ~n7660 & ~n7661;
  assign n7663 = n7484 & ~n7662;
  assign n7664 = n7647 ^ n7488;
  assign n7665 = n7664 ^ n7647;
  assign n7666 = n7482 & n7494;
  assign n7667 = n7666 ^ n7647;
  assign n7668 = n7665 & n7667;
  assign n7669 = n7668 ^ n7647;
  assign n7670 = n7200 & n7669;
  assign n7671 = ~n7663 & ~n7670;
  assign n7672 = ~n7659 & n7671;
  assign n7673 = ~n7642 & n7672;
  assign n4217 = x395 & x396;
  assign n4216 = x393 & x394;
  assign n4218 = n4217 ^ n4216;
  assign n4219 = ~x395 & ~x396;
  assign n4220 = ~x393 & ~x394;
  assign n4221 = ~n4219 & ~n4220;
  assign n4222 = n4221 ^ n4216;
  assign n4223 = n4222 ^ n4216;
  assign n4224 = n4216 ^ x392;
  assign n4225 = n4224 ^ n4216;
  assign n4226 = n4223 & n4225;
  assign n4227 = n4226 ^ n4216;
  assign n4228 = n4218 & ~n4227;
  assign n4229 = n4228 ^ n4217;
  assign n4230 = n4220 ^ n4219;
  assign n4231 = ~n4216 & ~n4217;
  assign n4232 = n4231 ^ n4220;
  assign n4233 = n4232 ^ n4220;
  assign n4234 = n4220 ^ x392;
  assign n4235 = n4234 ^ n4220;
  assign n4236 = n4233 & ~n4235;
  assign n4237 = n4236 ^ n4220;
  assign n4238 = n4230 & ~n4237;
  assign n4239 = n4238 ^ n4219;
  assign n4240 = ~n4229 & ~n4239;
  assign n4241 = ~x391 & ~n4240;
  assign n2875 = x392 ^ x391;
  assign n4242 = n4221 & ~n4231;
  assign n4243 = n2875 & n4242;
  assign n4244 = ~n4221 & n4231;
  assign n4245 = x391 & x392;
  assign n4246 = n4216 & n4245;
  assign n4247 = x396 & n4246;
  assign n4248 = n4247 ^ n4245;
  assign n4249 = ~n4244 & n4248;
  assign n4250 = ~n4243 & ~n4249;
  assign n2874 = x394 ^ x393;
  assign n4251 = n4245 ^ x394;
  assign n4252 = n4251 ^ n4245;
  assign n4253 = ~x392 & ~x396;
  assign n4254 = n4253 ^ n4245;
  assign n4255 = ~n4252 & n4254;
  assign n4256 = n4255 ^ n4245;
  assign n4257 = ~n2874 & n4256;
  assign n4258 = ~x395 & n4257;
  assign n4259 = n4250 & ~n4258;
  assign n4260 = ~n4241 & n4259;
  assign n4189 = x401 & x402;
  assign n4190 = ~x399 & ~x400;
  assign n4191 = ~n4189 & n4190;
  assign n4192 = ~x401 & ~x402;
  assign n4193 = x398 & ~n4192;
  assign n4194 = n4191 & ~n4193;
  assign n4195 = x399 & x400;
  assign n4196 = n4189 & n4195;
  assign n4197 = ~n4194 & ~n4196;
  assign n4198 = ~x397 & ~n4197;
  assign n2881 = x402 ^ x401;
  assign n2880 = x398 ^ x397;
  assign n2882 = n2881 ^ n2880;
  assign n2879 = x400 ^ x399;
  assign n2883 = n2882 ^ n2879;
  assign n4199 = ~x398 & n4192;
  assign n4200 = ~n4195 & n4199;
  assign n4201 = n2883 & n4200;
  assign n4202 = x397 & x398;
  assign n4203 = n4195 & n4202;
  assign n4204 = ~n4189 & n4203;
  assign n4205 = ~n4201 & ~n4204;
  assign n4206 = ~n4198 & n4205;
  assign n4207 = ~n4195 & n4202;
  assign n4208 = ~n4191 & n4207;
  assign n4209 = n4189 ^ x400;
  assign n4210 = n2879 & n4209;
  assign n4211 = n4210 ^ x400;
  assign n4212 = n2880 & n4211;
  assign n4213 = ~n4208 & ~n4212;
  assign n4214 = ~n4192 & ~n4213;
  assign n4215 = n4206 & ~n4214;
  assign n4261 = n4260 ^ n4215;
  assign n2876 = n2875 ^ n2874;
  assign n2873 = x396 ^ x395;
  assign n2877 = n2876 ^ n2873;
  assign n6171 = n2877 & n2883;
  assign n6172 = n4261 & n6171;
  assign n6173 = n4215 & n4260;
  assign n6174 = ~n6172 & ~n6173;
  assign n6169 = ~n4229 & n4250;
  assign n6167 = ~n4196 & ~n4203;
  assign n6168 = ~n4214 & n6167;
  assign n6170 = n6169 ^ n6168;
  assign n6175 = n6174 ^ n6170;
  assign n4303 = x407 & x408;
  assign n4302 = x405 & x406;
  assign n4304 = n4303 ^ n4302;
  assign n4305 = ~x407 & ~x408;
  assign n4306 = ~x405 & ~x406;
  assign n4307 = ~n4305 & ~n4306;
  assign n4308 = n4307 ^ n4302;
  assign n4309 = n4308 ^ n4302;
  assign n4310 = n4302 ^ x404;
  assign n4311 = n4310 ^ n4302;
  assign n4312 = n4309 & n4311;
  assign n4313 = n4312 ^ n4302;
  assign n4314 = n4304 & ~n4313;
  assign n4315 = n4314 ^ n4303;
  assign n2870 = x404 ^ x403;
  assign n4317 = ~n4302 & ~n4303;
  assign n4328 = n4307 & ~n4317;
  assign n4329 = n2870 & n4328;
  assign n4330 = ~n4307 & n4317;
  assign n4331 = x403 & x404;
  assign n4332 = n4302 & n4331;
  assign n4333 = x408 & n4332;
  assign n4334 = n4333 ^ n4331;
  assign n4335 = ~n4330 & n4334;
  assign n4336 = ~n4329 & ~n4335;
  assign n6162 = ~n4315 & n4336;
  assign n4272 = ~x413 & ~x414;
  assign n4273 = ~x411 & ~x412;
  assign n4274 = ~n4272 & ~n4273;
  assign n4275 = x410 & n4274;
  assign n4271 = x413 & x414;
  assign n4276 = n4275 ^ n4271;
  assign n4277 = x411 & x412;
  assign n4278 = n4277 ^ n4271;
  assign n4279 = n4276 & ~n4278;
  assign n4280 = n4279 ^ n4275;
  assign n2886 = x414 ^ x413;
  assign n2885 = x412 ^ x411;
  assign n2887 = n2886 ^ n2885;
  assign n2884 = x410 ^ x409;
  assign n2888 = n2887 ^ n2884;
  assign n4270 = x409 & ~n2888;
  assign n4282 = ~n4271 & ~n4277;
  assign n4295 = ~n4274 & n4282;
  assign n6163 = n4270 & ~n4295;
  assign n6164 = ~n4280 & ~n6163;
  assign n7091 = ~n6162 & ~n6164;
  assign n7092 = n6175 & ~n7091;
  assign n2869 = x406 ^ x405;
  assign n2871 = n2870 ^ n2869;
  assign n2868 = x408 ^ x407;
  assign n2872 = n2871 ^ n2868;
  assign n4263 = n2872 & n2877;
  assign n2889 = n2888 ^ n2883;
  assign n2878 = n2877 ^ n2872;
  assign n4265 = n2883 ^ n2878;
  assign n4266 = n2889 & n4265;
  assign n4267 = n4266 ^ n2883;
  assign n4268 = ~n4263 & ~n4267;
  assign n4316 = n4306 ^ n4305;
  assign n4318 = n4317 ^ n4306;
  assign n4319 = n4318 ^ n4306;
  assign n4320 = n4306 ^ x404;
  assign n4321 = n4320 ^ n4306;
  assign n4322 = n4319 & ~n4321;
  assign n4323 = n4322 ^ n4306;
  assign n4324 = n4316 & ~n4323;
  assign n4325 = n4324 ^ n4305;
  assign n4326 = ~n4315 & ~n4325;
  assign n4327 = ~x403 & ~n4326;
  assign n4337 = n4331 ^ x406;
  assign n4338 = n4337 ^ n4331;
  assign n4339 = ~x404 & ~x408;
  assign n4340 = n4339 ^ n4331;
  assign n4341 = ~n4338 & n4340;
  assign n4342 = n4341 ^ n4331;
  assign n4343 = ~n2869 & n4342;
  assign n4344 = ~x407 & n4343;
  assign n4345 = n4336 & ~n4344;
  assign n4346 = ~n4327 & n4345;
  assign n4292 = n4271 & n4277;
  assign n4281 = n4273 ^ n4272;
  assign n4283 = n4282 ^ n4273;
  assign n4284 = n4283 ^ n4273;
  assign n4285 = n4273 ^ x410;
  assign n4286 = n4285 ^ n4273;
  assign n4287 = n4284 & ~n4286;
  assign n4288 = n4287 ^ n4273;
  assign n4289 = n4281 & ~n4288;
  assign n4290 = n4289 ^ n4272;
  assign n4291 = ~n4280 & ~n4290;
  assign n4293 = n4292 ^ n4291;
  assign n4294 = n4293 ^ n4291;
  assign n4296 = n4295 ^ n4291;
  assign n4297 = n4296 ^ n4291;
  assign n4298 = ~n4294 & ~n4297;
  assign n4299 = n4298 ^ n4291;
  assign n4300 = n4270 & ~n4299;
  assign n4301 = n4300 ^ n4291;
  assign n4347 = n4346 ^ n4301;
  assign n6177 = n4268 & ~n4347;
  assign n6158 = n2872 & n2888;
  assign n6178 = n4347 & n6158;
  assign n4262 = n2883 & n2888;
  assign n4264 = n4262 & n4263;
  assign n4269 = ~n4264 & ~n4268;
  assign n4348 = n4347 ^ n4269;
  assign n4349 = n4348 ^ n4261;
  assign n6179 = n4349 ^ n4348;
  assign n6180 = n6171 ^ n4348;
  assign n6181 = n6179 & n6180;
  assign n6182 = n6181 ^ n4348;
  assign n6183 = ~n6178 & ~n6182;
  assign n6184 = ~n6177 & n6183;
  assign n6159 = n6158 ^ n4346;
  assign n6160 = n4347 & ~n6159;
  assign n6161 = n6160 ^ n4301;
  assign n7090 = n6184 ^ n6161;
  assign n7093 = n7092 ^ n6161;
  assign n7094 = n7093 ^ n7092;
  assign n7095 = n6162 & n6164;
  assign n7096 = ~n6175 & ~n7095;
  assign n7097 = n7096 ^ n7092;
  assign n7098 = n7094 & n7097;
  assign n7099 = n7098 ^ n7092;
  assign n7100 = ~n7090 & n7099;
  assign n7101 = ~n6161 & ~n6184;
  assign n7102 = ~n6175 & ~n7101;
  assign n7103 = n7102 ^ n7091;
  assign n7104 = n7103 ^ n7091;
  assign n6165 = n6164 ^ n6162;
  assign n6166 = n6165 ^ n6161;
  assign n6176 = n6175 ^ n6166;
  assign n6185 = n6184 ^ n6176;
  assign n7105 = ~n6185 & n7095;
  assign n7106 = n7105 ^ n7091;
  assign n7107 = ~n7104 & n7106;
  assign n7108 = n7107 ^ n7091;
  assign n7109 = ~n7100 & ~n7108;
  assign n7087 = n6174 ^ n6169;
  assign n7088 = ~n6170 & n7087;
  assign n7089 = n7088 ^ n6174;
  assign n7110 = n7109 ^ n7089;
  assign n7437 = n7092 & ~n7110;
  assign n7438 = n7091 & n7102;
  assign n7439 = n6161 & n6184;
  assign n7440 = n7089 & ~n7439;
  assign n7441 = ~n7438 & n7440;
  assign n7442 = ~n7105 & ~n7441;
  assign n7443 = ~n7437 & n7442;
  assign n4477 = x389 & x390;
  assign n4476 = x387 & x388;
  assign n4478 = n4477 ^ n4476;
  assign n4479 = ~x389 & ~x390;
  assign n4480 = ~x387 & ~x388;
  assign n4481 = ~n4479 & ~n4480;
  assign n4482 = n4481 ^ n4476;
  assign n4483 = n4482 ^ n4476;
  assign n4484 = n4476 ^ x386;
  assign n4485 = n4484 ^ n4476;
  assign n4486 = n4483 & n4485;
  assign n4487 = n4486 ^ n4476;
  assign n4488 = n4478 & ~n4487;
  assign n4489 = n4488 ^ n4477;
  assign n4490 = n4480 ^ n4479;
  assign n4491 = ~n4476 & ~n4477;
  assign n4492 = n4491 ^ n4480;
  assign n4493 = n4492 ^ n4480;
  assign n4494 = n4480 ^ x386;
  assign n4495 = n4494 ^ n4480;
  assign n4496 = n4493 & ~n4495;
  assign n4497 = n4496 ^ n4480;
  assign n4498 = n4490 & ~n4497;
  assign n4499 = n4498 ^ n4479;
  assign n4500 = ~n4489 & ~n4499;
  assign n4501 = ~x385 & ~n4500;
  assign n2863 = x386 ^ x385;
  assign n4502 = n4481 & ~n4491;
  assign n4503 = n2863 & n4502;
  assign n4504 = ~n4481 & n4491;
  assign n4505 = x385 & x386;
  assign n4506 = n4476 & n4505;
  assign n4507 = x390 & n4506;
  assign n4508 = n4507 ^ n4505;
  assign n4509 = ~n4504 & n4508;
  assign n4510 = ~n4503 & ~n4509;
  assign n2862 = x388 ^ x387;
  assign n4511 = n4505 ^ x388;
  assign n4512 = n4511 ^ n4505;
  assign n4513 = ~x386 & ~x390;
  assign n4514 = n4513 ^ n4505;
  assign n4515 = ~n4512 & n4514;
  assign n4516 = n4515 ^ n4505;
  assign n4517 = ~n2862 & n4516;
  assign n4518 = ~x389 & n4517;
  assign n4519 = n4510 & ~n4518;
  assign n4520 = ~n4501 & n4519;
  assign n4447 = ~x381 & ~x382;
  assign n4448 = ~x383 & ~x384;
  assign n4449 = ~n4447 & ~n4448;
  assign n4450 = x381 & x382;
  assign n4451 = x383 & x384;
  assign n4452 = ~n4450 & ~n4451;
  assign n4453 = ~n4449 & n4452;
  assign n4454 = ~x380 & n4453;
  assign n4455 = n4450 & n4451;
  assign n4456 = ~n4454 & ~n4455;
  assign n4457 = ~x379 & ~n4456;
  assign n4458 = x379 & x380;
  assign n4459 = n4447 & ~n4458;
  assign n4460 = n4448 & n4459;
  assign n4461 = ~n4455 & n4458;
  assign n4462 = n4461 ^ n4452;
  assign n2858 = x380 ^ x379;
  assign n4463 = n4461 ^ n2858;
  assign n4464 = n4452 ^ n4449;
  assign n4465 = n4464 ^ n4461;
  assign n4466 = ~n4461 & ~n4465;
  assign n4467 = n4466 ^ n4461;
  assign n4468 = n4463 & ~n4467;
  assign n4469 = n4468 ^ n4466;
  assign n4470 = n4469 ^ n4461;
  assign n4471 = n4470 ^ n4464;
  assign n4472 = ~n4462 & ~n4471;
  assign n4473 = n4472 ^ n4461;
  assign n4474 = ~n4460 & ~n4473;
  assign n4475 = ~n4457 & n4474;
  assign n4521 = n4520 ^ n4475;
  assign n2852 = x372 ^ x371;
  assign n2851 = x368 ^ x367;
  assign n2853 = n2852 ^ n2851;
  assign n2850 = x370 ^ x369;
  assign n2854 = n2853 ^ n2850;
  assign n2847 = x378 ^ x377;
  assign n2846 = x374 ^ x373;
  assign n2848 = n2847 ^ n2846;
  assign n2845 = x376 ^ x375;
  assign n2849 = n2848 ^ n2845;
  assign n2855 = n2854 ^ n2849;
  assign n2864 = n2863 ^ n2862;
  assign n2861 = x390 ^ x389;
  assign n2865 = n2864 ^ n2861;
  assign n2857 = x384 ^ x383;
  assign n2859 = n2858 ^ n2857;
  assign n2856 = x382 ^ x381;
  assign n2860 = n2859 ^ n2856;
  assign n2866 = n2865 ^ n2860;
  assign n4442 = n2855 & n2866;
  assign n4444 = n2860 & n2865;
  assign n4443 = n2849 & n2854;
  assign n4445 = n4444 ^ n4443;
  assign n4446 = ~n4442 & ~n4445;
  assign n4522 = n4521 ^ n4446;
  assign n4397 = x371 & x372;
  assign n4396 = x369 & x370;
  assign n4398 = n4397 ^ n4396;
  assign n4399 = ~x371 & ~x372;
  assign n4400 = ~x369 & ~x370;
  assign n4401 = ~n4399 & ~n4400;
  assign n4402 = n4401 ^ n4396;
  assign n4403 = n4402 ^ n4396;
  assign n4404 = n4396 ^ x368;
  assign n4405 = n4404 ^ n4396;
  assign n4406 = n4403 & n4405;
  assign n4407 = n4406 ^ n4396;
  assign n4408 = n4398 & ~n4407;
  assign n4409 = n4408 ^ n4397;
  assign n4410 = n4400 ^ n4399;
  assign n4411 = ~n4396 & ~n4397;
  assign n4412 = n4411 ^ n4400;
  assign n4413 = n4412 ^ n4400;
  assign n4414 = n4400 ^ x368;
  assign n4415 = n4414 ^ n4400;
  assign n4416 = n4413 & ~n4415;
  assign n4417 = n4416 ^ n4400;
  assign n4418 = n4410 & ~n4417;
  assign n4419 = n4418 ^ n4399;
  assign n4420 = ~n4409 & ~n4419;
  assign n4421 = ~x367 & ~n4420;
  assign n4422 = n4401 & ~n4411;
  assign n4423 = n2851 & n4422;
  assign n4424 = ~n4401 & n4411;
  assign n4425 = x367 & x368;
  assign n4426 = n4396 & n4425;
  assign n4427 = x372 & n4426;
  assign n4428 = n4427 ^ n4425;
  assign n4429 = ~n4424 & n4428;
  assign n4430 = ~n4423 & ~n4429;
  assign n4431 = n4425 ^ x370;
  assign n4432 = n4431 ^ n4425;
  assign n4433 = ~x368 & ~x372;
  assign n4434 = n4433 ^ n4425;
  assign n4435 = ~n4432 & n4434;
  assign n4436 = n4435 ^ n4425;
  assign n4437 = ~n2850 & n4436;
  assign n4438 = ~x371 & n4437;
  assign n4439 = n4430 & ~n4438;
  assign n4440 = ~n4421 & n4439;
  assign n4352 = x377 & x378;
  assign n4351 = x375 & x376;
  assign n4353 = n4352 ^ n4351;
  assign n4354 = ~x377 & ~x378;
  assign n4355 = ~x375 & ~x376;
  assign n4356 = ~n4354 & ~n4355;
  assign n4357 = n4356 ^ n4351;
  assign n4358 = n4357 ^ n4351;
  assign n4359 = n4351 ^ x374;
  assign n4360 = n4359 ^ n4351;
  assign n4361 = n4358 & n4360;
  assign n4362 = n4361 ^ n4351;
  assign n4363 = n4353 & ~n4362;
  assign n4364 = n4363 ^ n4352;
  assign n4365 = n4355 ^ n4354;
  assign n4366 = ~n4351 & ~n4352;
  assign n4367 = n4366 ^ n4355;
  assign n4368 = n4367 ^ n4355;
  assign n4369 = n4355 ^ x374;
  assign n4370 = n4369 ^ n4355;
  assign n4371 = n4368 & ~n4370;
  assign n4372 = n4371 ^ n4355;
  assign n4373 = n4365 & ~n4372;
  assign n4374 = n4373 ^ n4354;
  assign n4375 = ~n4364 & ~n4374;
  assign n4376 = ~x373 & ~n4375;
  assign n4377 = n4356 & ~n4366;
  assign n4378 = n2846 & n4377;
  assign n4379 = ~n4356 & n4366;
  assign n4380 = x373 & x374;
  assign n4381 = n4351 & n4380;
  assign n4382 = x378 & n4381;
  assign n4383 = n4382 ^ n4380;
  assign n4384 = ~n4379 & n4383;
  assign n4385 = ~n4378 & ~n4384;
  assign n4386 = n4380 ^ x376;
  assign n4387 = n4386 ^ n4380;
  assign n4388 = ~x374 & ~x378;
  assign n4389 = n4388 ^ n4380;
  assign n4390 = ~n4387 & n4389;
  assign n4391 = n4390 ^ n4380;
  assign n4392 = ~n2845 & n4391;
  assign n4393 = ~x377 & n4392;
  assign n4394 = n4385 & ~n4393;
  assign n4395 = ~n4376 & n4394;
  assign n4441 = n4440 ^ n4395;
  assign n4523 = n4522 ^ n4441;
  assign n6203 = ~n4441 & ~n4443;
  assign n6204 = n4523 & ~n6203;
  assign n6205 = ~n4521 & ~n6204;
  assign n6206 = ~n4441 & ~n4522;
  assign n6207 = n4444 & n4521;
  assign n6208 = n4441 & n4443;
  assign n6209 = ~n6207 & ~n6208;
  assign n6210 = ~n6206 & n6209;
  assign n6211 = ~n6205 & n6210;
  assign n6202 = ~n4364 & n4385;
  assign n6212 = n6211 ^ n6202;
  assign n6189 = n4443 ^ n4440;
  assign n6190 = ~n4441 & n6189;
  assign n6191 = n6190 ^ n4443;
  assign n7117 = n6202 ^ n6191;
  assign n7118 = ~n6212 & n7117;
  assign n7119 = n7118 ^ n6211;
  assign n6198 = ~n4489 & n4510;
  assign n6197 = ~n4455 & ~n4473;
  assign n6199 = n6198 ^ n6197;
  assign n6194 = n4475 ^ n4444;
  assign n6195 = n4521 & ~n6194;
  assign n6196 = n6195 ^ n4520;
  assign n6200 = n6199 ^ n6196;
  assign n6192 = ~n4409 & n4430;
  assign n7121 = n6200 ^ n6192;
  assign n6193 = n6192 ^ n6191;
  assign n6201 = n6200 ^ n6193;
  assign n6213 = n6212 ^ n6201;
  assign n7122 = n6213 ^ n6200;
  assign n7123 = ~n7121 & ~n7122;
  assign n7124 = n7123 ^ n6200;
  assign n7125 = ~n7119 & ~n7124;
  assign n7112 = n6198 ^ n6196;
  assign n7113 = ~n6199 & ~n7112;
  assign n7114 = n7113 ^ n6196;
  assign n7115 = n6192 & ~n6200;
  assign n7116 = ~n6213 & ~n7115;
  assign n7120 = n7116 & n7119;
  assign n7435 = ~n7114 & ~n7120;
  assign n7436 = ~n7125 & ~n7435;
  assign n7444 = n7443 ^ n7436;
  assign n2867 = n2866 ^ n2855;
  assign n2890 = n2889 ^ n2878;
  assign n4188 = n2867 & n2890;
  assign n4350 = n4349 ^ n4188;
  assign n6186 = n4523 ^ n4349;
  assign n6187 = ~n4350 & ~n6186;
  assign n6188 = n6187 ^ n4523;
  assign n6214 = n6213 ^ n6188;
  assign n7084 = n6188 ^ n6185;
  assign n7085 = ~n6214 & ~n7084;
  assign n7086 = n7085 ^ n6213;
  assign n7111 = n7110 ^ n7086;
  assign n7126 = ~n7120 & ~n7125;
  assign n7127 = n7126 ^ n7114;
  assign n7432 = n7127 ^ n7086;
  assign n7433 = n7111 & n7432;
  assign n7434 = n7433 ^ n7127;
  assign n7445 = n7444 ^ n7434;
  assign n2838 = x452 ^ x451;
  assign n2837 = x454 ^ x453;
  assign n4019 = x455 & x456;
  assign n4020 = n4019 ^ x454;
  assign n4021 = n2837 & ~n4020;
  assign n4022 = n4021 ^ x453;
  assign n4023 = n2838 & n4022;
  assign n4024 = ~x453 & ~x454;
  assign n4025 = ~n4019 & n4024;
  assign n4026 = x453 & x454;
  assign n4027 = x451 & x452;
  assign n4028 = ~n4026 & n4027;
  assign n4029 = ~n4025 & n4028;
  assign n4030 = ~n4023 & ~n4029;
  assign n4031 = ~x455 & ~x456;
  assign n4032 = ~n4030 & ~n4031;
  assign n4033 = n4026 & n4027;
  assign n4034 = ~x456 & n4033;
  assign n4035 = ~n4032 & ~n4034;
  assign n4036 = x452 & ~n4031;
  assign n4037 = n4019 & n4026;
  assign n4038 = ~n4036 & ~n4037;
  assign n4039 = n4022 & ~n4038;
  assign n4040 = n4031 ^ n4025;
  assign n4041 = n4031 ^ n4026;
  assign n4042 = n4025 ^ x452;
  assign n4043 = n4042 ^ n4031;
  assign n4044 = n4031 & ~n4043;
  assign n4045 = n4044 ^ n4031;
  assign n4046 = n4041 & n4045;
  assign n4047 = n4046 ^ n4044;
  assign n4048 = n4047 ^ n4031;
  assign n4049 = n4048 ^ n4042;
  assign n4050 = n4040 & ~n4049;
  assign n4051 = n4050 ^ n4025;
  assign n4052 = ~n4039 & ~n4051;
  assign n4053 = ~x451 & ~n4052;
  assign n4054 = ~x452 & ~x456;
  assign n4055 = n4024 & n4054;
  assign n4056 = ~n4033 & ~n4055;
  assign n4057 = ~x455 & ~n4056;
  assign n4058 = ~n4053 & ~n4057;
  assign n4059 = n4035 & n4058;
  assign n2833 = x458 ^ x457;
  assign n2832 = x460 ^ x459;
  assign n3978 = x461 & x462;
  assign n3979 = n3978 ^ x460;
  assign n3980 = n2832 & ~n3979;
  assign n3981 = n3980 ^ x459;
  assign n3982 = n2833 & n3981;
  assign n3983 = ~x459 & ~x460;
  assign n3984 = ~n3978 & n3983;
  assign n3985 = x459 & x460;
  assign n3986 = x457 & x458;
  assign n3987 = ~n3985 & n3986;
  assign n3988 = ~n3984 & n3987;
  assign n3989 = ~n3982 & ~n3988;
  assign n3990 = ~x461 & ~x462;
  assign n3991 = ~n3989 & ~n3990;
  assign n3992 = n3985 & n3986;
  assign n3993 = ~x462 & n3992;
  assign n3994 = ~n3991 & ~n3993;
  assign n3995 = x458 & ~n3990;
  assign n3996 = n3978 & n3985;
  assign n3997 = ~n3995 & ~n3996;
  assign n3998 = n3981 & ~n3997;
  assign n3999 = n3990 ^ n3984;
  assign n4000 = n3990 ^ n3985;
  assign n4001 = n3984 ^ x458;
  assign n4002 = n4001 ^ n3990;
  assign n4003 = n3990 & ~n4002;
  assign n4004 = n4003 ^ n3990;
  assign n4005 = n4000 & n4004;
  assign n4006 = n4005 ^ n4003;
  assign n4007 = n4006 ^ n3990;
  assign n4008 = n4007 ^ n4001;
  assign n4009 = n3999 & ~n4008;
  assign n4010 = n4009 ^ n3984;
  assign n4011 = ~n3998 & ~n4010;
  assign n4012 = ~x457 & ~n4011;
  assign n4013 = ~x458 & ~x462;
  assign n4014 = n3983 & n4013;
  assign n4015 = ~n3992 & ~n4014;
  assign n4016 = ~x461 & ~n4015;
  assign n4017 = ~n4012 & ~n4016;
  assign n4018 = n3994 & n4017;
  assign n4060 = n4059 ^ n4018;
  assign n2834 = x462 ^ x461;
  assign n2835 = n2834 ^ n2833;
  assign n2836 = n2835 ^ n2832;
  assign n2839 = x456 ^ x455;
  assign n2840 = n2839 ^ n2838;
  assign n2841 = n2840 ^ n2837;
  assign n4063 = n2836 & n2841;
  assign n6110 = n4063 ^ n4059;
  assign n6111 = ~n4060 & n6110;
  assign n6112 = n6111 ^ n4063;
  assign n4127 = x447 & x448;
  assign n4125 = ~x449 & ~x450;
  assign n4126 = x446 & ~n4125;
  assign n4128 = n4127 ^ n4126;
  assign n4129 = ~x447 & ~x448;
  assign n4130 = x449 & x450;
  assign n4131 = ~n4129 & n4130;
  assign n4132 = n4131 ^ n4126;
  assign n4133 = n4132 ^ n4131;
  assign n4134 = n4131 ^ n4130;
  assign n4135 = ~n4133 & ~n4134;
  assign n4136 = n4135 ^ n4131;
  assign n4137 = n4128 & n4136;
  assign n4138 = n4137 ^ n4127;
  assign n4139 = n4129 & ~n4130;
  assign n4140 = n4139 ^ n4125;
  assign n4141 = n4139 ^ n4127;
  assign n4142 = n4125 ^ x446;
  assign n4143 = n4142 ^ n4139;
  assign n4144 = ~n4139 & ~n4143;
  assign n4145 = n4144 ^ n4139;
  assign n4146 = ~n4141 & ~n4145;
  assign n4147 = n4146 ^ n4144;
  assign n4148 = n4147 ^ n4139;
  assign n4149 = n4148 ^ n4142;
  assign n4150 = n4140 & ~n4149;
  assign n4151 = n4150 ^ n4139;
  assign n4152 = ~n4138 & ~n4151;
  assign n4153 = ~x445 & ~n4152;
  assign n4154 = ~n4127 & ~n4131;
  assign n4155 = x445 & ~n4125;
  assign n4156 = ~n4154 & n4155;
  assign n4157 = x445 & x446;
  assign n4158 = ~n4156 & ~n4157;
  assign n4159 = n4127 ^ x450;
  assign n4161 = n4159 ^ n4129;
  assign n4160 = n4159 ^ x449;
  assign n4162 = n4161 ^ n4160;
  assign n4163 = n4159 ^ n4127;
  assign n4164 = n4163 ^ n4159;
  assign n4165 = n4164 ^ n4161;
  assign n4166 = ~n4161 & n4165;
  assign n4167 = n4166 ^ n4161;
  assign n4168 = ~n4162 & ~n4167;
  assign n4169 = n4168 ^ n4166;
  assign n4170 = n4169 ^ n4159;
  assign n4171 = n4170 ^ n4161;
  assign n4172 = x446 & n4171;
  assign n4173 = ~n4158 & ~n4172;
  assign n4174 = ~n4153 & ~n4173;
  assign n2828 = x448 ^ x447;
  assign n4175 = n4157 ^ x448;
  assign n4176 = n4175 ^ n4157;
  assign n4177 = ~x446 & ~x450;
  assign n4178 = n4177 ^ n4157;
  assign n4179 = ~n4176 & n4178;
  assign n4180 = n4179 ^ n4157;
  assign n4181 = ~n2828 & n4180;
  assign n4182 = ~x449 & n4181;
  assign n4183 = n4174 & ~n4182;
  assign n4068 = x441 & x442;
  assign n4066 = ~x443 & ~x444;
  assign n4067 = x440 & ~n4066;
  assign n4069 = n4068 ^ n4067;
  assign n4070 = ~x441 & ~x442;
  assign n4071 = x443 & x444;
  assign n4072 = ~n4070 & n4071;
  assign n4073 = n4072 ^ n4067;
  assign n4074 = n4073 ^ n4072;
  assign n4075 = n4072 ^ n4071;
  assign n4076 = ~n4074 & ~n4075;
  assign n4077 = n4076 ^ n4072;
  assign n4078 = n4069 & n4077;
  assign n4079 = n4078 ^ n4068;
  assign n4080 = n4070 & ~n4071;
  assign n4081 = n4080 ^ n4066;
  assign n4082 = n4080 ^ n4068;
  assign n4083 = n4066 ^ x440;
  assign n4084 = n4083 ^ n4080;
  assign n4085 = ~n4080 & ~n4084;
  assign n4086 = n4085 ^ n4080;
  assign n4087 = ~n4082 & ~n4086;
  assign n4088 = n4087 ^ n4085;
  assign n4089 = n4088 ^ n4080;
  assign n4090 = n4089 ^ n4083;
  assign n4091 = n4081 & ~n4090;
  assign n4092 = n4091 ^ n4080;
  assign n4093 = ~n4079 & ~n4092;
  assign n4094 = ~x439 & ~n4093;
  assign n4095 = ~n4068 & ~n4072;
  assign n4096 = x439 & ~n4066;
  assign n4097 = ~n4095 & n4096;
  assign n4098 = x439 & x440;
  assign n4099 = ~n4097 & ~n4098;
  assign n4100 = n4068 ^ x444;
  assign n4102 = n4100 ^ n4070;
  assign n4101 = n4100 ^ x443;
  assign n4103 = n4102 ^ n4101;
  assign n4104 = n4100 ^ n4068;
  assign n4105 = n4104 ^ n4100;
  assign n4106 = n4105 ^ n4102;
  assign n4107 = ~n4102 & n4106;
  assign n4108 = n4107 ^ n4102;
  assign n4109 = ~n4103 & ~n4108;
  assign n4110 = n4109 ^ n4107;
  assign n4111 = n4110 ^ n4100;
  assign n4112 = n4111 ^ n4102;
  assign n4113 = x440 & n4112;
  assign n4114 = ~n4099 & ~n4113;
  assign n4115 = ~n4094 & ~n4114;
  assign n2823 = x442 ^ x441;
  assign n4116 = n4098 ^ x442;
  assign n4117 = n4116 ^ n4098;
  assign n4118 = ~x440 & ~x444;
  assign n4119 = n4118 ^ n4098;
  assign n4120 = ~n4117 & n4119;
  assign n4121 = n4120 ^ n4098;
  assign n4122 = ~n2823 & n4121;
  assign n4123 = ~x443 & n4122;
  assign n4124 = n4115 & ~n4123;
  assign n4184 = n4183 ^ n4124;
  assign n2827 = x450 ^ x449;
  assign n2829 = n2828 ^ n2827;
  assign n2826 = x446 ^ x445;
  assign n2830 = n2829 ^ n2826;
  assign n2822 = x444 ^ x443;
  assign n2824 = n2823 ^ n2822;
  assign n2821 = x440 ^ x439;
  assign n2825 = n2824 ^ n2821;
  assign n2831 = n2830 ^ n2825;
  assign n2842 = n2841 ^ n2836;
  assign n4061 = n2831 & n2842;
  assign n4062 = n2825 & n2830;
  assign n4064 = n4063 ^ n4062;
  assign n4065 = ~n4061 & ~n4064;
  assign n4185 = n4184 ^ n4065;
  assign n4186 = n4185 ^ n4060;
  assign n6124 = n4060 & ~n4063;
  assign n6125 = ~n4186 & ~n6124;
  assign n6126 = n4184 ^ n4062;
  assign n6127 = ~n4061 & ~n6126;
  assign n6128 = ~n6125 & ~n6127;
  assign n6123 = n3994 & ~n3998;
  assign n6129 = n6128 ^ n6123;
  assign n6119 = ~n4079 & ~n4114;
  assign n6118 = ~n4138 & ~n4173;
  assign n6120 = n6119 ^ n6118;
  assign n6115 = n4124 ^ n4062;
  assign n6116 = n4184 & ~n6115;
  assign n6117 = n6116 ^ n4183;
  assign n6121 = n6120 ^ n6117;
  assign n6113 = n4035 & ~n4039;
  assign n6114 = n6113 ^ n6112;
  assign n6122 = n6121 ^ n6114;
  assign n6130 = n6129 ^ n6122;
  assign n7051 = ~n6112 & n6130;
  assign n7052 = n6123 ^ n6113;
  assign n7053 = ~n6129 & ~n7052;
  assign n7054 = n7053 ^ n6128;
  assign n7055 = n7051 & ~n7054;
  assign n7056 = n6123 & ~n6128;
  assign n7057 = n6113 & ~n6121;
  assign n7058 = n7056 & n7057;
  assign n7059 = ~n7055 & ~n7058;
  assign n7048 = n6119 ^ n6117;
  assign n7049 = ~n6120 & ~n7048;
  assign n7050 = n7049 ^ n6117;
  assign n7060 = n6121 & n7054;
  assign n7061 = ~n6130 & n7060;
  assign n7428 = ~n7050 & ~n7061;
  assign n7429 = n7059 & ~n7428;
  assign n2800 = x434 ^ x433;
  assign n2799 = x436 ^ x435;
  assign n2801 = n2800 ^ n2799;
  assign n2798 = x438 ^ x437;
  assign n2802 = n2801 ^ n2798;
  assign n2805 = x428 ^ x427;
  assign n2804 = x430 ^ x429;
  assign n2806 = n2805 ^ n2804;
  assign n2803 = x432 ^ x431;
  assign n2807 = n2806 ^ n2803;
  assign n3837 = n2802 & n2807;
  assign n3937 = x431 & x432;
  assign n3938 = x429 & x430;
  assign n3939 = ~n3937 & ~n3938;
  assign n3940 = ~x431 & ~x432;
  assign n3941 = ~x429 & ~x430;
  assign n3942 = ~n3940 & ~n3941;
  assign n3943 = n3939 & ~n3942;
  assign n3944 = x427 & x428;
  assign n3945 = n3938 & n3944;
  assign n3946 = x432 & n3945;
  assign n3947 = n3946 ^ n3944;
  assign n3948 = ~n3943 & n3947;
  assign n3949 = n3937 & n3938;
  assign n3950 = ~n3948 & ~n3949;
  assign n3951 = ~n3939 & n3942;
  assign n3952 = ~x428 & n3951;
  assign n3953 = ~x427 & n3952;
  assign n3954 = n3953 ^ n3951;
  assign n3955 = n3950 & ~n3954;
  assign n3956 = x431 ^ x428;
  assign n3957 = n2803 & n3956;
  assign n3958 = n3957 ^ x431;
  assign n3959 = n3941 & ~n3958;
  assign n3960 = n3955 & ~n3959;
  assign n3961 = x427 & ~n3948;
  assign n3962 = ~n3952 & n3961;
  assign n3963 = ~n3960 & ~n3962;
  assign n3964 = ~x428 & ~x432;
  assign n3965 = n3964 ^ n3944;
  assign n3966 = n3965 ^ n3944;
  assign n3967 = n3944 ^ n2806;
  assign n3968 = n3967 ^ n3944;
  assign n3969 = n3966 & n3968;
  assign n3970 = n3969 ^ n3944;
  assign n3971 = ~n3938 & n3970;
  assign n3972 = n3971 ^ n3944;
  assign n3973 = ~x431 & n3972;
  assign n3974 = ~n3963 & ~n3973;
  assign n3900 = x437 & x438;
  assign n3901 = x435 & x436;
  assign n3902 = n3900 & n3901;
  assign n3903 = ~n3900 & ~n3901;
  assign n3904 = ~x437 & ~x438;
  assign n3905 = ~x435 & ~x436;
  assign n3906 = ~n3904 & ~n3905;
  assign n3907 = ~n3903 & n3906;
  assign n3908 = ~x434 & n3907;
  assign n3909 = ~x433 & n3908;
  assign n3910 = n3909 ^ n3907;
  assign n3911 = ~n3902 & ~n3910;
  assign n3912 = x437 ^ x434;
  assign n3913 = n2798 & n3912;
  assign n3914 = n3913 ^ x437;
  assign n3915 = n3905 & ~n3914;
  assign n3916 = n3911 & ~n3915;
  assign n3917 = x433 & ~n3908;
  assign n3918 = ~n3916 & ~n3917;
  assign n3919 = x433 & x434;
  assign n3920 = n3919 ^ n2801;
  assign n3921 = n3920 ^ n3919;
  assign n3922 = ~x434 & ~x438;
  assign n3923 = n3922 ^ n3919;
  assign n3924 = n3923 ^ n3919;
  assign n3925 = n3921 & n3924;
  assign n3926 = n3925 ^ n3919;
  assign n3927 = ~n3901 & n3926;
  assign n3928 = n3927 ^ n3919;
  assign n3929 = ~x437 & n3928;
  assign n3930 = n3903 & ~n3906;
  assign n3931 = n3901 & n3919;
  assign n3932 = x438 & n3931;
  assign n3933 = n3932 ^ n3919;
  assign n3934 = ~n3930 & n3933;
  assign n3935 = ~n3929 & ~n3934;
  assign n3936 = ~n3918 & n3935;
  assign n3975 = n3974 ^ n3936;
  assign n6145 = ~n3837 & n3975;
  assign n6146 = ~n3936 & ~n3974;
  assign n6147 = ~n6145 & ~n6146;
  assign n3871 = x419 & x420;
  assign n3872 = ~x417 & ~x418;
  assign n3873 = ~n3871 & n3872;
  assign n3874 = ~x419 & ~x420;
  assign n3875 = x416 & ~n3874;
  assign n3876 = n3873 & ~n3875;
  assign n3877 = x417 & x418;
  assign n3878 = n3871 & n3877;
  assign n3879 = ~n3876 & ~n3878;
  assign n3880 = ~x415 & ~n3879;
  assign n2811 = x416 ^ x415;
  assign n2810 = x418 ^ x417;
  assign n2812 = n2811 ^ n2810;
  assign n3881 = ~x416 & n3874;
  assign n3882 = ~n3877 & n3881;
  assign n3883 = n2812 & n3882;
  assign n3884 = x415 & x416;
  assign n3885 = n3877 & n3884;
  assign n3886 = ~n3871 & n3885;
  assign n3887 = ~n3883 & ~n3886;
  assign n3888 = ~n3880 & n3887;
  assign n3889 = ~n3877 & n3884;
  assign n3890 = ~n3873 & n3889;
  assign n3891 = n3871 ^ x418;
  assign n3892 = n2810 & n3891;
  assign n3893 = n3892 ^ x418;
  assign n3894 = n2811 & n3893;
  assign n3895 = ~n3890 & ~n3894;
  assign n3896 = ~n3874 & ~n3895;
  assign n3897 = n3888 & ~n3896;
  assign n3841 = x423 & x424;
  assign n3842 = x425 & x426;
  assign n3843 = n3841 & n3842;
  assign n3844 = ~x423 & ~x424;
  assign n3845 = ~n3842 & n3844;
  assign n3846 = n3845 ^ x422;
  assign n3847 = ~x425 & ~x426;
  assign n3848 = n3847 ^ n3845;
  assign n3849 = n3848 ^ n3847;
  assign n3850 = ~n3841 & n3847;
  assign n3851 = n3850 ^ n3847;
  assign n3852 = ~n3849 & ~n3851;
  assign n3853 = n3852 ^ n3847;
  assign n3854 = ~n3846 & n3853;
  assign n3855 = n3854 ^ x422;
  assign n3856 = ~n3843 & n3855;
  assign n3857 = ~x421 & ~n3856;
  assign n2816 = x422 ^ x421;
  assign n3858 = n3842 & ~n3844;
  assign n3859 = n3841 & ~n3847;
  assign n3860 = ~n3858 & ~n3859;
  assign n3861 = n2816 & ~n3860;
  assign n3862 = x421 & x422;
  assign n3863 = ~n3845 & n3862;
  assign n3864 = ~n3843 & ~n3850;
  assign n3865 = n3863 & n3864;
  assign n3866 = ~n3861 & ~n3865;
  assign n3867 = ~x422 & n3850;
  assign n3868 = n3844 & n3867;
  assign n3869 = n3866 & ~n3868;
  assign n3870 = ~n3857 & n3869;
  assign n3898 = n3897 ^ n3870;
  assign n2809 = x420 ^ x419;
  assign n2813 = n2812 ^ n2809;
  assign n2815 = x426 ^ x425;
  assign n2817 = n2816 ^ n2815;
  assign n2814 = x424 ^ x423;
  assign n2818 = n2817 ^ n2814;
  assign n3833 = n2813 & n2818;
  assign n2808 = n2807 ^ n2802;
  assign n2819 = n2818 ^ n2813;
  assign n3834 = n2819 ^ n2807;
  assign n3835 = ~n2808 & n3834;
  assign n3836 = n3835 ^ n2819;
  assign n3838 = n3837 ^ n3836;
  assign n3839 = ~n3833 & ~n3838;
  assign n3840 = n3839 ^ n3837;
  assign n3899 = n3898 ^ n3840;
  assign n3976 = n3975 ^ n3899;
  assign n6148 = ~n3833 & n3898;
  assign n6149 = ~n3976 & ~n6148;
  assign n6150 = ~n3838 & ~n3975;
  assign n6151 = n6150 ^ n3837;
  assign n6152 = ~n6149 & ~n6151;
  assign n7071 = n6147 & n6152;
  assign n6134 = n3911 & ~n3934;
  assign n7072 = ~n3955 & ~n6134;
  assign n7073 = ~n7071 & ~n7072;
  assign n6141 = ~n3843 & n3866;
  assign n6139 = ~n3878 & ~n3885;
  assign n6140 = ~n3896 & n6139;
  assign n6142 = n6141 ^ n6140;
  assign n6136 = n3897 ^ n3833;
  assign n6137 = ~n3898 & n6136;
  assign n6138 = n6137 ^ n3833;
  assign n6143 = n6142 ^ n6138;
  assign n6135 = n6134 ^ n3955;
  assign n6144 = n6143 ^ n6135;
  assign n6153 = n6152 ^ n6147;
  assign n7075 = n6153 ^ n6143;
  assign n7076 = n6144 & n7075;
  assign n7077 = n7076 ^ n6143;
  assign n7078 = n7073 & ~n7077;
  assign n7067 = n6141 ^ n6138;
  assign n7068 = ~n6142 & ~n7067;
  assign n7069 = n7068 ^ n6138;
  assign n6154 = n6153 ^ n6144;
  assign n7070 = n6143 & ~n6154;
  assign n7074 = n7070 & ~n7073;
  assign n7426 = ~n7069 & ~n7074;
  assign n7427 = ~n7078 & ~n7426;
  assign n7430 = n7429 ^ n7427;
  assign n7079 = ~n7074 & ~n7078;
  assign n7080 = n7079 ^ n7069;
  assign n2820 = n2819 ^ n2808;
  assign n2843 = n2842 ^ n2831;
  assign n3832 = n2820 & n2843;
  assign n3977 = n3976 ^ n3832;
  assign n6131 = n4186 ^ n3832;
  assign n6132 = ~n3977 & n6131;
  assign n6133 = n6132 ^ n3976;
  assign n6155 = n6154 ^ n6133;
  assign n7064 = n6133 ^ n6130;
  assign n7065 = ~n6155 & n7064;
  assign n7066 = n7065 ^ n6154;
  assign n7081 = n7080 ^ n7066;
  assign n7062 = n7059 & ~n7061;
  assign n7063 = n7062 ^ n7050;
  assign n7423 = n7066 ^ n7063;
  assign n7424 = n7081 & ~n7423;
  assign n7425 = n7424 ^ n7080;
  assign n7431 = n7430 ^ n7425;
  assign n7446 = n7445 ^ n7431;
  assign n7082 = n7081 ^ n7063;
  assign n6156 = n6155 ^ n6130;
  assign n4524 = n4523 ^ n4350;
  assign n2844 = n2843 ^ n2820;
  assign n2891 = n2890 ^ n2867;
  assign n3829 = n2844 & n2891;
  assign n6106 = n4524 ^ n3829;
  assign n4187 = n4186 ^ n3977;
  assign n6107 = n4187 ^ n3829;
  assign n6108 = ~n6106 & ~n6107;
  assign n6109 = n6108 ^ n4524;
  assign n6157 = n6156 ^ n6109;
  assign n6215 = n6214 ^ n6185;
  assign n7045 = n6215 ^ n6156;
  assign n7046 = ~n6157 & ~n7045;
  assign n7047 = n7046 ^ n6215;
  assign n7083 = n7082 ^ n7047;
  assign n7128 = n7127 ^ n7111;
  assign n7420 = n7128 ^ n7047;
  assign n7421 = n7083 & n7420;
  assign n7422 = n7421 ^ n7082;
  assign n7613 = n7431 ^ n7422;
  assign n7614 = n7446 & ~n7613;
  assign n7615 = n7614 ^ n7445;
  assign n7616 = n7429 ^ n7425;
  assign n7617 = ~n7430 & n7616;
  assign n7618 = n7617 ^ n7425;
  assign n7619 = n7443 ^ n7434;
  assign n7620 = ~n7444 & n7619;
  assign n7621 = n7620 ^ n7434;
  assign n7712 = n7618 & n7621;
  assign n7713 = n7615 & n7712;
  assign n7718 = n7717 ^ n7713;
  assign n7719 = ~n7673 & ~n7718;
  assign n7447 = n7446 ^ n7422;
  assign n7129 = n7128 ^ n7083;
  assign n6216 = n6215 ^ n6157;
  assign n2892 = n2891 ^ n2844;
  assign n2987 = n2986 ^ n2939;
  assign n3830 = n2892 & n2987;
  assign n3186 = ~n3184 & ~n3185;
  assign n3500 = n3499 ^ n3186;
  assign n3828 = n3827 ^ n3500;
  assign n6097 = n3830 ^ n3828;
  assign n4525 = n4524 ^ n4187;
  assign n6098 = n4525 ^ n3829;
  assign n6099 = n6098 ^ n4525;
  assign n6100 = n4525 ^ n3828;
  assign n6101 = n6100 ^ n4525;
  assign n6102 = ~n6099 & ~n6101;
  assign n6103 = n6102 ^ n4525;
  assign n6104 = ~n6097 & n6103;
  assign n6105 = n6104 ^ n3830;
  assign n6217 = n6216 ^ n6105;
  assign n6337 = n6336 ^ n6274;
  assign n7042 = n6337 ^ n6105;
  assign n7043 = n6217 & n7042;
  assign n7044 = n7043 ^ n6216;
  assign n7130 = n7129 ^ n7044;
  assign n7210 = n7209 ^ n7161;
  assign n7417 = n7210 ^ n7044;
  assign n7418 = ~n7130 & n7417;
  assign n7419 = n7418 ^ n7129;
  assign n7448 = n7447 ^ n7419;
  assign n7485 = ~n7483 & ~n7484;
  assign n7497 = n7496 ^ n7485;
  assign n7624 = n7497 ^ n7447;
  assign n7625 = n7448 & n7624;
  assign n7626 = n7625 ^ n7497;
  assign n7723 = ~n7618 & ~n7621;
  assign n7724 = ~n7615 & n7723;
  assign n7622 = n7621 ^ n7618;
  assign n7720 = n7621 ^ n7615;
  assign n7721 = ~n7622 & n7720;
  assign n7722 = n7721 ^ n7615;
  assign n7725 = n7724 ^ n7722;
  assign n7726 = n7626 & n7725;
  assign n7727 = n7726 ^ n7724;
  assign n7728 = n7719 & ~n7727;
  assign n7747 = ~n7717 & n7728;
  assign n7731 = ~n7626 & ~n7722;
  assign n7748 = n7716 & ~n7731;
  assign n7749 = n7673 & ~n7748;
  assign n7750 = ~n7724 & ~n7749;
  assign n7751 = ~n7747 & n7750;
  assign n7605 = n7340 & ~n7591;
  assign n7606 = n7605 ^ n7604;
  assign n7607 = n7566 & n7606;
  assign n7608 = n7607 ^ n7604;
  assign n7609 = n7590 & ~n7608;
  assign n5682 = x171 & x172;
  assign n5681 = x173 & x174;
  assign n5683 = n5682 ^ n5681;
  assign n5684 = ~x171 & ~x172;
  assign n5685 = ~x173 & ~x174;
  assign n5686 = ~n5684 & ~n5685;
  assign n5687 = n5686 ^ n5681;
  assign n5688 = n5687 ^ n5681;
  assign n5689 = n5681 ^ x170;
  assign n5690 = n5689 ^ n5681;
  assign n5691 = n5688 & n5690;
  assign n5692 = n5691 ^ n5681;
  assign n5693 = n5683 & ~n5692;
  assign n5694 = n5693 ^ n5682;
  assign n5696 = ~n5681 & ~n5682;
  assign n5709 = n5686 & ~n5696;
  assign n5708 = x174 & n5682;
  assign n5710 = n5709 ^ n5708;
  assign n5711 = n5710 ^ n5709;
  assign n5712 = ~n5686 & n5696;
  assign n5713 = n5712 ^ n5709;
  assign n5714 = n5713 ^ n5709;
  assign n5715 = ~n5711 & ~n5714;
  assign n5716 = n5715 ^ n5709;
  assign n5717 = x170 & n5716;
  assign n5718 = n5717 ^ n5709;
  assign n6476 = x169 & n5718;
  assign n6477 = ~n5694 & ~n6476;
  assign n5726 = x165 & x166;
  assign n5727 = x167 & x168;
  assign n5731 = n5726 & n5727;
  assign n5735 = x163 & x164;
  assign n5737 = ~n5731 & n5735;
  assign n5728 = ~n5726 & ~n5727;
  assign n5738 = n5737 ^ n5728;
  assign n3149 = x164 ^ x163;
  assign n5739 = n5737 ^ n3149;
  assign n5723 = ~x165 & ~x166;
  assign n5724 = ~x167 & ~x168;
  assign n5725 = ~n5723 & ~n5724;
  assign n5740 = n5728 ^ n5725;
  assign n5741 = n5740 ^ n5737;
  assign n5742 = ~n5737 & ~n5741;
  assign n5743 = n5742 ^ n5737;
  assign n5744 = n5739 & ~n5743;
  assign n5745 = n5744 ^ n5742;
  assign n5746 = n5745 ^ n5737;
  assign n5747 = n5746 ^ n5740;
  assign n5748 = ~n5738 & ~n5747;
  assign n5749 = n5748 ^ n5737;
  assign n6475 = ~n5731 & ~n5749;
  assign n6478 = n6477 ^ n6475;
  assign n5729 = ~n5725 & n5728;
  assign n5730 = ~n3149 & n5729;
  assign n5732 = n5723 & n5724;
  assign n5733 = ~n5731 & ~n5732;
  assign n5734 = ~n5730 & n5733;
  assign n5736 = ~n5734 & ~n5735;
  assign n5750 = ~n5736 & ~n5749;
  assign n3144 = x172 ^ x171;
  assign n5672 = x169 & x170;
  assign n5673 = n5672 ^ x172;
  assign n5674 = n5673 ^ n5672;
  assign n5675 = ~x170 & ~x174;
  assign n5676 = n5675 ^ n5672;
  assign n5677 = ~n5674 & n5676;
  assign n5678 = n5677 ^ n5672;
  assign n5679 = ~n3144 & n5678;
  assign n5680 = ~x173 & n5679;
  assign n5695 = n5685 ^ n5684;
  assign n5697 = n5696 ^ n5685;
  assign n5698 = n5697 ^ n5685;
  assign n5699 = n5685 ^ x170;
  assign n5700 = n5699 ^ n5685;
  assign n5701 = n5698 & ~n5700;
  assign n5702 = n5701 ^ n5685;
  assign n5703 = n5695 & ~n5702;
  assign n5704 = n5703 ^ n5684;
  assign n5705 = ~n5694 & ~n5704;
  assign n5706 = n5705 ^ x169;
  assign n5707 = n5706 ^ n5705;
  assign n5719 = n5718 ^ n5705;
  assign n5720 = n5707 & ~n5719;
  assign n5721 = n5720 ^ n5705;
  assign n5722 = ~n5680 & n5721;
  assign n5751 = n5750 ^ n5722;
  assign n3143 = x174 ^ x173;
  assign n3145 = n3144 ^ n3143;
  assign n3142 = x170 ^ x169;
  assign n3146 = n3145 ^ n3142;
  assign n3148 = x166 ^ x165;
  assign n3150 = n3149 ^ n3148;
  assign n3147 = x168 ^ x167;
  assign n3151 = n3150 ^ n3147;
  assign n5671 = n3146 & n3151;
  assign n6472 = n5750 ^ n5671;
  assign n6473 = n5751 & ~n6472;
  assign n6474 = n6473 ^ n5722;
  assign n7012 = n6477 ^ n6474;
  assign n7013 = ~n6478 & ~n7012;
  assign n7014 = n7013 ^ n6474;
  assign n5444 = x147 & x148;
  assign n5443 = x149 & x150;
  assign n5445 = n5444 ^ n5443;
  assign n5446 = ~x147 & ~x148;
  assign n5447 = ~x149 & ~x150;
  assign n5448 = ~n5446 & ~n5447;
  assign n5449 = n5448 ^ n5443;
  assign n5450 = n5449 ^ n5443;
  assign n5451 = n5443 ^ x146;
  assign n5452 = n5451 ^ n5443;
  assign n5453 = n5450 & n5452;
  assign n5454 = n5453 ^ n5443;
  assign n5455 = n5445 & ~n5454;
  assign n5456 = n5455 ^ n5444;
  assign n3172 = x146 ^ x145;
  assign n5458 = ~n5443 & ~n5444;
  assign n5469 = n5448 & ~n5458;
  assign n5470 = n3172 & n5469;
  assign n5471 = ~n5448 & n5458;
  assign n5472 = x145 & x146;
  assign n5473 = n5444 & n5472;
  assign n5474 = x150 & n5473;
  assign n5475 = n5474 ^ n5472;
  assign n5476 = ~n5471 & n5475;
  assign n5477 = ~n5470 & ~n5476;
  assign n6425 = ~n5456 & n5477;
  assign n5399 = x141 & x142;
  assign n5398 = x143 & x144;
  assign n5400 = n5399 ^ n5398;
  assign n5401 = ~x141 & ~x142;
  assign n5402 = ~x143 & ~x144;
  assign n5403 = ~n5401 & ~n5402;
  assign n5404 = n5403 ^ n5398;
  assign n5405 = n5404 ^ n5398;
  assign n5406 = n5398 ^ x140;
  assign n5407 = n5406 ^ n5398;
  assign n5408 = n5405 & n5407;
  assign n5409 = n5408 ^ n5398;
  assign n5410 = n5400 & ~n5409;
  assign n5411 = n5410 ^ n5399;
  assign n3167 = x140 ^ x139;
  assign n5413 = ~n5398 & ~n5399;
  assign n5424 = n5403 & ~n5413;
  assign n5425 = n3167 & n5424;
  assign n5426 = ~n5403 & n5413;
  assign n5427 = x139 & x140;
  assign n5428 = n5399 & n5427;
  assign n5429 = x144 & n5428;
  assign n5430 = n5429 ^ n5427;
  assign n5431 = ~n5426 & n5430;
  assign n5432 = ~n5425 & ~n5431;
  assign n6426 = ~n5411 & n5432;
  assign n7030 = ~n6425 & ~n6426;
  assign n3156 = x134 ^ x133;
  assign n3155 = x136 ^ x135;
  assign n5531 = x137 & x138;
  assign n5532 = n5531 ^ x136;
  assign n5533 = n3155 & ~n5532;
  assign n5534 = n5533 ^ x135;
  assign n5535 = n3156 & n5534;
  assign n5536 = ~x135 & ~x136;
  assign n5537 = ~n5531 & n5536;
  assign n5538 = x135 & x136;
  assign n5539 = x133 & x134;
  assign n5540 = ~n5538 & n5539;
  assign n5541 = ~n5537 & n5540;
  assign n5542 = ~n5535 & ~n5541;
  assign n5543 = ~x137 & ~x138;
  assign n5544 = ~n5542 & ~n5543;
  assign n5545 = n5538 & n5539;
  assign n5546 = ~x138 & n5545;
  assign n5547 = ~n5544 & ~n5546;
  assign n5548 = x134 & ~n5543;
  assign n5549 = n5531 & n5538;
  assign n5550 = ~n5548 & ~n5549;
  assign n5551 = n5534 & ~n5550;
  assign n6433 = n5547 & ~n5551;
  assign n3161 = x128 ^ x127;
  assign n3159 = x130 ^ x129;
  assign n5490 = x131 & x132;
  assign n5491 = n5490 ^ x130;
  assign n5492 = n3159 & ~n5491;
  assign n5493 = n5492 ^ x129;
  assign n5494 = n3161 & n5493;
  assign n5495 = ~x129 & ~x130;
  assign n5496 = ~n5490 & n5495;
  assign n5497 = x129 & x130;
  assign n5498 = x127 & x128;
  assign n5499 = ~n5497 & n5498;
  assign n5500 = ~n5496 & n5499;
  assign n5501 = ~n5494 & ~n5500;
  assign n5502 = ~x131 & ~x132;
  assign n5503 = ~n5501 & ~n5502;
  assign n5504 = n5497 & n5498;
  assign n5505 = ~x132 & n5504;
  assign n5506 = ~n5503 & ~n5505;
  assign n5507 = x128 & ~n5502;
  assign n5508 = n5490 & n5497;
  assign n5509 = ~n5507 & ~n5508;
  assign n5510 = n5493 & ~n5509;
  assign n6432 = n5506 & ~n5510;
  assign n6434 = n6433 ^ n6432;
  assign n5552 = n5537 & ~n5548;
  assign n5553 = ~n5551 & ~n5552;
  assign n5554 = ~x133 & ~n5553;
  assign n5555 = n5547 & ~n5554;
  assign n5556 = ~x134 & ~x138;
  assign n5557 = n5556 ^ n5539;
  assign n5558 = n5557 ^ n5539;
  assign n3157 = n3156 ^ n3155;
  assign n5559 = n5539 ^ n3157;
  assign n5560 = n5559 ^ n5539;
  assign n5561 = n5558 & n5560;
  assign n5562 = n5561 ^ n5539;
  assign n5563 = ~n5538 & n5562;
  assign n5564 = n5563 ^ n5539;
  assign n5565 = ~x137 & n5564;
  assign n5566 = n5555 & ~n5565;
  assign n5511 = n5502 ^ n5496;
  assign n5512 = n5502 ^ n5497;
  assign n5513 = n5496 ^ x128;
  assign n5514 = n5513 ^ n5502;
  assign n5515 = n5502 & ~n5514;
  assign n5516 = n5515 ^ n5502;
  assign n5517 = n5512 & n5516;
  assign n5518 = n5517 ^ n5515;
  assign n5519 = n5518 ^ n5502;
  assign n5520 = n5519 ^ n5513;
  assign n5521 = n5511 & ~n5520;
  assign n5522 = n5521 ^ n5496;
  assign n5523 = ~n5510 & ~n5522;
  assign n5524 = ~x127 & ~n5523;
  assign n5525 = ~x128 & ~x132;
  assign n5526 = n5495 & n5525;
  assign n5527 = ~n5504 & ~n5526;
  assign n5528 = ~x131 & ~n5527;
  assign n5529 = ~n5524 & ~n5528;
  assign n5530 = n5506 & n5529;
  assign n5567 = n5566 ^ n5530;
  assign n3154 = x138 ^ x137;
  assign n3158 = n3157 ^ n3154;
  assign n3160 = x132 ^ x131;
  assign n3162 = n3161 ^ n3160;
  assign n3163 = n3162 ^ n3159;
  assign n6428 = n3158 & n3163;
  assign n6429 = n6428 ^ n5530;
  assign n6430 = n5567 & ~n6429;
  assign n6431 = n6430 ^ n5566;
  assign n6435 = n6434 ^ n6431;
  assign n5457 = n5447 ^ n5446;
  assign n5459 = n5458 ^ n5447;
  assign n5460 = n5459 ^ n5447;
  assign n5461 = n5447 ^ x146;
  assign n5462 = n5461 ^ n5447;
  assign n5463 = n5460 & ~n5462;
  assign n5464 = n5463 ^ n5447;
  assign n5465 = n5457 & ~n5464;
  assign n5466 = n5465 ^ n5446;
  assign n5467 = ~n5456 & ~n5466;
  assign n5468 = ~x145 & ~n5467;
  assign n3171 = x148 ^ x147;
  assign n5478 = n5472 ^ x148;
  assign n5479 = n5478 ^ n5472;
  assign n5480 = ~x146 & ~x150;
  assign n5481 = n5480 ^ n5472;
  assign n5482 = ~n5479 & n5481;
  assign n5483 = n5482 ^ n5472;
  assign n5484 = ~n3171 & n5483;
  assign n5485 = ~x149 & n5484;
  assign n5486 = n5477 & ~n5485;
  assign n5487 = ~n5468 & n5486;
  assign n5412 = n5402 ^ n5401;
  assign n5414 = n5413 ^ n5402;
  assign n5415 = n5414 ^ n5402;
  assign n5416 = n5402 ^ x140;
  assign n5417 = n5416 ^ n5402;
  assign n5418 = n5415 & ~n5417;
  assign n5419 = n5418 ^ n5402;
  assign n5420 = n5412 & ~n5419;
  assign n5421 = n5420 ^ n5401;
  assign n5422 = ~n5411 & ~n5421;
  assign n5423 = ~x139 & ~n5422;
  assign n3166 = x142 ^ x141;
  assign n5433 = n5427 ^ x142;
  assign n5434 = n5433 ^ n5427;
  assign n5435 = ~x140 & ~x144;
  assign n5436 = n5435 ^ n5427;
  assign n5437 = ~n5434 & n5436;
  assign n5438 = n5437 ^ n5427;
  assign n5439 = ~n3166 & n5438;
  assign n5440 = ~x143 & n5439;
  assign n5441 = n5432 & ~n5440;
  assign n5442 = ~n5423 & n5441;
  assign n5488 = n5487 ^ n5442;
  assign n3168 = n3167 ^ n3166;
  assign n3165 = x144 ^ x143;
  assign n3169 = n3168 ^ n3165;
  assign n3173 = n3172 ^ n3171;
  assign n3170 = x150 ^ x149;
  assign n3174 = n3173 ^ n3170;
  assign n6437 = n3169 & n3174;
  assign n6438 = n6437 ^ n5442;
  assign n6439 = n5488 & ~n6438;
  assign n6440 = n6439 ^ n5487;
  assign n5393 = n3169 ^ n3163;
  assign n5395 = n5393 ^ n3158;
  assign n5396 = ~n3174 & n5395;
  assign n3164 = n3163 ^ n3158;
  assign n5394 = ~n3164 & ~n5393;
  assign n5397 = n5396 ^ n5394;
  assign n5489 = n5488 ^ n5397;
  assign n6441 = ~n5489 & ~n5567;
  assign n3175 = n3174 ^ n3169;
  assign n3176 = n3175 ^ n3164;
  assign n6442 = ~n3163 & ~n6437;
  assign n6443 = n3176 & n6442;
  assign n6444 = ~n3169 & ~n3174;
  assign n6445 = ~n6443 & ~n6444;
  assign n6446 = ~n5488 & ~n6445;
  assign n6447 = n5488 & n6437;
  assign n6448 = ~n6446 & ~n6447;
  assign n6449 = ~n6441 & n6448;
  assign n6450 = n5567 & n6428;
  assign n6451 = n6449 & ~n6450;
  assign n7024 = ~n6440 & ~n6451;
  assign n7025 = ~n6435 & n7024;
  assign n6427 = n6426 ^ n6425;
  assign n7026 = n6440 & n6451;
  assign n7027 = n6427 & ~n7026;
  assign n7028 = ~n7025 & n7027;
  assign n7029 = n6435 & ~n7024;
  assign n7032 = n6425 & n6426;
  assign n7031 = ~n7026 & ~n7030;
  assign n7033 = n7032 ^ n7031;
  assign n7034 = ~n7029 & ~n7033;
  assign n7035 = n7034 ^ n7032;
  assign n7036 = ~n7028 & ~n7035;
  assign n7021 = n6433 ^ n6431;
  assign n7022 = ~n6434 & ~n7021;
  assign n7023 = n7022 ^ n6431;
  assign n7037 = n7036 ^ n7023;
  assign n7377 = ~n7030 & ~n7037;
  assign n7378 = ~n7023 & ~n7029;
  assign n7379 = ~n7377 & ~n7378;
  assign n6479 = n6478 ^ n6474;
  assign n5574 = x159 & x160;
  assign n5572 = ~x161 & ~x162;
  assign n5573 = x158 & ~n5572;
  assign n5575 = n5574 ^ n5573;
  assign n5576 = ~x159 & ~x160;
  assign n5577 = x161 & x162;
  assign n5578 = ~n5576 & n5577;
  assign n5579 = n5578 ^ n5573;
  assign n5580 = n5579 ^ n5578;
  assign n5581 = n5578 ^ n5577;
  assign n5582 = ~n5580 & ~n5581;
  assign n5583 = n5582 ^ n5578;
  assign n5584 = n5575 & n5583;
  assign n5585 = n5584 ^ n5574;
  assign n5586 = n5576 & ~n5577;
  assign n5587 = n5586 ^ n5572;
  assign n5588 = n5586 ^ n5574;
  assign n5589 = n5572 ^ x158;
  assign n5590 = n5589 ^ n5586;
  assign n5591 = ~n5586 & ~n5590;
  assign n5592 = n5591 ^ n5586;
  assign n5593 = ~n5588 & ~n5592;
  assign n5594 = n5593 ^ n5591;
  assign n5595 = n5594 ^ n5586;
  assign n5596 = n5595 ^ n5589;
  assign n5597 = n5587 & ~n5596;
  assign n5598 = n5597 ^ n5586;
  assign n5599 = ~n5585 & ~n5598;
  assign n5600 = ~x157 & ~n5599;
  assign n5601 = ~n5574 & ~n5578;
  assign n5602 = x157 & ~n5572;
  assign n5603 = ~n5601 & n5602;
  assign n5604 = x157 & x158;
  assign n5605 = ~n5603 & ~n5604;
  assign n5606 = n5574 ^ x162;
  assign n5608 = n5606 ^ n5576;
  assign n5607 = n5606 ^ x161;
  assign n5609 = n5608 ^ n5607;
  assign n5610 = n5606 ^ n5574;
  assign n5611 = n5610 ^ n5606;
  assign n5612 = n5611 ^ n5608;
  assign n5613 = ~n5608 & n5612;
  assign n5614 = n5613 ^ n5608;
  assign n5615 = ~n5609 & ~n5614;
  assign n5616 = n5615 ^ n5613;
  assign n5617 = n5616 ^ n5606;
  assign n5618 = n5617 ^ n5608;
  assign n5619 = x158 & n5618;
  assign n5620 = ~n5605 & ~n5619;
  assign n5621 = ~n5600 & ~n5620;
  assign n3133 = x160 ^ x159;
  assign n5622 = n5604 ^ x160;
  assign n5623 = n5622 ^ n5604;
  assign n5624 = ~x158 & ~x162;
  assign n5625 = n5624 ^ n5604;
  assign n5626 = ~n5623 & n5625;
  assign n5627 = n5626 ^ n5604;
  assign n5628 = ~n3133 & n5627;
  assign n5629 = ~x161 & n5628;
  assign n5630 = n5621 & ~n5629;
  assign n5631 = ~x155 & ~x156;
  assign n5632 = x152 & ~n5631;
  assign n5633 = x155 & x156;
  assign n5634 = ~x153 & ~x154;
  assign n5635 = ~n5633 & n5634;
  assign n5636 = ~n5632 & n5635;
  assign n5637 = x153 & x154;
  assign n5638 = n5637 ^ n5633;
  assign n5639 = n5637 ^ n5632;
  assign n5640 = n5638 & n5639;
  assign n5641 = n5640 ^ n5637;
  assign n5642 = ~n5634 & n5641;
  assign n5643 = ~n5636 & ~n5642;
  assign n5644 = ~x151 & ~n5643;
  assign n5645 = ~n5633 & ~n5637;
  assign n5646 = ~n5634 & ~n5645;
  assign n5647 = x151 & ~n5631;
  assign n5648 = n5646 & n5647;
  assign n5649 = x151 & x152;
  assign n5650 = ~n5648 & ~n5649;
  assign n5651 = ~n5631 & ~n5637;
  assign n5652 = ~n5635 & n5651;
  assign n5653 = ~x156 & n5637;
  assign n5654 = x152 & ~n5653;
  assign n5655 = ~n5652 & n5654;
  assign n5656 = ~n5650 & ~n5655;
  assign n5657 = ~n5644 & ~n5656;
  assign n5658 = ~x152 & ~x156;
  assign n5659 = n5658 ^ n5649;
  assign n5660 = n5659 ^ n5649;
  assign n5661 = x151 & ~n5634;
  assign n5662 = n5661 ^ n5649;
  assign n5663 = n5662 ^ n5649;
  assign n5664 = n5660 & ~n5663;
  assign n5665 = n5664 ^ n5649;
  assign n5666 = ~n5637 & n5665;
  assign n5667 = n5666 ^ n5649;
  assign n5668 = ~x155 & n5667;
  assign n5669 = n5657 & ~n5668;
  assign n6470 = n5630 & n5669;
  assign n6468 = ~n5642 & ~n5656;
  assign n6467 = ~n5585 & ~n5620;
  assign n6469 = n6468 ^ n6467;
  assign n6471 = n6470 ^ n6469;
  assign n6480 = n6479 ^ n6471;
  assign n5752 = n5751 ^ n5671;
  assign n5670 = n5669 ^ n5630;
  assign n5753 = n5752 ^ n5670;
  assign n3138 = x156 ^ x155;
  assign n3137 = x154 ^ x153;
  assign n3139 = n3138 ^ n3137;
  assign n3136 = x152 ^ x151;
  assign n3140 = n3139 ^ n3136;
  assign n3132 = x162 ^ x161;
  assign n3134 = n3133 ^ n3132;
  assign n3131 = x158 ^ x157;
  assign n3135 = n3134 ^ n3131;
  assign n3141 = n3140 ^ n3135;
  assign n3152 = n3151 ^ n3146;
  assign n5569 = n3152 ^ n3140;
  assign n5570 = ~n3141 & n5569;
  assign n5571 = n5570 ^ n3152;
  assign n6464 = n5670 ^ n5571;
  assign n6465 = n5753 & ~n6464;
  assign n6466 = n6465 ^ n5752;
  assign n6481 = n6480 ^ n6466;
  assign n5568 = n5567 ^ n5489;
  assign n3153 = n3152 ^ n3141;
  assign n5095 = n3153 & n3176;
  assign n6454 = n5568 ^ n5095;
  assign n6455 = n3135 & n3140;
  assign n6456 = n6455 ^ n5753;
  assign n6457 = n6456 ^ n5095;
  assign n6458 = n6457 ^ n6456;
  assign n5754 = n5753 ^ n5571;
  assign n6459 = n6456 ^ n5754;
  assign n6460 = ~n6458 & ~n6459;
  assign n6461 = n6460 ^ n6456;
  assign n6462 = ~n6454 & n6461;
  assign n6463 = n6462 ^ n5568;
  assign n6482 = n6481 ^ n6463;
  assign n6452 = n6451 ^ n6440;
  assign n6436 = n6435 ^ n6427;
  assign n6453 = n6452 ^ n6436;
  assign n7006 = n6463 ^ n6453;
  assign n7007 = ~n6482 & n7006;
  assign n7008 = n7007 ^ n6481;
  assign n7009 = n6479 ^ n6466;
  assign n7010 = ~n6480 & n7009;
  assign n7011 = n7010 ^ n6466;
  assign n7015 = n6470 ^ n6468;
  assign n7016 = ~n6469 & ~n7015;
  assign n7017 = n7016 ^ n6470;
  assign n7380 = ~n7011 & ~n7017;
  assign n7381 = ~n7008 & n7380;
  assign n7382 = ~n7037 & ~n7381;
  assign n7383 = ~n7379 & ~n7382;
  assign n7384 = ~n7014 & ~n7383;
  assign n7385 = n7379 & ~n7380;
  assign n7386 = n7011 & n7017;
  assign n7387 = n7008 & n7386;
  assign n7388 = ~n7385 & ~n7387;
  assign n7389 = n7384 & n7388;
  assign n7018 = n7017 ^ n7014;
  assign n7019 = n7018 ^ n7011;
  assign n7390 = n7019 & ~n7386;
  assign n7391 = ~n7008 & n7390;
  assign n7392 = ~n7378 & ~n7391;
  assign n7393 = n7037 & ~n7392;
  assign n7400 = n7011 ^ n7008;
  assign n7401 = n7017 ^ n7011;
  assign n7402 = n7400 & ~n7401;
  assign n7403 = n7402 ^ n7008;
  assign n7404 = ~n7379 & ~n7403;
  assign n7559 = ~n7393 & ~n7404;
  assign n7560 = ~n7389 & n7559;
  assign n5287 = x105 & x106;
  assign n5285 = ~x107 & ~x108;
  assign n5286 = x104 & ~n5285;
  assign n5288 = n5287 ^ n5286;
  assign n5289 = x107 & x108;
  assign n5290 = ~x105 & ~x106;
  assign n5291 = n5289 & ~n5290;
  assign n5292 = n5291 ^ n5286;
  assign n5293 = n5292 ^ n5291;
  assign n5294 = n5291 ^ n5289;
  assign n5295 = ~n5293 & ~n5294;
  assign n5296 = n5295 ^ n5291;
  assign n5297 = n5288 & n5296;
  assign n5298 = n5297 ^ n5287;
  assign n5314 = ~n5287 & ~n5291;
  assign n5315 = x103 & ~n5285;
  assign n5316 = ~n5314 & n5315;
  assign n5317 = x103 & x104;
  assign n5318 = ~n5316 & ~n5317;
  assign n5299 = ~n5289 & n5290;
  assign n5319 = ~n5285 & ~n5287;
  assign n5320 = ~n5299 & n5319;
  assign n5321 = ~x108 & n5287;
  assign n5322 = x104 & ~n5321;
  assign n5323 = ~n5320 & n5322;
  assign n5324 = ~n5318 & ~n5323;
  assign n6417 = ~n5298 & ~n5324;
  assign n5300 = n5299 ^ n5285;
  assign n5301 = n5299 ^ n5287;
  assign n5302 = n5285 ^ x104;
  assign n5303 = n5302 ^ n5299;
  assign n5304 = ~n5299 & ~n5303;
  assign n5305 = n5304 ^ n5299;
  assign n5306 = ~n5301 & ~n5305;
  assign n5307 = n5306 ^ n5304;
  assign n5308 = n5307 ^ n5299;
  assign n5309 = n5308 ^ n5302;
  assign n5310 = n5300 & ~n5309;
  assign n5311 = n5310 ^ n5299;
  assign n5312 = ~n5298 & ~n5311;
  assign n5313 = ~x103 & ~n5312;
  assign n5325 = ~n5313 & ~n5324;
  assign n3125 = x106 ^ x105;
  assign n5326 = n5317 ^ x106;
  assign n5327 = n5326 ^ n5317;
  assign n5328 = ~x104 & ~x108;
  assign n5329 = n5328 ^ n5317;
  assign n5330 = ~n5327 & n5329;
  assign n5331 = n5330 ^ n5317;
  assign n5332 = ~n3125 & n5331;
  assign n5333 = ~x107 & n5332;
  assign n5334 = n5325 & ~n5333;
  assign n5247 = ~x111 & ~x112;
  assign n5248 = ~x113 & ~x114;
  assign n5249 = ~n5247 & ~n5248;
  assign n5250 = x111 & x112;
  assign n5251 = x113 & x114;
  assign n5252 = ~n5250 & ~n5251;
  assign n5253 = ~n5249 & n5252;
  assign n3120 = x112 ^ x111;
  assign n3119 = x114 ^ x113;
  assign n3121 = n3120 ^ n3119;
  assign n5254 = x110 & n3121;
  assign n5255 = n5253 & ~n5254;
  assign n5256 = n5251 ^ n5250;
  assign n5257 = n5251 ^ n5249;
  assign n5258 = n5257 ^ n5251;
  assign n5259 = n5251 ^ x110;
  assign n5260 = n5259 ^ n5251;
  assign n5261 = n5258 & n5260;
  assign n5262 = n5261 ^ n5251;
  assign n5263 = n5256 & ~n5262;
  assign n5264 = n5263 ^ n5250;
  assign n5265 = ~n5255 & ~n5264;
  assign n5266 = ~x109 & ~n5265;
  assign n3118 = x110 ^ x109;
  assign n5267 = n5249 & ~n5252;
  assign n5268 = n3118 & n5267;
  assign n5269 = x109 & x110;
  assign n5270 = n5250 & n5269;
  assign n5271 = x114 & n5270;
  assign n5272 = n5271 ^ n5269;
  assign n5273 = ~n5253 & n5272;
  assign n5274 = ~n5268 & ~n5273;
  assign n5275 = n5269 ^ x112;
  assign n5276 = n5275 ^ n5269;
  assign n5277 = ~x110 & ~x114;
  assign n5278 = n5277 ^ n5269;
  assign n5279 = ~n5276 & n5278;
  assign n5280 = n5279 ^ n5269;
  assign n5281 = ~n3120 & n5280;
  assign n5282 = ~x113 & n5281;
  assign n5283 = n5274 & ~n5282;
  assign n5284 = ~n5266 & n5283;
  assign n5335 = n5334 ^ n5284;
  assign n3122 = n3121 ^ n3118;
  assign n3124 = x108 ^ x107;
  assign n3126 = n3125 ^ n3124;
  assign n3123 = x104 ^ x103;
  assign n3127 = n3126 ^ n3123;
  assign n6390 = n3122 & n3127;
  assign n6414 = n6390 ^ n5284;
  assign n6415 = n5335 & ~n6414;
  assign n6416 = n6415 ^ n5334;
  assign n6418 = n6417 ^ n6416;
  assign n6413 = ~n5264 & n5274;
  assign n6419 = n6418 ^ n6413;
  assign n5364 = x117 & x118;
  assign n5365 = x119 & x120;
  assign n5366 = ~n5364 & ~n5365;
  assign n5367 = ~x117 & ~x118;
  assign n5368 = ~x119 & ~x120;
  assign n5369 = ~n5367 & ~n5368;
  assign n5370 = ~n5366 & n5369;
  assign n5371 = x116 & n5370;
  assign n5372 = n5364 & n5365;
  assign n5373 = ~n5371 & ~n5372;
  assign n5374 = n5366 & ~n5369;
  assign n5375 = ~x116 & n5374;
  assign n5376 = n5373 & ~n5375;
  assign n5377 = ~x115 & ~n5376;
  assign n3109 = x116 ^ x115;
  assign n5378 = n5367 & n5368;
  assign n5379 = n3109 & n5378;
  assign n5380 = n5370 ^ x116;
  assign n5381 = n5380 ^ n5370;
  assign n5382 = ~n5372 & ~n5374;
  assign n5383 = n5382 ^ n5370;
  assign n5384 = n5381 & n5383;
  assign n5385 = n5384 ^ n5370;
  assign n5386 = x115 & n5385;
  assign n5387 = ~n5379 & ~n5386;
  assign n5388 = ~n5377 & n5387;
  assign n5337 = ~x123 & ~x124;
  assign n5338 = x125 & x126;
  assign n5339 = n5337 & ~n5338;
  assign n5340 = ~x125 & ~x126;
  assign n5341 = x122 & ~n5340;
  assign n5342 = n5339 & ~n5341;
  assign n5343 = x123 & x124;
  assign n5344 = n5338 & n5343;
  assign n5345 = ~n5342 & ~n5344;
  assign n5346 = ~x121 & ~n5345;
  assign n3114 = x122 ^ x121;
  assign n3113 = x126 ^ x125;
  assign n3115 = n3114 ^ n3113;
  assign n3112 = x124 ^ x123;
  assign n3116 = n3115 ^ n3112;
  assign n5347 = ~x122 & n5340;
  assign n5348 = ~n5343 & n5347;
  assign n5349 = n3116 & n5348;
  assign n5350 = x121 & x122;
  assign n5351 = n5343 & n5350;
  assign n5352 = ~n5338 & n5351;
  assign n5353 = ~n5349 & ~n5352;
  assign n5354 = ~n5346 & n5353;
  assign n5355 = ~n5343 & n5350;
  assign n5356 = ~n5339 & n5355;
  assign n5357 = n5338 ^ x124;
  assign n5358 = n3112 & n5357;
  assign n5359 = n5358 ^ x124;
  assign n5360 = n3114 & n5359;
  assign n5361 = ~n5356 & ~n5360;
  assign n5362 = ~n5340 & ~n5361;
  assign n5363 = n5354 & ~n5362;
  assign n5389 = n5388 ^ n5363;
  assign n3108 = x118 ^ x117;
  assign n3110 = n3109 ^ n3108;
  assign n3107 = x120 ^ x119;
  assign n3111 = n3110 ^ n3107;
  assign n6397 = n3111 & n3116;
  assign n6409 = n5389 & n6397;
  assign n6410 = n5363 & n5388;
  assign n6411 = ~n6409 & ~n6410;
  assign n6407 = n5373 & ~n5386;
  assign n6405 = ~n5344 & ~n5351;
  assign n6406 = ~n5362 & n6405;
  assign n6408 = n6407 ^ n6406;
  assign n6412 = n6411 ^ n6408;
  assign n6420 = n6419 ^ n6412;
  assign n6391 = n5335 & n6390;
  assign n3128 = n3127 ^ n3122;
  assign n3117 = n3116 ^ n3111;
  assign n3129 = n3128 ^ n3117;
  assign n6392 = ~n3111 & ~n6390;
  assign n6393 = n3129 & n6392;
  assign n6394 = ~n3122 & ~n3127;
  assign n6395 = ~n6393 & ~n6394;
  assign n6396 = ~n5335 & ~n6395;
  assign n6398 = n6397 ^ n5389;
  assign n6399 = n6398 ^ n6397;
  assign n5242 = n3122 ^ n3116;
  assign n5244 = n5242 ^ n3111;
  assign n5245 = ~n3127 & n5244;
  assign n5243 = ~n3117 & ~n5242;
  assign n5246 = n5245 ^ n5243;
  assign n5336 = n5335 ^ n5246;
  assign n6400 = n6397 ^ n5336;
  assign n6401 = ~n6399 & ~n6400;
  assign n6402 = n6401 ^ n6397;
  assign n6403 = ~n6396 & ~n6402;
  assign n6404 = ~n6391 & n6403;
  assign n6421 = n6420 ^ n6404;
  assign n6972 = n6417 ^ n6404;
  assign n6973 = ~n6418 & n6972;
  assign n6974 = n6973 ^ n6416;
  assign n6975 = n6413 & ~n6974;
  assign n6976 = ~n6421 & n6975;
  assign n6977 = ~n6416 & n6417;
  assign n6978 = n6412 & n6977;
  assign n6979 = ~n6404 & n6978;
  assign n6980 = ~n6976 & ~n6979;
  assign n6969 = n6411 ^ n6407;
  assign n6970 = ~n6408 & n6969;
  assign n6971 = n6970 ^ n6411;
  assign n6981 = ~n6412 & n6974;
  assign n6982 = n6421 & n6981;
  assign n7372 = n6971 & ~n6982;
  assign n7373 = n6980 & ~n7372;
  assign n3086 = x98 ^ x97;
  assign n3085 = x100 ^ x99;
  assign n3087 = n3086 ^ n3085;
  assign n3084 = x102 ^ x101;
  assign n3088 = n3087 ^ n3084;
  assign n3091 = x92 ^ x91;
  assign n3090 = x94 ^ x93;
  assign n3092 = n3091 ^ n3090;
  assign n3089 = x96 ^ x95;
  assign n3093 = n3092 ^ n3089;
  assign n5104 = n3088 & n3093;
  assign n5147 = x95 & x96;
  assign n5148 = ~x93 & ~x94;
  assign n5149 = ~n5147 & n5148;
  assign n5150 = ~x95 & ~x96;
  assign n5151 = x92 & ~n5150;
  assign n5152 = n5149 & ~n5151;
  assign n5153 = x93 & x94;
  assign n5154 = n5147 & n5153;
  assign n5155 = ~n5152 & ~n5154;
  assign n5156 = ~x91 & ~n5155;
  assign n5157 = ~x92 & n5150;
  assign n5158 = ~n5153 & n5157;
  assign n5159 = n3092 & n5158;
  assign n5160 = x91 & x92;
  assign n5161 = n5153 & n5160;
  assign n5162 = ~n5147 & n5161;
  assign n5163 = ~n5159 & ~n5162;
  assign n5164 = ~n5156 & n5163;
  assign n5165 = ~n5153 & n5160;
  assign n5166 = ~n5149 & n5165;
  assign n5167 = n5147 ^ x94;
  assign n5168 = n3090 & n5167;
  assign n5169 = n5168 ^ x94;
  assign n5170 = n3091 & n5169;
  assign n5171 = ~n5166 & ~n5170;
  assign n5172 = ~n5150 & ~n5171;
  assign n5173 = n5164 & ~n5172;
  assign n5120 = x101 & x102;
  assign n5121 = ~x99 & ~x100;
  assign n5122 = ~n5120 & n5121;
  assign n5123 = ~x101 & ~x102;
  assign n5124 = x98 & ~n5123;
  assign n5125 = n5122 & ~n5124;
  assign n5126 = x99 & x100;
  assign n5127 = n5120 & n5126;
  assign n5128 = ~n5125 & ~n5127;
  assign n5129 = ~x97 & ~n5128;
  assign n5130 = ~x98 & n5123;
  assign n5131 = ~n5126 & n5130;
  assign n5132 = n3087 & n5131;
  assign n5133 = x97 & x98;
  assign n5134 = n5126 & n5133;
  assign n5135 = ~n5120 & n5134;
  assign n5136 = ~n5132 & ~n5135;
  assign n5137 = ~n5129 & n5136;
  assign n5138 = ~n5126 & n5133;
  assign n5139 = ~n5122 & n5138;
  assign n5140 = n5120 ^ x100;
  assign n5141 = n3085 & n5140;
  assign n5142 = n5141 ^ x100;
  assign n5143 = n3086 & n5142;
  assign n5144 = ~n5139 & ~n5143;
  assign n5145 = ~n5123 & ~n5144;
  assign n5146 = n5137 & ~n5145;
  assign n5174 = n5173 ^ n5146;
  assign n6370 = n5104 & n5174;
  assign n6371 = n5146 & n5173;
  assign n6372 = ~n6370 & ~n6371;
  assign n6367 = ~n5154 & ~n5161;
  assign n6368 = ~n5172 & n6367;
  assign n6365 = ~n5127 & ~n5134;
  assign n6366 = ~n5145 & n6365;
  assign n6369 = n6368 ^ n6366;
  assign n6373 = n6372 ^ n6369;
  assign n5205 = x83 & x84;
  assign n5206 = x81 & x82;
  assign n5207 = n5205 & n5206;
  assign n5208 = ~x83 & ~x84;
  assign n5209 = x80 & ~n5208;
  assign n5210 = ~n5207 & ~n5209;
  assign n3101 = x82 ^ x81;
  assign n5211 = n5205 ^ x82;
  assign n5212 = n3101 & ~n5211;
  assign n5213 = n5212 ^ x81;
  assign n5214 = ~n5210 & n5213;
  assign n5225 = ~n5208 & n5213;
  assign n5226 = ~x80 & ~n5225;
  assign n5217 = ~x81 & ~x82;
  assign n5218 = ~n5205 & n5217;
  assign n5227 = ~n5207 & ~n5218;
  assign n5215 = ~n5206 & n5208;
  assign n5228 = n5227 ^ n5215;
  assign n5229 = n5227 ^ x79;
  assign n5230 = n5227 & n5229;
  assign n5231 = n5230 ^ n5227;
  assign n5232 = ~n5228 & n5231;
  assign n5233 = n5232 ^ n5230;
  assign n5234 = n5233 ^ n5227;
  assign n5235 = n5234 ^ x79;
  assign n5236 = x80 & n5235;
  assign n5237 = n5236 ^ x79;
  assign n5238 = ~n5226 & n5237;
  assign n6385 = ~n5214 & ~n5238;
  assign n5179 = x87 & x88;
  assign n5180 = x89 & x90;
  assign n5184 = n5179 & n5180;
  assign n5187 = x85 & x86;
  assign n5190 = ~n5184 & n5187;
  assign n5181 = ~n5179 & ~n5180;
  assign n5191 = n5190 ^ n5181;
  assign n3097 = x86 ^ x85;
  assign n5192 = n5190 ^ n3097;
  assign n5176 = ~x87 & ~x88;
  assign n5177 = ~x89 & ~x90;
  assign n5178 = ~n5176 & ~n5177;
  assign n5193 = n5181 ^ n5178;
  assign n5194 = n5193 ^ n3097;
  assign n5195 = ~n3097 & ~n5194;
  assign n5196 = n5195 ^ n3097;
  assign n5197 = n5192 & ~n5196;
  assign n5198 = n5197 ^ n5195;
  assign n5199 = n5198 ^ n3097;
  assign n5200 = n5199 ^ n5193;
  assign n5201 = ~n5191 & ~n5200;
  assign n5202 = n5201 ^ n5190;
  assign n6384 = ~n5184 & ~n5202;
  assign n6386 = n6385 ^ n6384;
  assign n5216 = ~x80 & n5215;
  assign n5219 = ~n5209 & n5218;
  assign n5220 = ~n5216 & ~n5219;
  assign n5221 = ~n5214 & n5220;
  assign n5222 = ~x79 & ~n5221;
  assign n5223 = n5216 & n5217;
  assign n5224 = ~n5222 & ~n5223;
  assign n5239 = n5224 & ~n5238;
  assign n5182 = ~n5178 & n5181;
  assign n5183 = ~x86 & n5182;
  assign n5185 = ~n5183 & ~n5184;
  assign n5186 = ~x85 & ~n5185;
  assign n5188 = n5176 & ~n5187;
  assign n5189 = n5177 & n5188;
  assign n5203 = ~n5189 & ~n5202;
  assign n5204 = ~n5186 & n5203;
  assign n5240 = n5239 ^ n5204;
  assign n3096 = x88 ^ x87;
  assign n3098 = n3097 ^ n3096;
  assign n3095 = x90 ^ x89;
  assign n3099 = n3098 ^ n3095;
  assign n3102 = x84 ^ x83;
  assign n3103 = n3102 ^ n3101;
  assign n3100 = x80 ^ x79;
  assign n3104 = n3103 ^ n3100;
  assign n5103 = n3099 & n3104;
  assign n6381 = n5204 ^ n5103;
  assign n6382 = n5240 & ~n6381;
  assign n6383 = n6382 ^ n5239;
  assign n6387 = n6386 ^ n6383;
  assign n6374 = n5103 & n5240;
  assign n5105 = n5103 & n5104;
  assign n3094 = n3093 ^ n3088;
  assign n5106 = n3104 ^ n3094;
  assign n3105 = n3104 ^ n3099;
  assign n5107 = n5106 ^ n3105;
  assign n5108 = n3099 ^ n3093;
  assign n5109 = n5108 ^ n3104;
  assign n5110 = n5109 ^ n3104;
  assign n5111 = ~n3094 & n5110;
  assign n5112 = n5111 ^ n3094;
  assign n5113 = n5109 & ~n5112;
  assign n5114 = n5113 ^ n3104;
  assign n5115 = n5107 & n5114;
  assign n5116 = n5115 ^ n5111;
  assign n5117 = n5116 ^ n3104;
  assign n5118 = n5117 ^ n3105;
  assign n5119 = ~n5105 & n5118;
  assign n5175 = n5174 ^ n5119;
  assign n6375 = n5175 & ~n5240;
  assign n6376 = n5118 ^ n5104;
  assign n6377 = ~n5174 & ~n6376;
  assign n6378 = n6377 ^ n5104;
  assign n6379 = ~n6375 & ~n6378;
  assign n6380 = ~n6374 & n6379;
  assign n6388 = n6387 ^ n6380;
  assign n6996 = n6373 & n6388;
  assign n6991 = ~n6383 & n6385;
  assign n6997 = n6996 ^ n6991;
  assign n6992 = ~n6380 & n6384;
  assign n6998 = n6992 ^ n6991;
  assign n6999 = n6997 & ~n6998;
  assign n7000 = n6999 ^ n6996;
  assign n6988 = n6372 ^ n6368;
  assign n6989 = ~n6369 & n6988;
  assign n6990 = n6989 ^ n6372;
  assign n6993 = ~n6991 & ~n6992;
  assign n6994 = ~n6373 & n6388;
  assign n6995 = n6993 & n6994;
  assign n7370 = n6990 & ~n6995;
  assign n7371 = ~n7000 & ~n7370;
  assign n7374 = n7373 ^ n7371;
  assign n7001 = ~n6995 & ~n7000;
  assign n7002 = n7001 ^ n6990;
  assign n6389 = n6388 ^ n6373;
  assign n6422 = n6421 ^ n6389;
  assign n5390 = n5389 ^ n5336;
  assign n5241 = n5240 ^ n5175;
  assign n5391 = n5390 ^ n5241;
  assign n3106 = n3105 ^ n3094;
  assign n5099 = n3106 & n3129;
  assign n6362 = n5241 ^ n5099;
  assign n6363 = ~n5391 & ~n6362;
  assign n6364 = n6363 ^ n5390;
  assign n6985 = n6389 ^ n6364;
  assign n6986 = n6422 & ~n6985;
  assign n6987 = n6986 ^ n6421;
  assign n7003 = n7002 ^ n6987;
  assign n6983 = n6980 & ~n6982;
  assign n6984 = n6983 ^ n6971;
  assign n7367 = n6987 ^ n6984;
  assign n7368 = n7003 & ~n7367;
  assign n7369 = n7368 ^ n7002;
  assign n7556 = n7373 ^ n7369;
  assign n7557 = ~n7374 & ~n7556;
  assign n7558 = n7557 ^ n7369;
  assign n7561 = n7560 ^ n7558;
  assign n7375 = n7374 ^ n7369;
  assign n7004 = n7003 ^ n6984;
  assign n6423 = n6422 ^ n6364;
  assign n6350 = n5099 & ~n5391;
  assign n6351 = n5095 & n5099;
  assign n3130 = n3129 ^ n3106;
  assign n3177 = n3176 ^ n3153;
  assign n5096 = n3177 ^ n3106;
  assign n5097 = n3130 & ~n5096;
  assign n5098 = n5097 ^ n3129;
  assign n5100 = n5099 ^ n5098;
  assign n5101 = ~n5095 & ~n5100;
  assign n5102 = n5101 ^ n5099;
  assign n6352 = ~n5102 & ~n5391;
  assign n6353 = ~n6351 & ~n6352;
  assign n5755 = n5754 ^ n5568;
  assign n6354 = n6353 ^ n5755;
  assign n6355 = n6354 ^ n6353;
  assign n6356 = ~n5098 & n5391;
  assign n6357 = ~n5095 & ~n6356;
  assign n6358 = n6357 ^ n6353;
  assign n6359 = ~n6355 & ~n6358;
  assign n6360 = n6359 ^ n6353;
  assign n6361 = ~n6350 & ~n6360;
  assign n6424 = n6423 ^ n6361;
  assign n6483 = n6482 ^ n6453;
  assign n6966 = n6483 ^ n6423;
  assign n6967 = ~n6424 & ~n6966;
  assign n6968 = n6967 ^ n6361;
  assign n7005 = n7004 ^ n6968;
  assign n7020 = n7019 ^ n7008;
  assign n7038 = n7037 ^ n7020;
  assign n7364 = n7038 ^ n6968;
  assign n7365 = ~n7005 & n7364;
  assign n7366 = n7365 ^ n7004;
  assign n7376 = n7375 ^ n7366;
  assign n7394 = n7378 & ~n7381;
  assign n7395 = n7037 & ~n7394;
  assign n7396 = n7014 & ~n7395;
  assign n7397 = n7396 ^ n7393;
  assign n7398 = n7379 & n7386;
  assign n7399 = n7398 ^ n7393;
  assign n7405 = n7404 ^ n7393;
  assign n7406 = ~n7393 & n7405;
  assign n7407 = n7406 ^ n7393;
  assign n7408 = ~n7399 & ~n7407;
  assign n7409 = n7408 ^ n7406;
  assign n7410 = n7409 ^ n7393;
  assign n7411 = n7410 ^ n7404;
  assign n7412 = n7397 & n7411;
  assign n7413 = n7412 ^ n7396;
  assign n7414 = ~n7389 & ~n7413;
  assign n7553 = n7414 ^ n7366;
  assign n7554 = ~n7376 & n7553;
  assign n7555 = n7554 ^ n7414;
  assign n7562 = n7561 ^ n7555;
  assign n7610 = n7609 ^ n7562;
  assign n7415 = n7414 ^ n7376;
  assign n7549 = n7415 ^ n7362;
  assign n6964 = n6963 ^ n6890;
  assign n6484 = n6483 ^ n6424;
  assign n6340 = n5093 ^ n4528;
  assign n5392 = n5391 ^ n5102;
  assign n5756 = n5755 ^ n5392;
  assign n6341 = n6340 ^ n5756;
  assign n6342 = n5756 ^ n4528;
  assign n6343 = n6342 ^ n5756;
  assign n3178 = n3177 ^ n3130;
  assign n4529 = ~n3035 & ~n3082;
  assign n4530 = n3178 & ~n4529;
  assign n6344 = n5756 ^ n4530;
  assign n6345 = n6344 ^ n5756;
  assign n6346 = ~n6343 & n6345;
  assign n6347 = n6346 ^ n5756;
  assign n6348 = n6341 & ~n6347;
  assign n6349 = n6348 ^ n5756;
  assign n6485 = n6484 ^ n6349;
  assign n6602 = n6601 ^ n6589;
  assign n6885 = n6602 ^ n6484;
  assign n6886 = n6485 & n6885;
  assign n6887 = n6886 ^ n6602;
  assign n6965 = n6964 ^ n6887;
  assign n7039 = n7038 ^ n7005;
  assign n7335 = n7039 ^ n6887;
  assign n7336 = n6965 & ~n7335;
  assign n7337 = n7336 ^ n6964;
  assign n7550 = n7415 ^ n7337;
  assign n7551 = n7549 & n7550;
  assign n7552 = n7551 ^ n7362;
  assign n7611 = n7610 ^ n7552;
  assign n7498 = n7497 ^ n7448;
  assign n7363 = n7362 ^ n7337;
  assign n7416 = n7415 ^ n7363;
  assign n7499 = n7498 ^ n7416;
  assign n7040 = n7039 ^ n6965;
  assign n6338 = n6337 ^ n6217;
  assign n4531 = ~n4528 & ~n4530;
  assign n5094 = n5093 ^ n4531;
  assign n5757 = n5756 ^ n5094;
  assign n2988 = n2987 ^ n2892;
  assign n3083 = n3082 ^ n3035;
  assign n3179 = n3178 ^ n3083;
  assign n3180 = n2988 & n3179;
  assign n6093 = n5757 ^ n3180;
  assign n3831 = ~n3829 & ~n3830;
  assign n4526 = n4525 ^ n3831;
  assign n4527 = n4526 ^ n3828;
  assign n6094 = n4527 ^ n3180;
  assign n6095 = ~n6093 & n6094;
  assign n6096 = n6095 ^ n5757;
  assign n6339 = n6338 ^ n6096;
  assign n6603 = n6602 ^ n6485;
  assign n6882 = n6603 ^ n6096;
  assign n6883 = n6339 & ~n6882;
  assign n6884 = n6883 ^ n6338;
  assign n7041 = n7040 ^ n6884;
  assign n7211 = n7210 ^ n7130;
  assign n7332 = n7211 ^ n6884;
  assign n7333 = ~n7041 & n7332;
  assign n7334 = n7333 ^ n7040;
  assign n7546 = n7416 ^ n7334;
  assign n7547 = ~n7499 & ~n7546;
  assign n7548 = n7547 ^ n7498;
  assign n7612 = n7611 ^ n7548;
  assign n7674 = n7673 ^ n7626;
  assign n7623 = n7622 ^ n7615;
  assign n7675 = n7674 ^ n7623;
  assign n7709 = n7675 ^ n7611;
  assign n7710 = ~n7612 & n7709;
  assign n7711 = n7710 ^ n7675;
  assign n7729 = ~n7672 & ~n7724;
  assign n7730 = ~n7642 & ~n7729;
  assign n7732 = ~n7724 & ~n7731;
  assign n7733 = n7732 ^ n7716;
  assign n7734 = n7730 & n7733;
  assign n7735 = ~n7728 & ~n7734;
  assign n7781 = ~n7711 & ~n7735;
  assign n7795 = ~n7751 & ~n7781;
  assign n7796 = n7700 & ~n7795;
  assign n7701 = n7560 ^ n7555;
  assign n7702 = n7561 & ~n7701;
  assign n7703 = n7702 ^ n7555;
  assign n7704 = n7562 ^ n7552;
  assign n7705 = n7610 & n7704;
  assign n7706 = n7705 ^ n7609;
  assign n7784 = ~n7703 & n7706;
  assign n7754 = n7711 & n7735;
  assign n7797 = n7751 & ~n7754;
  assign n7798 = ~n7784 & ~n7797;
  assign n7799 = ~n7796 & n7798;
  assign n7780 = n7703 & ~n7706;
  assign n7800 = n7780 ^ n7751;
  assign n7801 = n7700 & ~n7754;
  assign n7802 = n7801 ^ n7751;
  assign n7803 = n7802 ^ n7751;
  assign n7804 = n7781 ^ n7751;
  assign n7805 = n7804 ^ n7751;
  assign n7806 = ~n7803 & ~n7805;
  assign n7807 = n7806 ^ n7751;
  assign n7808 = ~n7800 & n7807;
  assign n7809 = n7808 ^ n7780;
  assign n7810 = ~n7799 & ~n7809;
  assign n2370 = x53 & x54;
  assign n2371 = x51 & x52;
  assign n2372 = ~n2370 & ~n2371;
  assign n2373 = ~x53 & ~x54;
  assign n2374 = ~x51 & ~x52;
  assign n2375 = ~n2373 & ~n2374;
  assign n2376 = ~n2372 & n2375;
  assign n2377 = x50 & n2376;
  assign n2378 = n2370 & n2371;
  assign n2379 = ~n2377 & ~n2378;
  assign n2380 = n2372 & ~n2375;
  assign n2381 = ~x50 & n2380;
  assign n2382 = n2379 & ~n2381;
  assign n2383 = ~x49 & ~n2382;
  assign n1146 = x50 ^ x49;
  assign n2384 = n2373 & n2374;
  assign n2385 = n1146 & n2384;
  assign n2386 = n2376 ^ x50;
  assign n2387 = n2386 ^ n2376;
  assign n2388 = ~n2378 & ~n2380;
  assign n2389 = n2388 ^ n2376;
  assign n2390 = n2387 & n2389;
  assign n2391 = n2390 ^ n2376;
  assign n2392 = x49 & n2391;
  assign n2393 = ~n2385 & ~n2392;
  assign n2394 = ~n2383 & n2393;
  assign n2326 = x47 & x48;
  assign n2325 = x45 & x46;
  assign n2327 = n2326 ^ n2325;
  assign n2328 = ~x47 & ~x48;
  assign n2329 = ~x45 & ~x46;
  assign n2330 = ~n2328 & ~n2329;
  assign n2331 = n2330 ^ n2325;
  assign n2332 = n2331 ^ n2325;
  assign n2333 = n2325 ^ x44;
  assign n2334 = n2333 ^ n2325;
  assign n2335 = n2332 & n2334;
  assign n2336 = n2335 ^ n2325;
  assign n2337 = n2327 & ~n2336;
  assign n2338 = n2337 ^ n2326;
  assign n2339 = n2329 ^ n2328;
  assign n2340 = ~n2325 & ~n2326;
  assign n2341 = n2340 ^ n2329;
  assign n2342 = n2341 ^ n2329;
  assign n2343 = n2329 ^ x44;
  assign n2344 = n2343 ^ n2329;
  assign n2345 = n2342 & ~n2344;
  assign n2346 = n2345 ^ n2329;
  assign n2347 = n2339 & ~n2346;
  assign n2348 = n2347 ^ n2328;
  assign n2349 = ~n2338 & ~n2348;
  assign n2350 = ~x43 & ~n2349;
  assign n1151 = x44 ^ x43;
  assign n2351 = n2330 & ~n2340;
  assign n2352 = n1151 & n2351;
  assign n2353 = ~n2330 & n2340;
  assign n2354 = x43 & x44;
  assign n2355 = n2325 & n2354;
  assign n2356 = x48 & n2355;
  assign n2357 = n2356 ^ n2354;
  assign n2358 = ~n2353 & n2357;
  assign n2359 = ~n2352 & ~n2358;
  assign n1150 = x46 ^ x45;
  assign n2360 = n2354 ^ x46;
  assign n2361 = n2360 ^ n2354;
  assign n2362 = ~x44 & ~x48;
  assign n2363 = n2362 ^ n2354;
  assign n2364 = ~n2361 & n2363;
  assign n2365 = n2364 ^ n2354;
  assign n2366 = ~n1150 & n2365;
  assign n2367 = ~x47 & n2366;
  assign n2368 = n2359 & ~n2367;
  assign n2369 = ~n2350 & n2368;
  assign n2395 = n2394 ^ n2369;
  assign n2465 = x39 & x40;
  assign n2464 = x41 & x42;
  assign n2466 = n2465 ^ n2464;
  assign n2467 = ~x39 & ~x40;
  assign n2468 = ~x41 & ~x42;
  assign n2469 = ~n2467 & ~n2468;
  assign n2470 = n2469 ^ n2464;
  assign n2471 = n2470 ^ n2464;
  assign n2472 = n2464 ^ x38;
  assign n2473 = n2472 ^ n2464;
  assign n2474 = n2471 & n2473;
  assign n2475 = n2474 ^ n2464;
  assign n2476 = n2466 & ~n2475;
  assign n2477 = n2476 ^ n2465;
  assign n1160 = x42 ^ x41;
  assign n2478 = x41 ^ x38;
  assign n2479 = n1160 & n2478;
  assign n2480 = n2479 ^ x41;
  assign n2481 = n2467 & ~n2480;
  assign n2482 = ~n2477 & ~n2481;
  assign n2483 = ~x37 & ~n2482;
  assign n2484 = x37 & x38;
  assign n1162 = x38 ^ x37;
  assign n1161 = x40 ^ x39;
  assign n1163 = n1162 ^ n1161;
  assign n2485 = n2484 ^ n1163;
  assign n2486 = n2485 ^ n2484;
  assign n2487 = ~x38 & ~x42;
  assign n2488 = n2487 ^ n2484;
  assign n2489 = n2488 ^ n2484;
  assign n2490 = n2486 & n2489;
  assign n2491 = n2490 ^ n2484;
  assign n2492 = ~n2465 & n2491;
  assign n2493 = n2492 ^ n2484;
  assign n2494 = ~x41 & n2493;
  assign n2495 = ~n2464 & ~n2465;
  assign n2496 = ~n2469 & n2495;
  assign n2497 = n2465 & n2484;
  assign n2498 = x42 & n2497;
  assign n2499 = n2498 ^ n2484;
  assign n2500 = ~n2496 & n2499;
  assign n2501 = n2469 & ~n2495;
  assign n2502 = n1162 & n2501;
  assign n2503 = ~n2500 & ~n2502;
  assign n2504 = ~n2494 & n2503;
  assign n2505 = ~n2483 & n2504;
  assign n1157 = x34 ^ x33;
  assign n2413 = x31 & x32;
  assign n2414 = n2413 ^ x34;
  assign n2415 = n2414 ^ n2413;
  assign n2416 = ~x32 & ~x36;
  assign n2417 = n2416 ^ n2413;
  assign n2418 = ~n2415 & n2417;
  assign n2419 = n2418 ^ n2413;
  assign n2420 = ~n1157 & n2419;
  assign n2421 = ~x35 & n2420;
  assign n2423 = x33 & x34;
  assign n2422 = x35 & x36;
  assign n2424 = n2423 ^ n2422;
  assign n2425 = ~x33 & ~x34;
  assign n2426 = ~x35 & ~x36;
  assign n2427 = ~n2425 & ~n2426;
  assign n2428 = n2427 ^ n2422;
  assign n2429 = n2428 ^ n2422;
  assign n2430 = n2422 ^ x32;
  assign n2431 = n2430 ^ n2422;
  assign n2432 = n2429 & n2431;
  assign n2433 = n2432 ^ n2422;
  assign n2434 = n2424 & ~n2433;
  assign n2435 = n2434 ^ n2423;
  assign n2436 = n2426 ^ n2425;
  assign n2437 = ~n2422 & ~n2423;
  assign n2438 = n2437 ^ n2426;
  assign n2439 = n2438 ^ n2426;
  assign n2440 = n2426 ^ x32;
  assign n2441 = n2440 ^ n2426;
  assign n2442 = n2439 & ~n2441;
  assign n2443 = n2442 ^ n2426;
  assign n2444 = n2436 & ~n2443;
  assign n2445 = n2444 ^ n2425;
  assign n2446 = ~n2435 & ~n2445;
  assign n2447 = n2446 ^ x31;
  assign n2448 = n2447 ^ n2446;
  assign n2450 = n2427 & ~n2437;
  assign n2449 = x36 & n2423;
  assign n2451 = n2450 ^ n2449;
  assign n2452 = n2451 ^ n2450;
  assign n2453 = ~n2427 & n2437;
  assign n2454 = n2453 ^ n2450;
  assign n2455 = n2454 ^ n2450;
  assign n2456 = ~n2452 & ~n2455;
  assign n2457 = n2456 ^ n2450;
  assign n2458 = x32 & n2457;
  assign n2459 = n2458 ^ n2450;
  assign n2460 = n2459 ^ n2446;
  assign n2461 = n2448 & ~n2460;
  assign n2462 = n2461 ^ n2446;
  assign n2463 = ~n2421 & n2462;
  assign n2506 = n2505 ^ n2463;
  assign n1156 = x36 ^ x35;
  assign n1158 = n1157 ^ n1156;
  assign n1155 = x32 ^ x31;
  assign n1159 = n1158 ^ n1155;
  assign n1164 = n1163 ^ n1160;
  assign n2396 = n1159 & n1164;
  assign n1145 = x52 ^ x51;
  assign n1147 = n1146 ^ n1145;
  assign n1144 = x54 ^ x53;
  assign n1148 = n1147 ^ n1144;
  assign n1152 = n1151 ^ n1150;
  assign n1149 = x48 ^ x47;
  assign n1153 = n1152 ^ n1149;
  assign n2397 = n1148 & n1153;
  assign n2398 = n2396 & n2397;
  assign n1154 = n1153 ^ n1148;
  assign n2399 = n1164 ^ n1154;
  assign n1165 = n1164 ^ n1159;
  assign n2400 = n2399 ^ n1165;
  assign n2401 = n1159 ^ n1153;
  assign n2402 = n2401 ^ n1164;
  assign n2403 = n2402 ^ n1164;
  assign n2404 = ~n1154 & n2403;
  assign n2405 = n2404 ^ n1154;
  assign n2406 = n2402 & ~n2405;
  assign n2407 = n2406 ^ n1164;
  assign n2408 = n2400 & n2407;
  assign n2409 = n2408 ^ n2404;
  assign n2410 = n2409 ^ n1164;
  assign n2411 = n2410 ^ n1165;
  assign n2412 = ~n2398 & n2411;
  assign n2507 = n2506 ^ n2412;
  assign n6001 = n2507 ^ n2397;
  assign n6002 = ~n2395 & n6001;
  assign n6003 = n6002 ^ n2397;
  assign n6004 = n2411 ^ n2396;
  assign n6005 = ~n2506 & ~n6004;
  assign n6006 = n6005 ^ n2396;
  assign n6007 = ~n6003 & ~n6006;
  assign n5997 = n2395 & ~n2397;
  assign n5998 = ~n2369 & ~n2394;
  assign n5999 = ~n5997 & ~n5998;
  assign n5995 = n2379 & ~n2392;
  assign n5994 = ~n2338 & n2359;
  assign n5996 = n5995 ^ n5994;
  assign n6000 = n5999 ^ n5996;
  assign n6008 = n6007 ^ n6000;
  assign n5989 = ~n2396 & n2506;
  assign n5990 = ~n2463 & ~n2505;
  assign n5991 = ~n5989 & ~n5990;
  assign n5987 = x31 & n2459;
  assign n5988 = ~n2435 & ~n5987;
  assign n5992 = n5991 ^ n5988;
  assign n5986 = ~n2477 & n2503;
  assign n5993 = n5992 ^ n5986;
  assign n6645 = n6000 ^ n5993;
  assign n6646 = n6008 & ~n6645;
  assign n6647 = n6646 ^ n6007;
  assign n6648 = n5999 ^ n5995;
  assign n6649 = ~n5996 & ~n6648;
  assign n6650 = n6649 ^ n5999;
  assign n6651 = n5988 ^ n5986;
  assign n6652 = ~n5992 & ~n6651;
  assign n6653 = n6652 ^ n5991;
  assign n7307 = n6650 & n6653;
  assign n7308 = n6647 & n7307;
  assign n1174 = x62 ^ x61;
  assign n2207 = x65 & x66;
  assign n2216 = ~x63 & ~x64;
  assign n2221 = n2207 & ~n2216;
  assign n2211 = x63 & x64;
  assign n2212 = ~x65 & ~x66;
  assign n2222 = n2211 & ~n2212;
  assign n2223 = ~n2221 & ~n2222;
  assign n2224 = n1174 & ~n2223;
  assign n1173 = x64 ^ x63;
  assign n2208 = n2207 ^ x64;
  assign n2209 = ~n1173 & ~n2208;
  assign n2213 = ~n2211 & n2212;
  assign n2225 = x61 & x62;
  assign n2226 = ~n2213 & n2225;
  assign n2227 = ~n2209 & n2226;
  assign n2228 = ~n2224 & ~n2227;
  assign n6013 = n2207 & n2211;
  assign n6014 = n2228 & ~n6013;
  assign n2210 = ~x61 & n2209;
  assign n2214 = ~x62 & n2213;
  assign n2215 = ~n2210 & ~n2214;
  assign n2217 = x61 & ~n2216;
  assign n2218 = x62 & ~n2212;
  assign n2219 = ~n2217 & ~n2218;
  assign n2220 = ~n2215 & n2219;
  assign n2229 = ~n2220 & n2228;
  assign n2177 = x57 & x58;
  assign n2178 = x59 & x60;
  assign n2179 = n2177 & n2178;
  assign n2180 = ~x57 & ~x58;
  assign n2181 = ~n2178 & n2180;
  assign n2182 = n2181 ^ x56;
  assign n2183 = ~x59 & ~x60;
  assign n2184 = n2183 ^ n2181;
  assign n2185 = n2184 ^ n2183;
  assign n2186 = ~n2177 & n2183;
  assign n2187 = n2186 ^ n2183;
  assign n2188 = ~n2185 & ~n2187;
  assign n2189 = n2188 ^ n2183;
  assign n2190 = ~n2182 & n2189;
  assign n2191 = n2190 ^ x56;
  assign n2192 = ~n2179 & n2191;
  assign n2193 = ~x55 & ~n2192;
  assign n2194 = ~n2179 & ~n2186;
  assign n2195 = x55 & x56;
  assign n2196 = ~n2181 & n2195;
  assign n2197 = n2194 & n2196;
  assign n1169 = x56 ^ x55;
  assign n2198 = n2178 & ~n2180;
  assign n2199 = n2177 & ~n2183;
  assign n2200 = ~n2198 & ~n2199;
  assign n2201 = n1169 & ~n2200;
  assign n2202 = ~n2197 & ~n2201;
  assign n2203 = ~x56 & n2186;
  assign n2204 = n2180 & n2203;
  assign n2205 = n2202 & ~n2204;
  assign n2206 = ~n2193 & n2205;
  assign n2230 = n2229 ^ n2206;
  assign n1168 = x58 ^ x57;
  assign n1170 = n1169 ^ n1168;
  assign n1167 = x60 ^ x59;
  assign n1171 = n1170 ^ n1167;
  assign n1175 = n1174 ^ n1173;
  assign n1172 = x66 ^ x65;
  assign n1176 = n1175 ^ n1172;
  assign n2173 = n1171 & n1176;
  assign n6010 = n2206 ^ n2173;
  assign n6011 = n2230 & ~n6010;
  assign n6012 = n6011 ^ n2229;
  assign n6015 = ~n2179 & n2202;
  assign n2278 = x75 & x76;
  assign n2277 = x77 & x78;
  assign n2279 = n2278 ^ n2277;
  assign n2280 = ~x75 & ~x76;
  assign n2281 = ~x77 & ~x78;
  assign n2282 = ~n2280 & ~n2281;
  assign n2283 = n2282 ^ n2277;
  assign n2284 = n2283 ^ n2277;
  assign n2285 = n2277 ^ x74;
  assign n2286 = n2285 ^ n2277;
  assign n2287 = n2284 & n2286;
  assign n2288 = n2287 ^ n2277;
  assign n2289 = n2279 & ~n2288;
  assign n2290 = n2289 ^ n2278;
  assign n2291 = n2281 ^ n2280;
  assign n2292 = ~n2277 & ~n2278;
  assign n2293 = n2292 ^ n2281;
  assign n2294 = n2293 ^ n2281;
  assign n2295 = n2281 ^ x74;
  assign n2296 = n2295 ^ n2281;
  assign n2297 = n2294 & ~n2296;
  assign n2298 = n2297 ^ n2281;
  assign n2299 = n2291 & ~n2298;
  assign n2300 = n2299 ^ n2280;
  assign n2301 = ~n2290 & ~n2300;
  assign n2302 = ~x73 & ~n2301;
  assign n1185 = x74 ^ x73;
  assign n2303 = n2282 & ~n2292;
  assign n2304 = n1185 & n2303;
  assign n2305 = ~n2282 & n2292;
  assign n2306 = x73 & x74;
  assign n2307 = n2278 & n2306;
  assign n2308 = x78 & n2307;
  assign n2309 = n2308 ^ n2306;
  assign n2310 = ~n2305 & n2309;
  assign n2311 = ~n2304 & ~n2310;
  assign n1184 = x76 ^ x75;
  assign n2312 = n2306 ^ x76;
  assign n2313 = n2312 ^ n2306;
  assign n2314 = ~x74 & ~x78;
  assign n2315 = n2314 ^ n2306;
  assign n2316 = ~n2313 & n2315;
  assign n2317 = n2316 ^ n2306;
  assign n2318 = ~n1184 & n2317;
  assign n2319 = ~x77 & n2318;
  assign n2320 = n2311 & ~n2319;
  assign n2321 = ~n2302 & n2320;
  assign n2233 = x69 & x70;
  assign n2232 = x71 & x72;
  assign n2234 = n2233 ^ n2232;
  assign n2235 = ~x69 & ~x70;
  assign n2236 = ~x71 & ~x72;
  assign n2237 = ~n2235 & ~n2236;
  assign n2238 = n2237 ^ n2232;
  assign n2239 = n2238 ^ n2232;
  assign n2240 = n2232 ^ x68;
  assign n2241 = n2240 ^ n2232;
  assign n2242 = n2239 & n2241;
  assign n2243 = n2242 ^ n2232;
  assign n2244 = n2234 & ~n2243;
  assign n2245 = n2244 ^ n2233;
  assign n2246 = n2236 ^ n2235;
  assign n2247 = ~n2232 & ~n2233;
  assign n2248 = n2247 ^ n2236;
  assign n2249 = n2248 ^ n2236;
  assign n2250 = n2236 ^ x68;
  assign n2251 = n2250 ^ n2236;
  assign n2252 = n2249 & ~n2251;
  assign n2253 = n2252 ^ n2236;
  assign n2254 = n2246 & ~n2253;
  assign n2255 = n2254 ^ n2235;
  assign n2256 = ~n2245 & ~n2255;
  assign n2257 = ~x67 & ~n2256;
  assign n1180 = x68 ^ x67;
  assign n2258 = n2237 & ~n2247;
  assign n2259 = n1180 & n2258;
  assign n2260 = ~n2237 & n2247;
  assign n2261 = x67 & x68;
  assign n2262 = n2233 & n2261;
  assign n2263 = x72 & n2262;
  assign n2264 = n2263 ^ n2261;
  assign n2265 = ~n2260 & n2264;
  assign n2266 = ~n2259 & ~n2265;
  assign n1179 = x70 ^ x69;
  assign n2267 = n2261 ^ x70;
  assign n2268 = n2267 ^ n2261;
  assign n2269 = ~x68 & ~x72;
  assign n2270 = n2269 ^ n2261;
  assign n2271 = ~n2268 & n2270;
  assign n2272 = n2271 ^ n2261;
  assign n2273 = ~n1179 & n2272;
  assign n2274 = ~x71 & n2273;
  assign n2275 = n2266 & ~n2274;
  assign n2276 = ~n2257 & n2275;
  assign n2322 = n2321 ^ n2276;
  assign n1177 = n1176 ^ n1171;
  assign n1186 = n1185 ^ n1184;
  assign n1183 = x78 ^ x77;
  assign n1187 = n1186 ^ n1183;
  assign n1181 = n1180 ^ n1179;
  assign n1178 = x72 ^ x71;
  assign n1182 = n1181 ^ n1178;
  assign n1188 = n1187 ^ n1182;
  assign n2172 = n1177 & n1188;
  assign n2174 = n1182 & n1187;
  assign n2175 = n2174 ^ n2173;
  assign n2176 = ~n2172 & ~n2175;
  assign n2231 = n2230 ^ n2176;
  assign n2323 = n2322 ^ n2231;
  assign n6026 = ~n2174 & ~n2322;
  assign n6027 = n2323 & ~n6026;
  assign n6028 = ~n2230 & ~n6027;
  assign n6029 = n2173 & n2230;
  assign n6030 = n2231 ^ n2174;
  assign n6031 = ~n2322 & ~n6030;
  assign n6032 = n6031 ^ n2174;
  assign n6033 = ~n6029 & ~n6032;
  assign n6034 = ~n6028 & n6033;
  assign n6660 = n6015 & ~n6034;
  assign n6661 = ~n6012 & n6660;
  assign n6662 = ~n6014 & ~n6661;
  assign n6021 = n2174 & n2322;
  assign n6022 = n2276 & n2321;
  assign n6023 = ~n6021 & ~n6022;
  assign n6019 = ~n2290 & n2311;
  assign n6018 = ~n2245 & n2266;
  assign n6020 = n6019 ^ n6018;
  assign n6024 = n6023 ^ n6020;
  assign n6016 = n6015 ^ n6014;
  assign n6017 = n6016 ^ n6012;
  assign n6025 = n6024 ^ n6017;
  assign n6035 = n6034 ^ n6025;
  assign n6663 = ~n6024 & n6035;
  assign n6664 = ~n6662 & ~n6663;
  assign n6665 = n6015 ^ n6012;
  assign n6666 = n6034 ^ n6015;
  assign n6667 = n6665 & ~n6666;
  assign n6668 = n6667 ^ n6034;
  assign n6669 = n6664 & ~n6668;
  assign n6670 = n6663 & n6668;
  assign n6671 = ~n6669 & ~n6670;
  assign n6657 = n6023 ^ n6019;
  assign n6658 = ~n6020 & n6657;
  assign n6659 = n6658 ^ n6023;
  assign n6672 = n6671 ^ n6659;
  assign n7303 = n6659 & ~n6670;
  assign n7304 = ~n6669 & ~n7303;
  assign n7305 = ~n6650 & ~n6653;
  assign n7306 = ~n6647 & n7305;
  assign n7309 = ~n7306 & ~n7308;
  assign n7310 = n7304 & n7309;
  assign n7311 = ~n6672 & ~n7310;
  assign n6009 = n6008 ^ n5993;
  assign n6036 = n6035 ^ n6009;
  assign n2508 = n2507 ^ n2395;
  assign n5982 = n2508 ^ n2323;
  assign n1166 = n1165 ^ n1154;
  assign n1189 = n1188 ^ n1177;
  assign n2171 = n1166 & n1189;
  assign n5983 = n2508 ^ n2171;
  assign n5984 = ~n5982 & ~n5983;
  assign n5985 = n5984 ^ n2323;
  assign n6642 = n6009 ^ n5985;
  assign n6643 = ~n6036 & n6642;
  assign n6644 = n6643 ^ n6035;
  assign n6654 = n6653 ^ n6650;
  assign n7312 = n6653 ^ n6647;
  assign n7313 = ~n6654 & n7312;
  assign n7314 = n7313 ^ n6647;
  assign n7315 = ~n6644 & n7314;
  assign n7316 = n7311 & ~n7315;
  assign n7510 = ~n7308 & n7316;
  assign n7319 = ~n6644 & ~n7306;
  assign n7320 = ~n7314 & ~n7319;
  assign n7511 = ~n6669 & ~n7320;
  assign n7512 = n6672 & ~n7511;
  assign n7513 = ~n7510 & ~n7512;
  assign n2511 = x995 & x996;
  assign n2510 = x993 & x994;
  assign n2512 = n2511 ^ n2510;
  assign n2513 = ~x995 & ~x996;
  assign n2514 = ~x993 & ~x994;
  assign n2515 = ~n2513 & ~n2514;
  assign n2516 = n2515 ^ n2510;
  assign n2517 = n2516 ^ n2510;
  assign n2518 = n2510 ^ x992;
  assign n2519 = n2518 ^ n2510;
  assign n2520 = n2517 & n2519;
  assign n2521 = n2520 ^ n2510;
  assign n2522 = n2512 & ~n2521;
  assign n2523 = n2522 ^ n2511;
  assign n1193 = x992 ^ x991;
  assign n2525 = ~n2510 & ~n2511;
  assign n2536 = n2515 & ~n2525;
  assign n2537 = n1193 & n2536;
  assign n2538 = ~n2515 & n2525;
  assign n2539 = x991 & x992;
  assign n2540 = n2510 & n2539;
  assign n2541 = x996 & n2540;
  assign n2542 = n2541 ^ n2539;
  assign n2543 = ~n2538 & n2542;
  assign n2544 = ~n2537 & ~n2543;
  assign n6042 = ~n2523 & n2544;
  assign n1196 = x5 ^ x4;
  assign n1197 = n1196 ^ x3;
  assign n1198 = x2 ^ x1;
  assign n1199 = n1198 ^ x0;
  assign n2560 = n1197 & n1199;
  assign n2570 = x1 ^ x0;
  assign n2571 = ~n1198 & n2570;
  assign n2572 = n2571 ^ x0;
  assign n2567 = x4 ^ x3;
  assign n2568 = ~n1196 & n2567;
  assign n2569 = n2568 ^ x3;
  assign n2573 = n2572 ^ n2569;
  assign n6043 = n2560 & n2573;
  assign n6044 = n2569 & n2572;
  assign n6045 = ~n6043 & ~n6044;
  assign n6631 = ~n6042 & ~n6045;
  assign n1201 = x999 ^ x998;
  assign n2564 = x998 ^ x997;
  assign n2565 = ~n1201 & n2564;
  assign n2566 = n2565 ^ x997;
  assign n2574 = n2573 ^ n2566;
  assign n1202 = n1201 ^ x997;
  assign n2556 = x6 & n1202;
  assign n1200 = n1199 ^ n1197;
  assign n1203 = n1202 ^ x6;
  assign n2557 = n1203 ^ n1199;
  assign n2558 = ~n1200 & n2557;
  assign n2559 = n2558 ^ n1203;
  assign n2561 = n2560 ^ n2559;
  assign n2562 = ~n2556 & ~n2561;
  assign n2563 = n2562 ^ n2560;
  assign n2575 = n2574 ^ n2563;
  assign n6050 = ~n2566 & ~n2575;
  assign n6051 = ~n2561 & ~n2573;
  assign n6052 = n6051 ^ n2560;
  assign n6053 = ~n2556 & n6052;
  assign n6054 = ~n6050 & ~n6053;
  assign n1192 = x994 ^ x993;
  assign n1194 = n1193 ^ n1192;
  assign n1191 = x996 ^ x995;
  assign n1195 = n1194 ^ n1191;
  assign n1204 = n1203 ^ n1200;
  assign n2555 = n1195 & n1204;
  assign n2576 = n2575 ^ n2555;
  assign n2524 = n2514 ^ n2513;
  assign n2526 = n2525 ^ n2514;
  assign n2527 = n2526 ^ n2514;
  assign n2528 = n2514 ^ x992;
  assign n2529 = n2528 ^ n2514;
  assign n2530 = n2527 & ~n2529;
  assign n2531 = n2530 ^ n2514;
  assign n2532 = n2524 & ~n2531;
  assign n2533 = n2532 ^ n2513;
  assign n2534 = ~n2523 & ~n2533;
  assign n2535 = ~x991 & ~n2534;
  assign n2545 = n2539 ^ x994;
  assign n2546 = n2545 ^ n2539;
  assign n2547 = ~x992 & ~x996;
  assign n2548 = n2547 ^ n2539;
  assign n2549 = ~n2546 & n2548;
  assign n2550 = n2549 ^ n2539;
  assign n2551 = ~n1192 & n2550;
  assign n2552 = ~x995 & n2551;
  assign n2553 = n2544 & ~n2552;
  assign n2554 = ~n2535 & n2553;
  assign n6047 = n2555 ^ n2554;
  assign n6048 = ~n2576 & ~n6047;
  assign n6049 = n6048 ^ n2575;
  assign n6055 = n6054 ^ n6049;
  assign n6046 = n6045 ^ n6042;
  assign n6633 = n6054 ^ n6046;
  assign n6634 = ~n6055 & n6633;
  assign n6635 = n6634 ^ n6054;
  assign n6636 = ~n6631 & ~n6635;
  assign n2583 = ~x11 & ~x12;
  assign n2584 = x8 & ~n2583;
  assign n2585 = ~x9 & ~x10;
  assign n2590 = n2584 & ~n2585;
  assign n2589 = x9 & x10;
  assign n2591 = n2590 ^ n2589;
  assign n2586 = x11 & x12;
  assign n2592 = n2589 ^ n2586;
  assign n2593 = n2591 & ~n2592;
  assign n2594 = n2593 ^ n2590;
  assign n2597 = ~n2586 & ~n2589;
  assign n2598 = ~n2583 & ~n2585;
  assign n2599 = n2598 ^ x8;
  assign n2600 = n2599 ^ n2598;
  assign n2601 = n2600 ^ x7;
  assign n2602 = x12 ^ x9;
  assign n2603 = x12 & n2602;
  assign n2604 = n2603 ^ n2598;
  assign n2605 = n2604 ^ x12;
  assign n2606 = n2601 & ~n2605;
  assign n2607 = n2606 ^ n2603;
  assign n2608 = n2607 ^ x12;
  assign n2609 = x7 & n2608;
  assign n2610 = n2609 ^ x7;
  assign n2611 = ~n2597 & n2610;
  assign n1213 = x10 ^ x9;
  assign n2612 = x7 & n1213;
  assign n2613 = n2584 & n2612;
  assign n2614 = ~n2611 & ~n2613;
  assign n6082 = ~n2594 & n2614;
  assign n2626 = ~x15 & ~x16;
  assign n2627 = x17 & x18;
  assign n2628 = ~n2626 & n2627;
  assign n2629 = x15 & x16;
  assign n2630 = ~n2628 & ~n2629;
  assign n2631 = ~x17 & ~x18;
  assign n2632 = x13 & ~n2631;
  assign n2633 = ~n2630 & n2632;
  assign n2634 = x13 & x14;
  assign n2635 = ~n2633 & ~n2634;
  assign n2636 = n2629 ^ x18;
  assign n2638 = n2636 ^ n2626;
  assign n2637 = n2636 ^ x17;
  assign n2639 = n2638 ^ n2637;
  assign n2640 = n2636 ^ n2629;
  assign n2641 = n2640 ^ n2636;
  assign n2642 = n2641 ^ n2638;
  assign n2643 = ~n2638 & n2642;
  assign n2644 = n2643 ^ n2638;
  assign n2645 = ~n2639 & ~n2644;
  assign n2646 = n2645 ^ n2643;
  assign n2647 = n2646 ^ n2636;
  assign n2648 = n2647 ^ n2638;
  assign n2649 = x14 & n2648;
  assign n2650 = ~n2635 & ~n2649;
  assign n2651 = x14 & ~n2631;
  assign n2652 = n2651 ^ n2629;
  assign n2653 = n2651 ^ n2628;
  assign n2654 = n2653 ^ n2628;
  assign n2655 = n2628 ^ n2627;
  assign n2656 = ~n2654 & ~n2655;
  assign n2657 = n2656 ^ n2628;
  assign n2658 = n2652 & n2657;
  assign n2659 = n2658 ^ n2629;
  assign n6081 = ~n2650 & ~n2659;
  assign n6083 = n6082 ^ n6081;
  assign n2660 = n2626 & ~n2627;
  assign n2661 = n2660 ^ n2631;
  assign n2662 = n2660 ^ n2629;
  assign n2663 = n2631 ^ x14;
  assign n2664 = n2663 ^ n2660;
  assign n2665 = ~n2660 & ~n2664;
  assign n2666 = n2665 ^ n2660;
  assign n2667 = ~n2662 & ~n2666;
  assign n2668 = n2667 ^ n2665;
  assign n2669 = n2668 ^ n2660;
  assign n2670 = n2669 ^ n2663;
  assign n2671 = n2661 & ~n2670;
  assign n2672 = n2671 ^ n2660;
  assign n2673 = ~n2659 & ~n2672;
  assign n2674 = ~x13 & ~n2673;
  assign n2675 = ~n2650 & ~n2674;
  assign n1208 = x16 ^ x15;
  assign n2676 = n2634 ^ x16;
  assign n2677 = n2676 ^ n2634;
  assign n2678 = ~x14 & ~x18;
  assign n2679 = n2678 ^ n2634;
  assign n2680 = ~n2677 & n2679;
  assign n2681 = n2680 ^ n2634;
  assign n2682 = ~n1208 & n2681;
  assign n2683 = ~x17 & n2682;
  assign n2684 = n2675 & ~n2683;
  assign n2587 = n2585 & ~n2586;
  assign n2588 = ~n2584 & n2587;
  assign n2595 = ~n2588 & ~n2594;
  assign n2596 = ~x7 & ~n2595;
  assign n2615 = ~x11 & ~n2612;
  assign n2616 = n2589 ^ x8;
  assign n2617 = x12 ^ x7;
  assign n2618 = n2589 ^ x7;
  assign n2619 = n2618 ^ x7;
  assign n2620 = ~n2617 & ~n2619;
  assign n2621 = n2620 ^ x7;
  assign n2622 = ~n2616 & n2621;
  assign n2623 = n2615 & n2622;
  assign n2624 = n2614 & ~n2623;
  assign n2625 = ~n2596 & n2624;
  assign n2685 = n2684 ^ n2625;
  assign n1207 = x18 ^ x17;
  assign n1209 = n1208 ^ n1207;
  assign n1206 = x14 ^ x13;
  assign n1210 = n1209 ^ n1206;
  assign n1212 = x8 ^ x7;
  assign n1214 = n1213 ^ n1212;
  assign n1211 = x12 ^ x11;
  assign n1215 = n1214 ^ n1211;
  assign n6057 = n1210 & n1215;
  assign n6078 = n6057 ^ n2684;
  assign n6079 = ~n2685 & n6078;
  assign n6080 = n6079 ^ n6057;
  assign n6084 = n6083 ^ n6080;
  assign n2687 = ~x27 & ~x28;
  assign n2688 = x29 & x30;
  assign n2689 = ~n2687 & n2688;
  assign n2690 = x27 & x28;
  assign n2691 = ~n2689 & ~n2690;
  assign n2692 = ~x29 & ~x30;
  assign n2693 = x25 & ~n2692;
  assign n2694 = ~n2691 & n2693;
  assign n2695 = x25 & x26;
  assign n2696 = ~n2694 & ~n2695;
  assign n2697 = n2690 ^ x30;
  assign n2699 = n2697 ^ n2687;
  assign n2698 = n2697 ^ x29;
  assign n2700 = n2699 ^ n2698;
  assign n2701 = n2697 ^ n2690;
  assign n2702 = n2701 ^ n2697;
  assign n2703 = n2702 ^ n2699;
  assign n2704 = ~n2699 & n2703;
  assign n2705 = n2704 ^ n2699;
  assign n2706 = ~n2700 & ~n2705;
  assign n2707 = n2706 ^ n2704;
  assign n2708 = n2707 ^ n2697;
  assign n2709 = n2708 ^ n2699;
  assign n2710 = x26 & n2709;
  assign n2711 = ~n2696 & ~n2710;
  assign n2712 = x26 & ~n2692;
  assign n2713 = n2712 ^ n2690;
  assign n2714 = n2712 ^ n2689;
  assign n2715 = n2714 ^ n2689;
  assign n2716 = n2689 ^ n2688;
  assign n2717 = ~n2715 & ~n2716;
  assign n2718 = n2717 ^ n2689;
  assign n2719 = n2713 & n2718;
  assign n2720 = n2719 ^ n2690;
  assign n6075 = ~n2711 & ~n2720;
  assign n2747 = x23 & x24;
  assign n2746 = x21 & x22;
  assign n2748 = n2747 ^ n2746;
  assign n2749 = ~x23 & ~x24;
  assign n2750 = ~x21 & ~x22;
  assign n2751 = ~n2749 & ~n2750;
  assign n2752 = n2751 ^ n2746;
  assign n2753 = n2752 ^ n2746;
  assign n2754 = n2746 ^ x20;
  assign n2755 = n2754 ^ n2746;
  assign n2756 = n2753 & n2755;
  assign n2757 = n2756 ^ n2746;
  assign n2758 = n2748 & ~n2757;
  assign n2759 = n2758 ^ n2747;
  assign n2761 = ~n2746 & ~n2747;
  assign n2772 = n2751 & ~n2761;
  assign n2773 = ~x20 & ~n2772;
  assign n2774 = ~n2751 & n2761;
  assign n2775 = x19 & ~n2774;
  assign n2776 = ~n2773 & n2775;
  assign n6074 = ~n2759 & ~n2776;
  assign n6076 = n6075 ^ n6074;
  assign n2760 = n2750 ^ n2749;
  assign n2762 = n2761 ^ n2750;
  assign n2763 = n2762 ^ n2750;
  assign n2764 = n2750 ^ x20;
  assign n2765 = n2764 ^ n2750;
  assign n2766 = n2763 & ~n2765;
  assign n2767 = n2766 ^ n2750;
  assign n2768 = n2760 & ~n2767;
  assign n2769 = n2768 ^ n2749;
  assign n2770 = ~n2759 & ~n2769;
  assign n2771 = ~x19 & ~n2770;
  assign n2777 = x20 & x24;
  assign n2778 = n2746 & n2777;
  assign n2779 = n2776 & ~n2778;
  assign n2780 = x24 ^ x20;
  assign n2781 = n2746 ^ x24;
  assign n2782 = n2781 ^ n2746;
  assign n2783 = n2750 ^ n2746;
  assign n2784 = ~n2782 & n2783;
  assign n2785 = n2784 ^ n2746;
  assign n2786 = ~n2780 & n2785;
  assign n2787 = ~x23 & n2786;
  assign n2788 = ~n2779 & ~n2787;
  assign n2789 = ~n2771 & n2788;
  assign n2721 = n2687 & ~n2688;
  assign n2722 = n2721 ^ n2692;
  assign n2723 = n2721 ^ n2690;
  assign n2724 = n2692 ^ x26;
  assign n2725 = n2724 ^ n2721;
  assign n2726 = ~n2721 & ~n2725;
  assign n2727 = n2726 ^ n2721;
  assign n2728 = ~n2723 & ~n2727;
  assign n2729 = n2728 ^ n2726;
  assign n2730 = n2729 ^ n2721;
  assign n2731 = n2730 ^ n2724;
  assign n2732 = n2722 & ~n2731;
  assign n2733 = n2732 ^ n2721;
  assign n2734 = ~n2720 & ~n2733;
  assign n2735 = ~x25 & ~n2734;
  assign n2736 = ~n2711 & ~n2735;
  assign n1224 = x28 ^ x27;
  assign n2737 = n2695 ^ x28;
  assign n2738 = n2737 ^ n2695;
  assign n2739 = ~x26 & ~x30;
  assign n2740 = n2739 ^ n2695;
  assign n2741 = ~n2738 & n2740;
  assign n2742 = n2741 ^ n2695;
  assign n2743 = ~n1224 & n2742;
  assign n2744 = ~x29 & n2743;
  assign n2745 = n2736 & ~n2744;
  assign n2790 = n2789 ^ n2745;
  assign n1219 = x22 ^ x21;
  assign n1218 = x20 ^ x19;
  assign n1220 = n1219 ^ n1218;
  assign n1217 = x24 ^ x23;
  assign n1221 = n1220 ^ n1217;
  assign n1223 = x30 ^ x29;
  assign n1225 = n1224 ^ n1223;
  assign n1222 = x26 ^ x25;
  assign n1226 = n1225 ^ n1222;
  assign n2686 = n1221 & n1226;
  assign n6071 = n2745 ^ n2686;
  assign n6072 = n2790 & ~n6071;
  assign n6073 = n6072 ^ n2789;
  assign n6077 = n6076 ^ n6073;
  assign n6085 = n6084 ^ n6077;
  assign n6058 = n2685 & ~n6057;
  assign n1216 = n1215 ^ n1210;
  assign n1227 = n1226 ^ n1221;
  assign n2578 = n1227 ^ n1215;
  assign n2579 = ~n1216 & n2578;
  assign n2580 = n2579 ^ n1227;
  assign n6059 = n6058 ^ n2580;
  assign n6060 = n6058 ^ n2685;
  assign n2791 = n2790 ^ n2686;
  assign n6061 = n2791 ^ n2580;
  assign n6062 = n6061 ^ n6058;
  assign n6063 = ~n6058 & n6062;
  assign n6064 = n6063 ^ n6058;
  assign n6065 = ~n6060 & ~n6064;
  assign n6066 = n6065 ^ n6063;
  assign n6067 = n6066 ^ n6058;
  assign n6068 = n6067 ^ n6061;
  assign n6069 = n6059 & n6068;
  assign n6070 = n6069 ^ n6058;
  assign n6086 = n6085 ^ n6070;
  assign n6056 = n6055 ^ n6046;
  assign n6087 = n6086 ^ n6056;
  assign n2792 = n2791 ^ n2685;
  assign n1205 = n1204 ^ n1195;
  assign n1228 = n1227 ^ n1216;
  assign n2581 = n1205 & n1228;
  assign n2582 = n2581 ^ n2580;
  assign n2793 = n2792 ^ n2582;
  assign n2577 = n2576 ^ n2554;
  assign n6039 = n2581 ^ n2577;
  assign n6040 = n2793 & ~n6039;
  assign n6041 = n6040 ^ n2581;
  assign n6617 = n6056 ^ n6041;
  assign n6618 = ~n6087 & n6617;
  assign n6619 = n6618 ^ n6086;
  assign n6630 = ~n6049 & n6054;
  assign n6632 = n6630 & n6631;
  assign n7274 = ~n6619 & ~n6632;
  assign n6626 = n6075 ^ n6073;
  assign n6627 = ~n6076 & ~n6626;
  assign n6628 = n6627 ^ n6073;
  assign n7285 = n7274 ^ n6628;
  assign n6623 = n6082 ^ n6080;
  assign n6624 = ~n6083 & ~n6623;
  assign n6625 = n6624 ^ n6080;
  assign n6620 = n6084 ^ n6070;
  assign n6621 = ~n6085 & n6620;
  assign n6622 = n6621 ^ n6070;
  assign n7283 = n6625 ^ n6622;
  assign n7284 = n7283 ^ n7274;
  assign n7286 = n7285 ^ n7284;
  assign n6629 = n6628 ^ n6625;
  assign n7287 = n7274 ^ n6629;
  assign n7288 = n7287 ^ n7274;
  assign n7289 = ~n7283 & n7288;
  assign n7290 = n7289 ^ n7283;
  assign n7291 = n7287 & ~n7290;
  assign n7292 = n7291 ^ n7274;
  assign n7293 = ~n7286 & n7292;
  assign n7294 = n7293 ^ n7289;
  assign n7295 = n7294 ^ n7274;
  assign n7296 = n7295 ^ n7285;
  assign n7297 = ~n6636 & n7296;
  assign n7514 = n7513 ^ n7297;
  assign n7272 = ~n6628 & n6636;
  assign n6637 = ~n6632 & ~n6636;
  assign n6638 = n6637 ^ n6629;
  assign n6639 = n6638 ^ n6622;
  assign n6640 = n6639 ^ n6619;
  assign n7271 = ~n6625 & n6640;
  assign n7273 = n7272 ^ n7271;
  assign n7275 = n7274 ^ n7271;
  assign n7276 = n7275 ^ n7274;
  assign n7277 = n7274 ^ n6619;
  assign n7278 = ~n7276 & n7277;
  assign n7279 = n7278 ^ n7274;
  assign n7280 = n7273 & n7279;
  assign n7281 = n7280 ^ n7272;
  assign n7282 = ~n6622 & n7281;
  assign n7298 = ~n6619 & n7272;
  assign n7299 = ~n6625 & n7298;
  assign n7300 = ~n7297 & ~n7299;
  assign n7301 = ~n7282 & n7300;
  assign n6655 = n6654 ^ n6647;
  assign n6656 = n6655 ^ n6644;
  assign n6673 = n6672 ^ n6656;
  assign n6037 = n6036 ^ n5985;
  assign n1190 = n1189 ^ n1166;
  assign n1229 = n1228 ^ n1205;
  assign n5909 = n1190 & n1229;
  assign n2794 = n2793 ^ n2577;
  assign n5978 = n5909 ^ n2794;
  assign n2324 = n2323 ^ n2171;
  assign n2509 = n2508 ^ n2324;
  assign n5979 = n5909 ^ n2509;
  assign n5980 = ~n5978 & n5979;
  assign n5981 = n5980 ^ n2794;
  assign n6038 = n6037 ^ n5981;
  assign n6088 = n6087 ^ n6041;
  assign n6614 = n6088 ^ n5981;
  assign n6615 = ~n6038 & ~n6614;
  assign n6616 = n6615 ^ n6037;
  assign n7267 = n6673 ^ n6616;
  assign n7268 = n6673 ^ n6640;
  assign n7269 = ~n7267 & n7268;
  assign n7270 = n7269 ^ n6640;
  assign n7302 = n7301 ^ n7270;
  assign n7317 = ~n7304 & n7308;
  assign n7318 = n7316 & ~n7317;
  assign n7321 = n7320 ^ n6669;
  assign n7322 = n6672 & n7321;
  assign n7323 = ~n7318 & ~n7322;
  assign n7324 = n6644 & n7306;
  assign n7325 = ~n7304 & n7324;
  assign n7326 = ~n7323 & ~n7325;
  assign n7507 = n7326 ^ n7301;
  assign n7508 = ~n7302 & n7507;
  assign n7509 = n7508 ^ n7326;
  assign n7515 = n7514 ^ n7509;
  assign n7683 = ~n7297 & ~n7513;
  assign n7684 = ~n7515 & ~n7683;
  assign n2031 = ~x989 & ~x990;
  assign n2032 = x985 & ~n2031;
  assign n1132 = x988 ^ x987;
  assign n2033 = x989 & x990;
  assign n2034 = n2033 ^ x988;
  assign n2035 = n1132 & ~n2034;
  assign n2036 = n2035 ^ x987;
  assign n2037 = n2032 & n2036;
  assign n2038 = x985 & x986;
  assign n2039 = ~n2037 & ~n2038;
  assign n2040 = ~x987 & ~x988;
  assign n2041 = ~n2033 & n2040;
  assign n2042 = x987 & x988;
  assign n2043 = ~n2031 & ~n2042;
  assign n2044 = ~n2041 & n2043;
  assign n2045 = ~x990 & n2042;
  assign n2046 = x986 & ~n2045;
  assign n2047 = ~n2044 & n2046;
  assign n2048 = ~n2039 & ~n2047;
  assign n2049 = n2033 & n2042;
  assign n2050 = x986 & ~n2031;
  assign n2051 = ~n2049 & ~n2050;
  assign n2052 = n2036 & ~n2051;
  assign n5971 = ~n2048 & ~n2052;
  assign n1997 = ~x983 & ~x984;
  assign n1137 = x982 ^ x981;
  assign n1998 = x983 & x984;
  assign n1999 = n1998 ^ x982;
  assign n2000 = n1137 & ~n1999;
  assign n2001 = n2000 ^ x981;
  assign n2002 = ~n1997 & n2001;
  assign n2003 = ~x980 & ~n2002;
  assign n2008 = ~x981 & ~x982;
  assign n2009 = ~n1998 & n2008;
  assign n2004 = x981 & x982;
  assign n2005 = n1997 & ~n2004;
  assign n2006 = n1998 & n2004;
  assign n2007 = ~n2005 & ~n2006;
  assign n2010 = n2009 ^ n2007;
  assign n2011 = n2007 ^ x979;
  assign n2012 = n2007 & n2011;
  assign n2013 = n2012 ^ n2007;
  assign n2014 = ~n2010 & n2013;
  assign n2015 = n2014 ^ n2012;
  assign n2016 = n2015 ^ n2007;
  assign n2017 = n2016 ^ x979;
  assign n2018 = x980 & n2017;
  assign n2019 = n2018 ^ x979;
  assign n2020 = ~n2003 & n2019;
  assign n2021 = x980 & ~n1997;
  assign n2022 = ~n2006 & ~n2021;
  assign n2023 = n2001 & ~n2022;
  assign n5970 = ~n2020 & ~n2023;
  assign n5972 = n5971 ^ n5970;
  assign n2053 = n2041 & ~n2050;
  assign n2054 = ~n2052 & ~n2053;
  assign n2055 = ~x985 & ~n2054;
  assign n2056 = ~n2048 & ~n2055;
  assign n2057 = ~x986 & ~x990;
  assign n2058 = n2057 ^ n2038;
  assign n2059 = n2058 ^ n2038;
  assign n1133 = x986 ^ x985;
  assign n1134 = n1133 ^ n1132;
  assign n2060 = n2038 ^ n1134;
  assign n2061 = n2060 ^ n2038;
  assign n2062 = n2059 & n2061;
  assign n2063 = n2062 ^ n2038;
  assign n2064 = ~n2042 & n2063;
  assign n2065 = n2064 ^ n2038;
  assign n2066 = ~x989 & n2065;
  assign n2067 = n2056 & ~n2066;
  assign n2024 = n2009 & ~n2021;
  assign n2025 = ~n2023 & ~n2024;
  assign n2026 = ~x979 & ~n2025;
  assign n2027 = ~n2020 & ~n2026;
  assign n1138 = x984 ^ x983;
  assign n1139 = n1138 ^ n1137;
  assign n1136 = x980 ^ x979;
  assign n1140 = n1139 ^ n1136;
  assign n2028 = ~x980 & n2005;
  assign n2029 = n1140 & n2028;
  assign n2030 = n2027 & ~n2029;
  assign n2068 = n2067 ^ n2030;
  assign n1131 = x990 ^ x989;
  assign n1135 = n1134 ^ n1131;
  assign n2069 = n1135 & n1140;
  assign n5967 = n2069 ^ n2067;
  assign n5968 = ~n2068 & n5967;
  assign n5969 = n5968 ^ n2069;
  assign n5973 = n5972 ^ n5969;
  assign n1127 = x974 ^ x973;
  assign n1125 = x976 ^ x975;
  assign n2124 = x977 & x978;
  assign n2125 = n2124 ^ x976;
  assign n2126 = n1125 & ~n2125;
  assign n2127 = n2126 ^ x975;
  assign n2128 = n1127 & n2127;
  assign n2129 = ~x975 & ~x976;
  assign n2130 = ~n2124 & n2129;
  assign n2131 = x975 & x976;
  assign n2132 = x973 & x974;
  assign n2133 = ~n2131 & n2132;
  assign n2134 = ~n2130 & n2133;
  assign n2135 = ~n2128 & ~n2134;
  assign n2136 = ~x977 & ~x978;
  assign n2137 = ~n2135 & ~n2136;
  assign n2138 = n2131 & n2132;
  assign n2139 = ~x978 & n2138;
  assign n2140 = ~n2137 & ~n2139;
  assign n2141 = n2124 & n2131;
  assign n2142 = x974 & ~n2136;
  assign n2143 = ~n2141 & ~n2142;
  assign n2144 = n2127 & ~n2143;
  assign n5964 = n2140 & ~n2144;
  assign n2090 = x971 & x972;
  assign n2089 = x969 & x970;
  assign n2095 = n2090 ^ n2089;
  assign n2086 = ~x969 & ~x970;
  assign n2087 = ~x971 & ~x972;
  assign n2088 = ~n2086 & ~n2087;
  assign n2096 = n2090 ^ n2088;
  assign n2097 = n2096 ^ n2090;
  assign n2098 = n2090 ^ x968;
  assign n2099 = n2098 ^ n2090;
  assign n2100 = n2097 & n2099;
  assign n2101 = n2100 ^ n2090;
  assign n2102 = n2095 & ~n2101;
  assign n2103 = n2102 ^ n2089;
  assign n1120 = x968 ^ x967;
  assign n2091 = ~n2089 & ~n2090;
  assign n2106 = n2088 & ~n2091;
  assign n2107 = n1120 & n2106;
  assign n2092 = ~n2088 & n2091;
  assign n2108 = x967 & x968;
  assign n2109 = n2089 & n2108;
  assign n2110 = x972 & n2109;
  assign n2111 = n2110 ^ n2108;
  assign n2112 = ~n2092 & n2111;
  assign n2113 = ~n2107 & ~n2112;
  assign n5963 = ~n2103 & n2113;
  assign n5965 = n5964 ^ n5963;
  assign n2145 = n2136 ^ n2130;
  assign n2146 = n2136 ^ n2131;
  assign n2147 = n2130 ^ x974;
  assign n2148 = n2147 ^ n2136;
  assign n2149 = n2136 & ~n2148;
  assign n2150 = n2149 ^ n2136;
  assign n2151 = n2146 & n2150;
  assign n2152 = n2151 ^ n2149;
  assign n2153 = n2152 ^ n2136;
  assign n2154 = n2153 ^ n2147;
  assign n2155 = n2145 & ~n2154;
  assign n2156 = n2155 ^ n2130;
  assign n2157 = ~n2144 & ~n2156;
  assign n2158 = ~x973 & ~n2157;
  assign n2159 = ~x974 & ~x978;
  assign n2160 = n2129 & n2159;
  assign n2161 = ~n2138 & ~n2160;
  assign n2162 = ~x977 & ~n2161;
  assign n2163 = ~n2158 & ~n2162;
  assign n2164 = n2140 & n2163;
  assign n1122 = x970 ^ x969;
  assign n1121 = x972 ^ x971;
  assign n1123 = n1122 ^ n1121;
  assign n2093 = x968 & n1123;
  assign n2094 = n2092 & ~n2093;
  assign n2104 = ~n2094 & ~n2103;
  assign n2105 = ~x967 & ~n2104;
  assign n2114 = n2108 ^ x970;
  assign n2115 = n2114 ^ n2108;
  assign n2116 = ~x968 & ~x972;
  assign n2117 = n2116 ^ n2108;
  assign n2118 = ~n2115 & n2117;
  assign n2119 = n2118 ^ n2108;
  assign n2120 = ~n1122 & n2119;
  assign n2121 = ~x971 & n2120;
  assign n2122 = n2113 & ~n2121;
  assign n2123 = ~n2105 & n2122;
  assign n2165 = n2164 ^ n2123;
  assign n1124 = n1123 ^ n1120;
  assign n1126 = x978 ^ x977;
  assign n1128 = n1127 ^ n1126;
  assign n1129 = n1128 ^ n1125;
  assign n2070 = n1124 & n1129;
  assign n5960 = n2123 ^ n2070;
  assign n5961 = n2165 & ~n5960;
  assign n5962 = n5961 ^ n2164;
  assign n5966 = n5965 ^ n5962;
  assign n5974 = n5973 ^ n5966;
  assign n5953 = n2070 & n2165;
  assign n2071 = n2069 & n2070;
  assign n1130 = n1129 ^ n1124;
  assign n2072 = n1140 ^ n1130;
  assign n1141 = n1140 ^ n1135;
  assign n2073 = n2072 ^ n1141;
  assign n2074 = n1135 ^ n1129;
  assign n2075 = n2074 ^ n1140;
  assign n2076 = n2075 ^ n1140;
  assign n2077 = ~n1130 & n2076;
  assign n2078 = n2077 ^ n1130;
  assign n2079 = n2075 & ~n2078;
  assign n2080 = n2079 ^ n1140;
  assign n2081 = n2073 & n2080;
  assign n2082 = n2081 ^ n2077;
  assign n2083 = n2082 ^ n1140;
  assign n2084 = n2083 ^ n1141;
  assign n2085 = ~n2071 & n2084;
  assign n2166 = n2165 ^ n2085;
  assign n5954 = ~n2068 & n2166;
  assign n5955 = n2068 & n2069;
  assign n5956 = ~n2084 & ~n2165;
  assign n5957 = ~n5955 & ~n5956;
  assign n5958 = ~n5954 & n5957;
  assign n5959 = ~n5953 & n5958;
  assign n5975 = n5974 ^ n5959;
  assign n6702 = n5963 & n5964;
  assign n6703 = ~n5962 & n6702;
  assign n6704 = n5975 & n6703;
  assign n6705 = n5964 ^ n5962;
  assign n6706 = ~n5965 & ~n6705;
  assign n6707 = n6706 ^ n5962;
  assign n6708 = n6707 ^ n5973;
  assign n6709 = n6707 ^ n5959;
  assign n6710 = n6709 ^ n5959;
  assign n6711 = n5975 ^ n5959;
  assign n6712 = n6710 & n6711;
  assign n6713 = n6712 ^ n5959;
  assign n6714 = ~n6708 & ~n6713;
  assign n6715 = ~n6704 & ~n6714;
  assign n6699 = n5971 ^ n5969;
  assign n6700 = ~n5972 & ~n6699;
  assign n6701 = n6700 ^ n5969;
  assign n6716 = n6715 ^ n6701;
  assign n7258 = ~n5963 & ~n5964;
  assign n7259 = n6716 & ~n7258;
  assign n7260 = n5973 & n6707;
  assign n7261 = ~n5975 & n7260;
  assign n7262 = ~n6701 & ~n7261;
  assign n7263 = ~n7259 & ~n7262;
  assign n1856 = x951 & x952;
  assign n1855 = x953 & x954;
  assign n1857 = n1856 ^ n1855;
  assign n1858 = ~x951 & ~x952;
  assign n1859 = ~x953 & ~x954;
  assign n1860 = ~n1858 & ~n1859;
  assign n1861 = n1860 ^ n1855;
  assign n1862 = n1861 ^ n1855;
  assign n1863 = n1855 ^ x950;
  assign n1864 = n1863 ^ n1855;
  assign n1865 = n1862 & n1864;
  assign n1866 = n1865 ^ n1855;
  assign n1867 = n1857 & ~n1866;
  assign n1868 = n1867 ^ n1856;
  assign n1875 = ~n1855 & ~n1856;
  assign n1876 = ~n1860 & n1875;
  assign n1877 = x949 & x950;
  assign n1878 = n1856 & n1877;
  assign n1879 = x954 & n1878;
  assign n1880 = n1879 ^ n1877;
  assign n1881 = ~n1876 & n1880;
  assign n1110 = x950 ^ x949;
  assign n1882 = n1860 & ~n1875;
  assign n1883 = n1110 & n1882;
  assign n1884 = ~n1881 & ~n1883;
  assign n5928 = ~n1868 & n1884;
  assign n1814 = x945 & x946;
  assign n1813 = x947 & x948;
  assign n1815 = n1814 ^ n1813;
  assign n1816 = ~x945 & ~x946;
  assign n1817 = ~x947 & ~x948;
  assign n1818 = ~n1816 & ~n1817;
  assign n1819 = n1818 ^ n1813;
  assign n1820 = n1819 ^ n1813;
  assign n1821 = n1813 ^ x944;
  assign n1822 = n1821 ^ n1813;
  assign n1823 = n1820 & n1822;
  assign n1824 = n1823 ^ n1813;
  assign n1825 = n1815 & ~n1824;
  assign n1826 = n1825 ^ n1814;
  assign n1833 = ~n1813 & ~n1814;
  assign n1834 = ~n1818 & n1833;
  assign n1835 = x943 & x944;
  assign n1836 = n1814 & n1835;
  assign n1837 = x948 & n1836;
  assign n1838 = n1837 ^ n1835;
  assign n1839 = ~n1834 & n1838;
  assign n1115 = x944 ^ x943;
  assign n1840 = n1818 & ~n1833;
  assign n1841 = n1115 & n1840;
  assign n1842 = ~n1839 & ~n1841;
  assign n5929 = ~n1826 & n1842;
  assign n6689 = ~n5928 & ~n5929;
  assign n1957 = ~x957 & ~x958;
  assign n1960 = x957 & x958;
  assign n1956 = x959 & x960;
  assign n1961 = n1960 ^ n1956;
  assign n1954 = ~x959 & ~x960;
  assign n1955 = x956 & ~n1954;
  assign n1962 = n1960 ^ n1955;
  assign n1963 = n1961 & n1962;
  assign n1964 = n1963 ^ n1960;
  assign n1965 = ~n1957 & n1964;
  assign n1968 = ~n1956 & ~n1960;
  assign n1969 = ~n1957 & ~n1968;
  assign n1970 = x955 & ~n1954;
  assign n1971 = n1969 & n1970;
  assign n1972 = x955 & x956;
  assign n1973 = ~n1971 & ~n1972;
  assign n1958 = ~n1956 & n1957;
  assign n1974 = ~n1954 & ~n1960;
  assign n1975 = ~n1958 & n1974;
  assign n1976 = ~x960 & n1960;
  assign n1977 = x956 & ~n1976;
  assign n1978 = ~n1975 & n1977;
  assign n1979 = ~n1973 & ~n1978;
  assign n5939 = ~n1965 & ~n1979;
  assign n1918 = ~x963 & ~x964;
  assign n1921 = x963 & x964;
  assign n1917 = x965 & x966;
  assign n1922 = n1921 ^ n1917;
  assign n1915 = ~x965 & ~x966;
  assign n1916 = x962 & ~n1915;
  assign n1923 = n1921 ^ n1916;
  assign n1924 = n1922 & n1923;
  assign n1925 = n1924 ^ n1921;
  assign n1926 = ~n1918 & n1925;
  assign n1929 = ~n1917 & ~n1921;
  assign n1930 = ~n1918 & ~n1929;
  assign n1931 = x961 & ~n1915;
  assign n1932 = n1930 & n1931;
  assign n1933 = x961 & x962;
  assign n1934 = ~n1932 & ~n1933;
  assign n1919 = ~n1917 & n1918;
  assign n1935 = ~n1915 & ~n1921;
  assign n1936 = ~n1919 & n1935;
  assign n1937 = ~x966 & n1921;
  assign n1938 = x962 & ~n1937;
  assign n1939 = ~n1936 & n1938;
  assign n1940 = ~n1934 & ~n1939;
  assign n5938 = ~n1926 & ~n1940;
  assign n5940 = n5939 ^ n5938;
  assign n1959 = ~n1955 & n1958;
  assign n1966 = ~n1959 & ~n1965;
  assign n1967 = ~x955 & ~n1966;
  assign n1980 = ~n1967 & ~n1979;
  assign n1981 = ~x956 & ~x960;
  assign n1982 = n1981 ^ n1972;
  assign n1983 = n1982 ^ n1972;
  assign n1984 = x955 & ~n1957;
  assign n1985 = n1984 ^ n1972;
  assign n1986 = n1985 ^ n1972;
  assign n1987 = n1983 & ~n1986;
  assign n1988 = n1987 ^ n1972;
  assign n1989 = ~n1960 & n1988;
  assign n1990 = n1989 ^ n1972;
  assign n1991 = ~x959 & n1990;
  assign n1992 = n1980 & ~n1991;
  assign n1920 = ~n1916 & n1919;
  assign n1927 = ~n1920 & ~n1926;
  assign n1928 = ~x961 & ~n1927;
  assign n1941 = ~n1928 & ~n1940;
  assign n1942 = ~x962 & ~x966;
  assign n1943 = n1942 ^ n1933;
  assign n1944 = n1943 ^ n1933;
  assign n1945 = x961 & ~n1918;
  assign n1946 = n1945 ^ n1933;
  assign n1947 = n1946 ^ n1933;
  assign n1948 = n1944 & ~n1947;
  assign n1949 = n1948 ^ n1933;
  assign n1950 = ~n1921 & n1949;
  assign n1951 = n1950 ^ n1933;
  assign n1952 = ~x965 & n1951;
  assign n1953 = n1941 & ~n1952;
  assign n1993 = n1992 ^ n1953;
  assign n1099 = x960 ^ x959;
  assign n1098 = x958 ^ x957;
  assign n1100 = n1099 ^ n1098;
  assign n1097 = x956 ^ x955;
  assign n1101 = n1100 ^ n1097;
  assign n1104 = x966 ^ x965;
  assign n1103 = x964 ^ x963;
  assign n1105 = n1104 ^ n1103;
  assign n1102 = x962 ^ x961;
  assign n1106 = n1105 ^ n1102;
  assign n1898 = n1101 & n1106;
  assign n5935 = n1953 ^ n1898;
  assign n5936 = n1993 & ~n5935;
  assign n5937 = n5936 ^ n1992;
  assign n5941 = n5940 ^ n5937;
  assign n1108 = x954 ^ x953;
  assign n1869 = x953 ^ x950;
  assign n1870 = n1108 & n1869;
  assign n1871 = n1870 ^ x953;
  assign n1872 = n1858 & ~n1871;
  assign n1873 = ~n1868 & ~n1872;
  assign n1874 = ~x949 & ~n1873;
  assign n1885 = ~x950 & ~x954;
  assign n1886 = n1885 ^ n1877;
  assign n1887 = n1886 ^ n1877;
  assign n1109 = x952 ^ x951;
  assign n1111 = n1110 ^ n1109;
  assign n1888 = n1877 ^ n1111;
  assign n1889 = n1888 ^ n1877;
  assign n1890 = n1887 & n1889;
  assign n1891 = n1890 ^ n1877;
  assign n1892 = ~n1856 & n1891;
  assign n1893 = n1892 ^ n1877;
  assign n1894 = ~x953 & n1893;
  assign n1895 = n1884 & ~n1894;
  assign n1896 = ~n1874 & n1895;
  assign n1113 = x948 ^ x947;
  assign n1827 = x947 ^ x944;
  assign n1828 = n1113 & n1827;
  assign n1829 = n1828 ^ x947;
  assign n1830 = n1816 & ~n1829;
  assign n1831 = ~n1826 & ~n1830;
  assign n1832 = ~x943 & ~n1831;
  assign n1843 = ~x944 & ~x948;
  assign n1844 = n1843 ^ n1835;
  assign n1845 = n1844 ^ n1835;
  assign n1114 = x946 ^ x945;
  assign n1116 = n1115 ^ n1114;
  assign n1846 = n1835 ^ n1116;
  assign n1847 = n1846 ^ n1835;
  assign n1848 = n1845 & n1847;
  assign n1849 = n1848 ^ n1835;
  assign n1850 = ~n1814 & n1849;
  assign n1851 = n1850 ^ n1835;
  assign n1852 = ~x947 & n1851;
  assign n1853 = n1842 & ~n1852;
  assign n1854 = ~n1832 & n1853;
  assign n1897 = n1896 ^ n1854;
  assign n1112 = n1111 ^ n1108;
  assign n1117 = n1116 ^ n1113;
  assign n1899 = n1112 & n1117;
  assign n5931 = n1897 & n1899;
  assign n5932 = n1854 & n1896;
  assign n5933 = ~n5931 & ~n5932;
  assign n5943 = n1898 & n1993;
  assign n1107 = n1106 ^ n1101;
  assign n1901 = n1117 ^ n1107;
  assign n1118 = n1117 ^ n1112;
  assign n1902 = n1901 ^ n1118;
  assign n1903 = n1112 ^ n1106;
  assign n1904 = n1903 ^ n1117;
  assign n1905 = n1904 ^ n1117;
  assign n1906 = ~n1107 & n1905;
  assign n1907 = n1906 ^ n1107;
  assign n1908 = n1904 & ~n1907;
  assign n1909 = n1908 ^ n1117;
  assign n1910 = n1902 & n1909;
  assign n1911 = n1910 ^ n1906;
  assign n1912 = n1911 ^ n1117;
  assign n1913 = n1912 ^ n1118;
  assign n5944 = ~n1913 & ~n1993;
  assign n1900 = n1898 & n1899;
  assign n1914 = ~n1900 & n1913;
  assign n1994 = n1993 ^ n1914;
  assign n1995 = n1994 ^ n1897;
  assign n5945 = n1995 ^ n1994;
  assign n5946 = n1994 ^ n1899;
  assign n5947 = n5945 & n5946;
  assign n5948 = n5947 ^ n1994;
  assign n5949 = ~n5944 & ~n5948;
  assign n5950 = ~n5943 & n5949;
  assign n6679 = n5933 & ~n5950;
  assign n6680 = n5941 & ~n6679;
  assign n6681 = ~n5933 & n5950;
  assign n6682 = ~n6680 & ~n6681;
  assign n6683 = n5928 & n5929;
  assign n6684 = n6682 & n6683;
  assign n6685 = n6679 ^ n5941;
  assign n5930 = n5929 ^ n5928;
  assign n5934 = n5933 ^ n5930;
  assign n5942 = n5941 ^ n5934;
  assign n5951 = n5950 ^ n5942;
  assign n6686 = n5951 & ~n6683;
  assign n6687 = n6686 ^ n6679;
  assign n6688 = n6687 ^ n6686;
  assign n6690 = n6689 ^ n6686;
  assign n6691 = n6688 & ~n6690;
  assign n6692 = n6691 ^ n6686;
  assign n6693 = n6685 & n6692;
  assign n6694 = ~n6684 & ~n6693;
  assign n6676 = n5939 ^ n5937;
  assign n6677 = ~n5940 & ~n6676;
  assign n6678 = n6677 ^ n5937;
  assign n6695 = n6694 ^ n6678;
  assign n7255 = ~n6689 & n6695;
  assign n7256 = ~n6678 & n6682;
  assign n7257 = ~n7255 & ~n7256;
  assign n7264 = n7263 ^ n7257;
  assign n2167 = n2166 ^ n2068;
  assign n1119 = n1118 ^ n1107;
  assign n1142 = n1141 ^ n1130;
  assign n1996 = n1119 & n1142;
  assign n2168 = n2167 ^ n1996;
  assign n5925 = n1996 ^ n1995;
  assign n5926 = n2168 & ~n5925;
  assign n5927 = n5926 ^ n2167;
  assign n5952 = n5951 ^ n5927;
  assign n6696 = n5975 ^ n5951;
  assign n6697 = n5952 & ~n6696;
  assign n6698 = n6697 ^ n5975;
  assign n6717 = n6716 ^ n6698;
  assign n7252 = n6698 ^ n6695;
  assign n7253 = n6717 & ~n7252;
  assign n7254 = n7253 ^ n6716;
  assign n7516 = n7257 ^ n7254;
  assign n7517 = n7264 & ~n7516;
  assign n7518 = n7517 ^ n7263;
  assign n7265 = n7264 ^ n7254;
  assign n6641 = n6640 ^ n6616;
  assign n6674 = n6673 ^ n6641;
  assign n5976 = n5975 ^ n5952;
  assign n2169 = n2168 ^ n1995;
  assign n5913 = n5909 ^ n2169;
  assign n2795 = n2794 ^ n2509;
  assign n5910 = n5909 ^ n2795;
  assign n1230 = n1229 ^ n1190;
  assign n1143 = n1142 ^ n1119;
  assign n1810 = n1190 ^ n1143;
  assign n1811 = n1230 & ~n1810;
  assign n1812 = n1811 ^ n1229;
  assign n5911 = n5910 ^ n1812;
  assign n5912 = n5911 ^ n5909;
  assign n5914 = n5913 ^ n5912;
  assign n2170 = n2169 ^ n1812;
  assign n5915 = n5909 ^ n2170;
  assign n5916 = n5915 ^ n5909;
  assign n5917 = ~n5911 & n5916;
  assign n5918 = n5917 ^ n5911;
  assign n5919 = n5915 & ~n5918;
  assign n5920 = n5919 ^ n5909;
  assign n5921 = ~n5914 & n5920;
  assign n5922 = n5921 ^ n5917;
  assign n5923 = n5922 ^ n5909;
  assign n5924 = n5923 ^ n5913;
  assign n5977 = n5976 ^ n5924;
  assign n6089 = n6088 ^ n6038;
  assign n6611 = n6089 ^ n5924;
  assign n6612 = n5977 & n6611;
  assign n6613 = n6612 ^ n6089;
  assign n6675 = n6674 ^ n6613;
  assign n6718 = n6717 ^ n6695;
  assign n7249 = n6718 ^ n6613;
  assign n7250 = n6675 & ~n7249;
  assign n7251 = n7250 ^ n6674;
  assign n7266 = n7265 ^ n7251;
  assign n7327 = n7326 ^ n7302;
  assign n7519 = n7327 ^ n7251;
  assign n7520 = ~n7266 & n7519;
  assign n7521 = n7520 ^ n7327;
  assign n7689 = n7518 & n7521;
  assign n7690 = n7684 & n7689;
  assign n7522 = n7521 ^ n7518;
  assign n7685 = n7518 ^ n7515;
  assign n7686 = n7522 & ~n7685;
  assign n7687 = n7686 ^ n7521;
  assign n7688 = ~n7684 & ~n7687;
  assign n1434 = x863 & x864;
  assign n1433 = x861 & x862;
  assign n1435 = n1434 ^ n1433;
  assign n1436 = ~x863 & ~x864;
  assign n1437 = ~x861 & ~x862;
  assign n1438 = ~n1436 & ~n1437;
  assign n1439 = n1438 ^ n1433;
  assign n1440 = n1439 ^ n1433;
  assign n1441 = n1433 ^ x860;
  assign n1442 = n1441 ^ n1433;
  assign n1443 = n1440 & n1442;
  assign n1444 = n1443 ^ n1433;
  assign n1445 = n1435 & ~n1444;
  assign n1446 = n1445 ^ n1434;
  assign n1027 = x860 ^ x859;
  assign n1448 = ~n1433 & ~n1434;
  assign n1459 = n1438 & ~n1448;
  assign n1460 = n1027 & n1459;
  assign n1461 = ~n1438 & n1448;
  assign n1462 = x859 & x860;
  assign n1463 = n1433 & n1462;
  assign n1464 = x864 & n1463;
  assign n1465 = n1464 ^ n1462;
  assign n1466 = ~n1461 & n1465;
  assign n1467 = ~n1460 & ~n1466;
  assign n5824 = ~n1446 & n1467;
  assign n1389 = x869 & x870;
  assign n1388 = x867 & x868;
  assign n1390 = n1389 ^ n1388;
  assign n1391 = ~x869 & ~x870;
  assign n1392 = ~x867 & ~x868;
  assign n1393 = ~n1391 & ~n1392;
  assign n1394 = n1393 ^ n1388;
  assign n1395 = n1394 ^ n1388;
  assign n1396 = n1388 ^ x866;
  assign n1397 = n1396 ^ n1388;
  assign n1398 = n1395 & n1397;
  assign n1399 = n1398 ^ n1388;
  assign n1400 = n1390 & ~n1399;
  assign n1401 = n1400 ^ n1389;
  assign n1032 = x866 ^ x865;
  assign n1403 = ~n1388 & ~n1389;
  assign n1414 = n1393 & ~n1403;
  assign n1415 = n1032 & n1414;
  assign n1416 = ~n1393 & n1403;
  assign n1417 = x865 & x866;
  assign n1418 = n1388 & n1417;
  assign n1419 = x870 & n1418;
  assign n1420 = n1419 ^ n1417;
  assign n1421 = ~n1416 & n1420;
  assign n1422 = ~n1415 & ~n1421;
  assign n5823 = ~n1401 & n1422;
  assign n5825 = n5824 ^ n5823;
  assign n1447 = n1437 ^ n1436;
  assign n1449 = n1448 ^ n1437;
  assign n1450 = n1449 ^ n1437;
  assign n1451 = n1437 ^ x860;
  assign n1452 = n1451 ^ n1437;
  assign n1453 = n1450 & ~n1452;
  assign n1454 = n1453 ^ n1437;
  assign n1455 = n1447 & ~n1454;
  assign n1456 = n1455 ^ n1436;
  assign n1457 = ~n1446 & ~n1456;
  assign n1458 = ~x859 & ~n1457;
  assign n1026 = x862 ^ x861;
  assign n1468 = n1462 ^ x862;
  assign n1469 = n1468 ^ n1462;
  assign n1470 = ~x860 & ~x864;
  assign n1471 = n1470 ^ n1462;
  assign n1472 = ~n1469 & n1471;
  assign n1473 = n1472 ^ n1462;
  assign n1474 = ~n1026 & n1473;
  assign n1475 = ~x863 & n1474;
  assign n1476 = n1467 & ~n1475;
  assign n1477 = ~n1458 & n1476;
  assign n1402 = n1392 ^ n1391;
  assign n1404 = n1403 ^ n1392;
  assign n1405 = n1404 ^ n1392;
  assign n1406 = n1392 ^ x866;
  assign n1407 = n1406 ^ n1392;
  assign n1408 = n1405 & ~n1407;
  assign n1409 = n1408 ^ n1392;
  assign n1410 = n1402 & ~n1409;
  assign n1411 = n1410 ^ n1391;
  assign n1412 = ~n1401 & ~n1411;
  assign n1413 = ~x865 & ~n1412;
  assign n1031 = x868 ^ x867;
  assign n1423 = n1417 ^ x868;
  assign n1424 = n1423 ^ n1417;
  assign n1425 = ~x866 & ~x870;
  assign n1426 = n1425 ^ n1417;
  assign n1427 = ~n1424 & n1426;
  assign n1428 = n1427 ^ n1417;
  assign n1429 = ~n1031 & n1428;
  assign n1430 = ~x869 & n1429;
  assign n1431 = n1422 & ~n1430;
  assign n1432 = ~n1413 & n1431;
  assign n1478 = n1477 ^ n1432;
  assign n1028 = n1027 ^ n1026;
  assign n1025 = x864 ^ x863;
  assign n1029 = n1028 ^ n1025;
  assign n1033 = n1032 ^ n1031;
  assign n1030 = x870 ^ x869;
  assign n1034 = n1033 ^ n1030;
  assign n1386 = n1029 & n1034;
  assign n5820 = n1432 ^ n1386;
  assign n5821 = n1478 & ~n5820;
  assign n5822 = n5821 ^ n1477;
  assign n5826 = n5825 ^ n5822;
  assign n1038 = x854 ^ x853;
  assign n1037 = x856 ^ x855;
  assign n1506 = x857 & x858;
  assign n1507 = n1506 ^ x856;
  assign n1508 = n1037 & ~n1507;
  assign n1509 = n1508 ^ x855;
  assign n1510 = n1038 & n1509;
  assign n1511 = ~x855 & ~x856;
  assign n1512 = ~n1506 & n1511;
  assign n1513 = x855 & x856;
  assign n1514 = x853 & x854;
  assign n1515 = ~n1513 & n1514;
  assign n1516 = ~n1512 & n1515;
  assign n1517 = ~n1510 & ~n1516;
  assign n1518 = ~x857 & ~x858;
  assign n1519 = ~n1517 & ~n1518;
  assign n1520 = n1513 & n1514;
  assign n1521 = ~x858 & n1520;
  assign n1522 = ~n1519 & ~n1521;
  assign n1523 = ~x854 & ~x858;
  assign n1524 = n1523 ^ n1514;
  assign n1525 = n1524 ^ n1514;
  assign n1039 = n1038 ^ n1037;
  assign n1526 = n1514 ^ n1039;
  assign n1527 = n1526 ^ n1514;
  assign n1528 = n1525 & n1527;
  assign n1529 = n1528 ^ n1514;
  assign n1530 = ~n1513 & n1529;
  assign n1531 = n1530 ^ n1514;
  assign n1532 = ~x857 & n1531;
  assign n1533 = n1522 & ~n1532;
  assign n1534 = x854 & ~n1518;
  assign n1535 = n1506 & n1513;
  assign n1536 = ~n1534 & ~n1535;
  assign n1537 = n1509 & ~n1536;
  assign n1538 = n1512 & ~n1534;
  assign n1539 = ~n1537 & ~n1538;
  assign n1540 = ~x853 & ~n1539;
  assign n1541 = n1533 & ~n1540;
  assign n1481 = ~x851 & ~x852;
  assign n1482 = ~x849 & ~x850;
  assign n1483 = ~n1481 & ~n1482;
  assign n1484 = x851 & x852;
  assign n1485 = x849 & x850;
  assign n1486 = ~n1484 & ~n1485;
  assign n1487 = n1483 & ~n1486;
  assign n1488 = x848 & n1487;
  assign n1489 = n1484 & n1485;
  assign n1490 = ~n1488 & ~n1489;
  assign n1491 = ~n1483 & n1486;
  assign n1492 = ~x848 & n1491;
  assign n1493 = n1490 & ~n1492;
  assign n1494 = ~x847 & ~n1493;
  assign n1043 = x848 ^ x847;
  assign n1495 = n1481 & n1482;
  assign n1496 = n1043 & n1495;
  assign n1497 = n1487 ^ x848;
  assign n1498 = n1497 ^ n1487;
  assign n1499 = ~n1489 & ~n1491;
  assign n1500 = n1499 ^ n1487;
  assign n1501 = n1498 & n1500;
  assign n1502 = n1501 ^ n1487;
  assign n1503 = x847 & n1502;
  assign n1504 = ~n1496 & ~n1503;
  assign n1505 = ~n1494 & n1504;
  assign n1542 = n1541 ^ n1505;
  assign n1036 = x858 ^ x857;
  assign n1040 = n1039 ^ n1036;
  assign n1042 = x850 ^ x849;
  assign n1044 = n1043 ^ n1042;
  assign n1041 = x852 ^ x851;
  assign n1045 = n1044 ^ n1041;
  assign n1480 = n1040 & n1045;
  assign n5828 = n1505 ^ n1480;
  assign n5829 = n1542 & ~n5828;
  assign n5830 = n5829 ^ n1541;
  assign n1543 = n1542 ^ n1480;
  assign n1035 = n1034 ^ n1029;
  assign n1046 = n1045 ^ n1040;
  assign n1385 = n1035 & n1046;
  assign n5831 = n1543 ^ n1385;
  assign n5832 = n1478 ^ n1386;
  assign n5833 = n5832 ^ n1478;
  assign n5834 = n1478 ^ n1385;
  assign n5835 = n5834 ^ n1478;
  assign n5836 = ~n5833 & ~n5835;
  assign n5837 = n5836 ^ n1478;
  assign n5838 = n5831 & n5837;
  assign n5839 = n5838 ^ n1543;
  assign n6727 = ~n5830 & ~n5839;
  assign n6728 = n5826 & ~n6727;
  assign n6729 = n5830 & n5839;
  assign n6730 = ~n6728 & ~n6729;
  assign n5818 = n1522 & ~n1537;
  assign n5817 = n1490 & ~n1503;
  assign n5819 = n5818 ^ n5817;
  assign n6731 = n6727 ^ n5817;
  assign n6732 = n6731 ^ n5817;
  assign n6733 = n5826 ^ n5817;
  assign n6734 = n6733 ^ n5817;
  assign n6735 = n6732 & ~n6734;
  assign n6736 = n6735 ^ n5817;
  assign n6737 = n5819 & ~n6736;
  assign n6738 = n6737 ^ n5818;
  assign n6739 = n6730 & n6738;
  assign n6740 = ~n5817 & ~n5818;
  assign n6741 = n6728 & n6740;
  assign n6742 = n5817 & n5818;
  assign n6743 = n5826 & ~n6742;
  assign n6744 = n6729 & n6743;
  assign n6745 = ~n6741 & ~n6744;
  assign n6746 = ~n6739 & n6745;
  assign n6724 = n5824 ^ n5822;
  assign n6725 = ~n5825 & ~n6724;
  assign n6726 = n6725 ^ n5822;
  assign n6747 = n6746 ^ n6726;
  assign n5840 = n5839 ^ n5830;
  assign n5827 = n5826 ^ n5819;
  assign n5841 = n5840 ^ n5827;
  assign n1344 = x875 & x876;
  assign n1345 = x873 & x874;
  assign n1346 = ~n1344 & ~n1345;
  assign n1347 = ~x875 & ~x876;
  assign n1348 = ~x873 & ~x874;
  assign n1349 = ~n1347 & ~n1348;
  assign n1350 = n1346 & ~n1349;
  assign n1351 = x871 & x872;
  assign n1352 = n1345 & n1351;
  assign n1353 = x876 & n1352;
  assign n1354 = n1353 ^ n1351;
  assign n1355 = ~n1350 & n1354;
  assign n1356 = n1344 & n1345;
  assign n1357 = ~n1355 & ~n1356;
  assign n1358 = ~n1346 & n1349;
  assign n1359 = ~x872 & n1358;
  assign n1360 = ~x871 & n1359;
  assign n1361 = n1360 ^ n1358;
  assign n1362 = n1357 & ~n1361;
  assign n1002 = x876 ^ x875;
  assign n1363 = x875 ^ x872;
  assign n1364 = n1002 & n1363;
  assign n1365 = n1364 ^ x875;
  assign n1366 = n1348 & ~n1365;
  assign n1367 = n1362 & ~n1366;
  assign n1368 = x871 & ~n1355;
  assign n1369 = ~n1359 & n1368;
  assign n1370 = ~n1367 & ~n1369;
  assign n1371 = ~x872 & ~x876;
  assign n1372 = n1371 ^ n1351;
  assign n1373 = n1372 ^ n1351;
  assign n1004 = x872 ^ x871;
  assign n1003 = x874 ^ x873;
  assign n1005 = n1004 ^ n1003;
  assign n1374 = n1351 ^ n1005;
  assign n1375 = n1374 ^ n1351;
  assign n1376 = n1373 & n1375;
  assign n1377 = n1376 ^ n1351;
  assign n1378 = ~n1345 & n1377;
  assign n1379 = n1378 ^ n1351;
  assign n1380 = ~x875 & n1379;
  assign n1381 = ~n1370 & ~n1380;
  assign n1319 = ~x881 & ~x882;
  assign n1320 = ~x879 & ~x880;
  assign n1321 = ~n1319 & ~n1320;
  assign n1322 = x881 & x882;
  assign n1323 = x879 & x880;
  assign n1324 = ~n1322 & ~n1323;
  assign n1325 = n1321 & ~n1324;
  assign n1326 = x878 & n1325;
  assign n1327 = n1322 & n1323;
  assign n1328 = ~n1326 & ~n1327;
  assign n1329 = ~n1321 & n1324;
  assign n1330 = ~x878 & n1329;
  assign n1331 = n1328 & ~n1330;
  assign n1332 = ~x877 & ~n1331;
  assign n1009 = x878 ^ x877;
  assign n1333 = n1319 & n1320;
  assign n1334 = n1009 & n1333;
  assign n1335 = n1325 ^ x878;
  assign n1336 = n1335 ^ n1325;
  assign n1337 = ~n1327 & ~n1329;
  assign n1338 = n1337 ^ n1325;
  assign n1339 = n1336 & n1338;
  assign n1340 = n1339 ^ n1325;
  assign n1341 = x877 & n1340;
  assign n1342 = ~n1334 & ~n1341;
  assign n1343 = ~n1332 & n1342;
  assign n1382 = n1381 ^ n1343;
  assign n1281 = x887 & x888;
  assign n1282 = x885 & x886;
  assign n1283 = n1281 & n1282;
  assign n1284 = ~n1281 & ~n1282;
  assign n1285 = ~x887 & ~x888;
  assign n1286 = ~x885 & ~x886;
  assign n1287 = ~n1285 & ~n1286;
  assign n1288 = ~n1284 & n1287;
  assign n1289 = ~x884 & n1288;
  assign n1290 = ~x883 & n1289;
  assign n1291 = n1290 ^ n1288;
  assign n1292 = ~n1283 & ~n1291;
  assign n1013 = x888 ^ x887;
  assign n1293 = x887 ^ x884;
  assign n1294 = n1013 & n1293;
  assign n1295 = n1294 ^ x887;
  assign n1296 = n1286 & ~n1295;
  assign n1297 = n1292 & ~n1296;
  assign n1298 = x883 & ~n1289;
  assign n1299 = ~n1297 & ~n1298;
  assign n1300 = x883 & x884;
  assign n1015 = x884 ^ x883;
  assign n1014 = x886 ^ x885;
  assign n1016 = n1015 ^ n1014;
  assign n1301 = n1300 ^ n1016;
  assign n1302 = n1301 ^ n1300;
  assign n1303 = ~x884 & ~x888;
  assign n1304 = n1303 ^ n1300;
  assign n1305 = n1304 ^ n1300;
  assign n1306 = n1302 & n1305;
  assign n1307 = n1306 ^ n1300;
  assign n1308 = ~n1282 & n1307;
  assign n1309 = n1308 ^ n1300;
  assign n1310 = ~x887 & n1309;
  assign n1311 = n1284 & ~n1287;
  assign n1312 = n1282 & n1300;
  assign n1313 = x888 & n1312;
  assign n1314 = n1313 ^ n1300;
  assign n1315 = ~n1311 & n1314;
  assign n1316 = ~n1310 & ~n1315;
  assign n1317 = ~n1299 & n1316;
  assign n1256 = x893 & x894;
  assign n1257 = x891 & x892;
  assign n1258 = ~n1256 & ~n1257;
  assign n1259 = ~x893 & ~x894;
  assign n1260 = ~x891 & ~x892;
  assign n1261 = ~n1259 & ~n1260;
  assign n1262 = ~n1258 & n1261;
  assign n1263 = x890 & n1262;
  assign n1264 = n1256 & n1257;
  assign n1265 = ~n1263 & ~n1264;
  assign n1266 = n1258 & ~n1261;
  assign n1267 = ~x890 & n1266;
  assign n1268 = n1265 & ~n1267;
  assign n1269 = ~x889 & ~n1268;
  assign n1020 = x890 ^ x889;
  assign n1270 = n1259 & n1260;
  assign n1271 = n1020 & n1270;
  assign n1272 = n1262 ^ x890;
  assign n1273 = n1272 ^ n1262;
  assign n1274 = ~n1264 & ~n1266;
  assign n1275 = n1274 ^ n1262;
  assign n1276 = n1273 & n1275;
  assign n1277 = n1276 ^ n1262;
  assign n1278 = x889 & n1277;
  assign n1279 = ~n1271 & ~n1278;
  assign n1280 = ~n1269 & n1279;
  assign n1318 = n1317 ^ n1280;
  assign n1383 = n1382 ^ n1318;
  assign n1017 = n1016 ^ n1013;
  assign n1019 = x892 ^ x891;
  assign n1021 = n1020 ^ n1019;
  assign n1018 = x894 ^ x893;
  assign n1022 = n1021 ^ n1018;
  assign n1235 = n1017 & n1022;
  assign n1008 = x880 ^ x879;
  assign n1010 = n1009 ^ n1008;
  assign n1007 = x882 ^ x881;
  assign n1011 = n1010 ^ n1007;
  assign n1006 = n1005 ^ n1002;
  assign n1012 = n1011 ^ n1006;
  assign n1023 = n1022 ^ n1017;
  assign n1236 = n1023 ^ n1006;
  assign n1237 = n1012 & ~n1236;
  assign n1238 = n1237 ^ n1011;
  assign n1239 = ~n1235 & ~n1238;
  assign n1024 = n1023 ^ n1012;
  assign n1047 = n1046 ^ n1035;
  assign n1240 = n1024 & n1047;
  assign n1241 = ~n1239 & n1240;
  assign n1242 = ~n1006 & ~n1011;
  assign n1243 = ~n1017 & ~n1022;
  assign n1244 = n1242 & n1243;
  assign n1245 = ~n1241 & ~n1244;
  assign n1246 = n1006 & n1011;
  assign n1247 = n1246 ^ n1047;
  assign n1248 = n1247 ^ n1246;
  assign n1249 = n1246 ^ n1238;
  assign n1250 = n1249 ^ n1246;
  assign n1251 = ~n1248 & ~n1250;
  assign n1252 = n1251 ^ n1246;
  assign n1253 = ~n1235 & n1252;
  assign n1254 = n1253 ^ n1246;
  assign n1255 = n1245 & ~n1254;
  assign n1384 = n1383 ^ n1255;
  assign n1387 = ~n1385 & ~n1386;
  assign n1479 = n1478 ^ n1387;
  assign n1544 = n1543 ^ n1479;
  assign n5814 = n1544 ^ n1240;
  assign n5815 = ~n1384 & ~n5814;
  assign n5816 = n5815 ^ n1544;
  assign n5842 = n5841 ^ n5816;
  assign n5802 = ~n1235 & ~n1318;
  assign n5803 = n5802 ^ n1246;
  assign n5804 = n5803 ^ n1246;
  assign n5805 = n1250 & ~n5804;
  assign n5806 = n5805 ^ n1246;
  assign n5807 = ~n1382 & ~n5806;
  assign n5808 = n5807 ^ n1246;
  assign n5809 = n1239 ^ n1235;
  assign n5810 = ~n1318 & n5809;
  assign n5811 = n5810 ^ n1235;
  assign n5812 = ~n5808 & ~n5811;
  assign n5797 = ~n1235 & n1318;
  assign n5798 = ~n1280 & ~n1317;
  assign n5799 = ~n5797 & ~n5798;
  assign n5794 = n1328 & ~n1341;
  assign n5795 = n5794 ^ n1362;
  assign n5792 = n1265 & ~n1278;
  assign n5791 = n1292 & ~n1315;
  assign n5793 = n5792 ^ n5791;
  assign n5796 = n5795 ^ n5793;
  assign n5800 = n5799 ^ n5796;
  assign n5788 = ~n1246 & n1382;
  assign n5789 = ~n1343 & ~n1381;
  assign n5790 = ~n5788 & ~n5789;
  assign n5801 = n5800 ^ n5790;
  assign n5813 = n5812 ^ n5801;
  assign n6721 = n5816 ^ n5813;
  assign n6722 = ~n5842 & n6721;
  assign n6723 = n6722 ^ n5841;
  assign n6748 = n6747 ^ n6723;
  assign n6750 = ~n5792 & n5799;
  assign n6751 = ~n5791 & n6750;
  assign n6749 = n1362 & n5794;
  assign n6752 = n6751 ^ n6749;
  assign n6753 = n5799 ^ n5792;
  assign n6754 = ~n5793 & ~n6753;
  assign n6755 = n6754 ^ n5799;
  assign n6756 = n6755 ^ n6749;
  assign n6757 = n5791 & n5792;
  assign n6758 = ~n5799 & n6757;
  assign n6759 = ~n1362 & ~n5794;
  assign n6760 = ~n6758 & n6759;
  assign n6761 = ~n6750 & n6760;
  assign n6762 = n6761 ^ n6755;
  assign n6763 = ~n6755 & n6762;
  assign n6764 = n6763 ^ n6755;
  assign n6765 = n6756 & ~n6764;
  assign n6766 = n6765 ^ n6763;
  assign n6767 = n6766 ^ n6755;
  assign n6768 = n6767 ^ n6761;
  assign n6769 = ~n6752 & n6768;
  assign n6770 = n6769 ^ n6761;
  assign n6771 = n6770 ^ n5790;
  assign n6772 = n6771 ^ n6770;
  assign n6773 = ~n5790 & n5794;
  assign n6774 = ~n6755 & n6773;
  assign n6775 = ~n5794 & n6751;
  assign n6776 = ~n6774 & ~n6775;
  assign n6777 = n1362 & ~n6776;
  assign n6778 = n6758 & n6773;
  assign n6779 = n5790 & ~n5794;
  assign n6780 = n6751 ^ n1362;
  assign n6781 = n6780 ^ n6751;
  assign n6782 = n6758 ^ n6751;
  assign n6783 = n6781 & n6782;
  assign n6784 = n6783 ^ n6751;
  assign n6785 = ~n6779 & n6784;
  assign n6786 = ~n6778 & ~n6785;
  assign n6787 = ~n6777 & n6786;
  assign n6788 = n6787 ^ n6770;
  assign n6789 = n6788 ^ n6770;
  assign n6790 = ~n6772 & n6789;
  assign n6791 = n6790 ^ n6770;
  assign n6792 = ~n5812 & ~n6791;
  assign n6793 = n6792 ^ n6770;
  assign n6794 = n5800 & ~n6793;
  assign n6795 = n5790 & n5812;
  assign n6796 = n6795 ^ n6787;
  assign n6797 = ~n6770 & n6796;
  assign n6798 = ~n6794 & ~n6797;
  assign n7238 = n6798 ^ n6747;
  assign n7239 = ~n6748 & ~n7238;
  assign n7240 = n7239 ^ n6798;
  assign n1074 = x902 ^ x901;
  assign n1073 = x904 ^ x903;
  assign n1075 = n1074 ^ n1073;
  assign n1072 = x906 ^ x905;
  assign n1076 = n1075 ^ n1072;
  assign n1079 = x896 ^ x895;
  assign n1078 = x898 ^ x897;
  assign n1080 = n1079 ^ n1078;
  assign n1077 = x900 ^ x899;
  assign n1081 = n1080 ^ n1077;
  assign n1752 = n1076 & n1081;
  assign n1779 = x899 & x900;
  assign n1780 = x897 & x898;
  assign n1781 = ~n1779 & ~n1780;
  assign n1782 = ~x899 & ~x900;
  assign n1783 = ~x897 & ~x898;
  assign n1784 = ~n1782 & ~n1783;
  assign n1785 = ~n1781 & n1784;
  assign n1786 = x896 & n1785;
  assign n1787 = n1779 & n1780;
  assign n1788 = ~n1786 & ~n1787;
  assign n1789 = n1781 & ~n1784;
  assign n1790 = ~x896 & n1789;
  assign n1791 = n1788 & ~n1790;
  assign n1792 = ~x895 & ~n1791;
  assign n1793 = n1782 & n1783;
  assign n1794 = n1079 & n1793;
  assign n1795 = n1785 ^ x896;
  assign n1796 = n1795 ^ n1785;
  assign n1797 = ~n1787 & ~n1789;
  assign n1798 = n1797 ^ n1785;
  assign n1799 = n1796 & n1798;
  assign n1800 = n1799 ^ n1785;
  assign n1801 = x895 & n1800;
  assign n1802 = ~n1794 & ~n1801;
  assign n1803 = ~n1792 & n1802;
  assign n1756 = x905 & x906;
  assign n1757 = n1756 ^ x904;
  assign n1758 = ~n1073 & ~n1757;
  assign n1759 = ~x901 & n1758;
  assign n1760 = x903 & x904;
  assign n1761 = ~x905 & ~x906;
  assign n1762 = ~n1760 & n1761;
  assign n1763 = ~x902 & n1762;
  assign n1764 = ~n1759 & ~n1763;
  assign n1765 = ~x903 & ~x904;
  assign n1766 = x901 & ~n1765;
  assign n1767 = x902 & ~n1761;
  assign n1768 = ~n1766 & ~n1767;
  assign n1769 = ~n1764 & n1768;
  assign n1770 = n1756 & ~n1765;
  assign n1771 = n1760 & ~n1761;
  assign n1772 = ~n1770 & ~n1771;
  assign n1773 = n1074 & ~n1772;
  assign n1774 = x901 & x902;
  assign n1775 = ~n1762 & n1774;
  assign n1776 = ~n1758 & n1775;
  assign n1777 = ~n1773 & ~n1776;
  assign n1778 = ~n1769 & n1777;
  assign n1804 = n1803 ^ n1778;
  assign n5864 = n1752 & n1804;
  assign n1082 = n1081 ^ n1076;
  assign n1090 = x908 ^ x907;
  assign n1089 = x912 ^ x911;
  assign n1091 = n1090 ^ n1089;
  assign n1088 = x910 ^ x909;
  assign n1092 = n1091 ^ n1088;
  assign n1085 = x914 ^ x913;
  assign n1084 = x918 ^ x917;
  assign n1086 = n1085 ^ n1084;
  assign n1083 = x916 ^ x915;
  assign n1087 = n1086 ^ n1083;
  assign n1093 = n1092 ^ n1087;
  assign n1749 = n1093 ^ n1081;
  assign n1750 = ~n1082 & n1749;
  assign n1751 = n1750 ^ n1093;
  assign n5865 = ~n1751 & ~n1804;
  assign n1748 = n1087 & n1092;
  assign n1753 = n1752 ^ n1751;
  assign n1754 = ~n1748 & ~n1753;
  assign n1755 = n1754 ^ n1752;
  assign n1805 = n1804 ^ n1755;
  assign n1722 = x909 & x910;
  assign n1723 = x911 & x912;
  assign n1724 = ~n1722 & ~n1723;
  assign n1725 = ~x909 & ~x910;
  assign n1726 = ~x911 & ~x912;
  assign n1727 = ~n1725 & ~n1726;
  assign n1728 = ~n1724 & n1727;
  assign n1729 = x908 & n1728;
  assign n1730 = n1722 & n1723;
  assign n1731 = ~n1729 & ~n1730;
  assign n1732 = n1724 & ~n1727;
  assign n1733 = ~x908 & n1732;
  assign n1734 = n1731 & ~n1733;
  assign n1735 = ~x907 & ~n1734;
  assign n1736 = n1725 & n1726;
  assign n1737 = n1090 & n1736;
  assign n1738 = n1728 ^ x908;
  assign n1739 = n1738 ^ n1728;
  assign n1740 = ~n1730 & ~n1732;
  assign n1741 = n1740 ^ n1728;
  assign n1742 = n1739 & n1741;
  assign n1743 = n1742 ^ n1728;
  assign n1744 = x907 & n1743;
  assign n1745 = ~n1737 & ~n1744;
  assign n1746 = ~n1735 & n1745;
  assign n1680 = x915 & x916;
  assign n1679 = x917 & x918;
  assign n1681 = n1680 ^ n1679;
  assign n1682 = ~x915 & ~x916;
  assign n1683 = ~x917 & ~x918;
  assign n1684 = ~n1682 & ~n1683;
  assign n1685 = n1684 ^ n1679;
  assign n1686 = n1685 ^ n1679;
  assign n1687 = n1679 ^ x914;
  assign n1688 = n1687 ^ n1679;
  assign n1689 = n1686 & n1688;
  assign n1690 = n1689 ^ n1679;
  assign n1691 = n1681 & ~n1690;
  assign n1692 = n1691 ^ n1680;
  assign n1693 = x917 ^ x914;
  assign n1694 = n1084 & n1693;
  assign n1695 = n1694 ^ x917;
  assign n1696 = n1682 & ~n1695;
  assign n1697 = ~n1692 & ~n1696;
  assign n1698 = ~x913 & ~n1697;
  assign n1700 = x913 & ~n1682;
  assign n1699 = x913 & x914;
  assign n1701 = n1700 ^ n1699;
  assign n1702 = n1701 ^ n1699;
  assign n1703 = ~x914 & ~x918;
  assign n1704 = n1703 ^ n1699;
  assign n1705 = n1704 ^ n1699;
  assign n1706 = ~n1702 & n1705;
  assign n1707 = n1706 ^ n1699;
  assign n1708 = ~n1680 & n1707;
  assign n1709 = n1708 ^ n1699;
  assign n1710 = ~x917 & n1709;
  assign n1711 = ~n1679 & ~n1680;
  assign n1712 = n1684 & ~n1711;
  assign n1713 = n1085 & n1712;
  assign n1714 = ~n1684 & n1711;
  assign n1715 = n1680 & n1699;
  assign n1716 = x918 & n1715;
  assign n1717 = n1716 ^ n1699;
  assign n1718 = ~n1714 & n1717;
  assign n1719 = ~n1713 & ~n1718;
  assign n1720 = ~n1710 & n1719;
  assign n1721 = ~n1698 & n1720;
  assign n1747 = n1746 ^ n1721;
  assign n1806 = n1805 ^ n1747;
  assign n5866 = n1806 ^ n1805;
  assign n5867 = n1805 ^ n1748;
  assign n5868 = n5866 & ~n5867;
  assign n5869 = n5868 ^ n1805;
  assign n5870 = ~n5865 & n5869;
  assign n5871 = ~n5864 & n5870;
  assign n5848 = n1778 ^ n1752;
  assign n5849 = n1804 & ~n5848;
  assign n5850 = n5849 ^ n1803;
  assign n5854 = n1788 & ~n1801;
  assign n5852 = n1756 & n1760;
  assign n5853 = n1777 & ~n5852;
  assign n5855 = n5854 ^ n5853;
  assign n5851 = ~n1692 & n1719;
  assign n5858 = n1731 & ~n1744;
  assign n5859 = n1747 & n1748;
  assign n5860 = n1721 & n1746;
  assign n5861 = ~n5859 & ~n5860;
  assign n6834 = ~n5858 & ~n5861;
  assign n6835 = ~n5851 & n6834;
  assign n6836 = n6835 ^ n5853;
  assign n6837 = n6836 ^ n6835;
  assign n6838 = n5858 & n5861;
  assign n6839 = n5851 & n6838;
  assign n6840 = n6839 ^ n6835;
  assign n6841 = n6840 ^ n6835;
  assign n6842 = n6837 & n6841;
  assign n6843 = n6842 ^ n6835;
  assign n6844 = ~n5855 & n6843;
  assign n6845 = n6844 ^ n6835;
  assign n5862 = n5861 ^ n5858;
  assign n5856 = n5855 ^ n5851;
  assign n5857 = n5856 ^ n5850;
  assign n5863 = n5862 ^ n5857;
  assign n6846 = n6845 ^ n5863;
  assign n6847 = n6846 ^ n6845;
  assign n6848 = ~n5853 & ~n5854;
  assign n6849 = ~n6834 & n6848;
  assign n6850 = ~n6839 & n6849;
  assign n6853 = ~n5851 & n5855;
  assign n6851 = n5853 & n5854;
  assign n6852 = n6851 ^ n5851;
  assign n6854 = n6853 ^ n6852;
  assign n6855 = n6854 ^ n6853;
  assign n6856 = n6853 ^ n5858;
  assign n6857 = n6856 ^ n6853;
  assign n6858 = n6855 & ~n6857;
  assign n6859 = n6858 ^ n6853;
  assign n6860 = ~n5862 & n6859;
  assign n6861 = n6860 ^ n6853;
  assign n6862 = ~n6850 & ~n6861;
  assign n6863 = n6862 ^ n6845;
  assign n6864 = n6863 ^ n6845;
  assign n6865 = ~n6847 & n6864;
  assign n6866 = n6865 ^ n6845;
  assign n6867 = ~n5850 & n6866;
  assign n6868 = n6867 ^ n6845;
  assign n6869 = n5871 & n6868;
  assign n6870 = ~n5863 & n5871;
  assign n6871 = ~n6845 & ~n6870;
  assign n6872 = ~n5850 & ~n5863;
  assign n6873 = n6872 ^ n6862;
  assign n6874 = n6871 & n6873;
  assign n6875 = ~n6869 & ~n6874;
  assign n5872 = n5871 ^ n5863;
  assign n1651 = x941 & x942;
  assign n1652 = x939 & x940;
  assign n1653 = ~n1651 & ~n1652;
  assign n1654 = ~x941 & ~x942;
  assign n1655 = ~x939 & ~x940;
  assign n1656 = ~n1654 & ~n1655;
  assign n1657 = ~n1653 & n1656;
  assign n1658 = x938 & n1657;
  assign n1659 = n1651 & n1652;
  assign n1660 = ~n1658 & ~n1659;
  assign n1661 = n1653 & ~n1656;
  assign n1662 = ~x938 & n1661;
  assign n1663 = n1660 & ~n1662;
  assign n1664 = ~x937 & ~n1663;
  assign n1056 = x938 ^ x937;
  assign n1665 = n1654 & n1655;
  assign n1666 = n1056 & n1665;
  assign n1667 = n1657 ^ x938;
  assign n1668 = n1667 ^ n1657;
  assign n1669 = ~n1659 & ~n1661;
  assign n1670 = n1669 ^ n1657;
  assign n1671 = n1668 & n1670;
  assign n1672 = n1671 ^ n1657;
  assign n1673 = x937 & n1672;
  assign n1674 = ~n1666 & ~n1673;
  assign n1675 = ~n1664 & n1674;
  assign n1621 = x933 & x934;
  assign n1622 = x935 & x936;
  assign n1623 = n1621 & n1622;
  assign n1624 = ~x933 & ~x934;
  assign n1625 = ~n1622 & n1624;
  assign n1626 = n1625 ^ x932;
  assign n1627 = ~x935 & ~x936;
  assign n1628 = n1627 ^ n1625;
  assign n1629 = n1628 ^ n1627;
  assign n1630 = ~n1621 & n1627;
  assign n1631 = n1630 ^ n1627;
  assign n1632 = ~n1629 & ~n1631;
  assign n1633 = n1632 ^ n1627;
  assign n1634 = ~n1626 & n1633;
  assign n1635 = n1634 ^ x932;
  assign n1636 = ~n1623 & n1635;
  assign n1637 = ~x931 & ~n1636;
  assign n1638 = x931 & x932;
  assign n1639 = ~n1625 & n1638;
  assign n1640 = ~n1623 & ~n1630;
  assign n1641 = n1639 & n1640;
  assign n1051 = x932 ^ x931;
  assign n1642 = n1622 & ~n1624;
  assign n1643 = n1621 & ~n1627;
  assign n1644 = ~n1642 & ~n1643;
  assign n1645 = n1051 & ~n1644;
  assign n1646 = ~n1641 & ~n1645;
  assign n1647 = ~x932 & n1630;
  assign n1648 = n1624 & n1647;
  assign n1649 = n1646 & ~n1648;
  assign n1650 = ~n1637 & n1649;
  assign n1676 = n1675 ^ n1650;
  assign n1579 = x929 & x930;
  assign n1578 = x927 & x928;
  assign n1580 = n1579 ^ n1578;
  assign n1581 = ~x929 & ~x930;
  assign n1582 = ~x927 & ~x928;
  assign n1583 = ~n1581 & ~n1582;
  assign n1584 = n1583 ^ n1578;
  assign n1585 = n1584 ^ n1578;
  assign n1586 = n1578 ^ x926;
  assign n1587 = n1586 ^ n1578;
  assign n1588 = n1585 & n1587;
  assign n1589 = n1588 ^ n1578;
  assign n1590 = n1580 & ~n1589;
  assign n1591 = n1590 ^ n1579;
  assign n1592 = ~n1578 & ~n1579;
  assign n1593 = n1582 ^ n1581;
  assign n1594 = n1581 ^ x926;
  assign n1595 = n1593 & ~n1594;
  assign n1596 = n1595 ^ n1581;
  assign n1597 = n1592 & n1596;
  assign n1598 = ~n1591 & ~n1597;
  assign n1599 = ~x925 & ~n1598;
  assign n1067 = x926 ^ x925;
  assign n1600 = n1583 & ~n1592;
  assign n1601 = n1067 & n1600;
  assign n1602 = ~n1583 & n1592;
  assign n1603 = x925 & x926;
  assign n1604 = n1578 & n1603;
  assign n1605 = x930 & n1604;
  assign n1606 = n1605 ^ n1603;
  assign n1607 = ~n1602 & n1606;
  assign n1608 = ~n1601 & ~n1607;
  assign n1066 = x928 ^ x927;
  assign n1609 = n1603 ^ x928;
  assign n1610 = n1609 ^ n1603;
  assign n1611 = ~x926 & ~x930;
  assign n1612 = n1611 ^ n1603;
  assign n1613 = ~n1610 & n1612;
  assign n1614 = n1613 ^ n1603;
  assign n1615 = ~n1066 & n1614;
  assign n1616 = ~x929 & n1615;
  assign n1617 = n1608 & ~n1616;
  assign n1618 = ~n1599 & n1617;
  assign n1062 = x920 ^ x919;
  assign n1555 = ~x921 & ~x922;
  assign n1556 = x923 & x924;
  assign n1557 = ~n1555 & n1556;
  assign n1558 = x921 & x922;
  assign n1559 = ~x923 & ~x924;
  assign n1560 = n1558 & ~n1559;
  assign n1561 = ~n1557 & ~n1560;
  assign n1562 = n1062 & ~n1561;
  assign n1563 = ~n1558 & n1559;
  assign n1564 = x919 & x920;
  assign n1565 = ~n1563 & n1564;
  assign n1061 = x922 ^ x921;
  assign n1566 = n1556 ^ x922;
  assign n1567 = ~n1061 & ~n1566;
  assign n1568 = n1565 & ~n1567;
  assign n1569 = ~n1562 & ~n1568;
  assign n1570 = ~x919 & n1567;
  assign n1571 = ~x920 & n1563;
  assign n1572 = ~n1570 & ~n1571;
  assign n1573 = x919 & ~n1555;
  assign n1574 = x920 & ~n1559;
  assign n1575 = ~n1573 & ~n1574;
  assign n1576 = ~n1572 & n1575;
  assign n1577 = n1569 & ~n1576;
  assign n1619 = n1618 ^ n1577;
  assign n1050 = x934 ^ x933;
  assign n1052 = n1051 ^ n1050;
  assign n1049 = x936 ^ x935;
  assign n1053 = n1052 ^ n1049;
  assign n1055 = x940 ^ x939;
  assign n1057 = n1056 ^ n1055;
  assign n1054 = x942 ^ x941;
  assign n1058 = n1057 ^ n1054;
  assign n1547 = n1053 & n1058;
  assign n1063 = n1062 ^ n1061;
  assign n1060 = x924 ^ x923;
  assign n1064 = n1063 ^ n1060;
  assign n1068 = n1067 ^ n1066;
  assign n1065 = x930 ^ x929;
  assign n1069 = n1068 ^ n1065;
  assign n1551 = n1064 & n1069;
  assign n1070 = n1069 ^ n1064;
  assign n1059 = n1058 ^ n1053;
  assign n1548 = n1064 ^ n1059;
  assign n1549 = n1070 & ~n1548;
  assign n1550 = n1549 ^ n1069;
  assign n1552 = n1551 ^ n1550;
  assign n1553 = ~n1547 & ~n1552;
  assign n1554 = n1553 ^ n1551;
  assign n1620 = n1619 ^ n1554;
  assign n1677 = n1676 ^ n1620;
  assign n1071 = n1070 ^ n1059;
  assign n1094 = n1093 ^ n1082;
  assign n1546 = n1071 & n1094;
  assign n1678 = n1677 ^ n1546;
  assign n5845 = n1806 ^ n1546;
  assign n5846 = ~n1678 & n5845;
  assign n5847 = n5846 ^ n1677;
  assign n5873 = n5872 ^ n5847;
  assign n5888 = n1660 & ~n1673;
  assign n5889 = ~n1623 & n1646;
  assign n5890 = ~n5888 & ~n5889;
  assign n5891 = n1650 ^ n1547;
  assign n5892 = n1676 & ~n5891;
  assign n5893 = n5892 ^ n1675;
  assign n5894 = n5890 & n5893;
  assign n5895 = n5893 ^ n5888;
  assign n5896 = n5889 ^ n5888;
  assign n5897 = ~n5895 & ~n5896;
  assign n5898 = n5897 ^ n5893;
  assign n5899 = ~n5894 & n5898;
  assign n5900 = n5888 & n5889;
  assign n5901 = ~n5893 & n5900;
  assign n5902 = ~n5899 & ~n5901;
  assign n5886 = ~n1591 & n1608;
  assign n5884 = n1556 & n1558;
  assign n5885 = n1569 & ~n5884;
  assign n5887 = n5886 ^ n5885;
  assign n5903 = n5902 ^ n5887;
  assign n5881 = n1577 ^ n1551;
  assign n5882 = n1619 & ~n5881;
  assign n5883 = n5882 ^ n1618;
  assign n5904 = n5903 ^ n5883;
  assign n5874 = n1551 & n1619;
  assign n5875 = ~n1620 & ~n1676;
  assign n5876 = n1547 & n1676;
  assign n5877 = ~n1550 & ~n1619;
  assign n5878 = ~n5876 & ~n5877;
  assign n5879 = ~n5875 & n5878;
  assign n5880 = ~n5874 & n5879;
  assign n5905 = n5904 ^ n5880;
  assign n6831 = n5905 ^ n5872;
  assign n6832 = ~n5873 & ~n6831;
  assign n6833 = n6832 ^ n5905;
  assign n6876 = n6875 ^ n6833;
  assign n6803 = n5901 ^ n5894;
  assign n6804 = n5886 & n6803;
  assign n6805 = n6804 ^ n5894;
  assign n6806 = n5904 & n6805;
  assign n6807 = ~n5883 & n5885;
  assign n6808 = ~n5898 & n6807;
  assign n6809 = ~n5886 & ~n5901;
  assign n6810 = n6808 & ~n6809;
  assign n6811 = n5887 & n5894;
  assign n6812 = ~n6810 & ~n6811;
  assign n6813 = ~n6806 & n6812;
  assign n6814 = n5880 & n5904;
  assign n6815 = ~n5883 & n5903;
  assign n6816 = ~n5885 & ~n5886;
  assign n6817 = ~n5890 & n6816;
  assign n6818 = ~n5901 & n6817;
  assign n6819 = n5885 & n5886;
  assign n6820 = n6819 ^ n5899;
  assign n6821 = n6820 ^ n5899;
  assign n6822 = n5899 ^ n5894;
  assign n6823 = n6821 & n6822;
  assign n6824 = n6823 ^ n5899;
  assign n6825 = ~n6818 & ~n6824;
  assign n6826 = ~n6815 & ~n6825;
  assign n6827 = ~n6814 & ~n6826;
  assign n6828 = n6827 ^ n6814;
  assign n6829 = n6813 & n6828;
  assign n6830 = n6829 ^ n6814;
  assign n6877 = n6876 ^ n6830;
  assign n5843 = n5842 ^ n5813;
  assign n1807 = n1806 ^ n1678;
  assign n1048 = n1047 ^ n1024;
  assign n1095 = n1094 ^ n1071;
  assign n1096 = n1048 & n1095;
  assign n5784 = n1807 ^ n1096;
  assign n1545 = n1544 ^ n1384;
  assign n5785 = n1545 ^ n1096;
  assign n5786 = n5784 & n5785;
  assign n5787 = n5786 ^ n1807;
  assign n5844 = n5843 ^ n5787;
  assign n5906 = n5905 ^ n5873;
  assign n6800 = n5906 ^ n5843;
  assign n6801 = n5844 & ~n6800;
  assign n6802 = n6801 ^ n5906;
  assign n6878 = n6877 ^ n6802;
  assign n6799 = n6798 ^ n6748;
  assign n7241 = n6802 ^ n6799;
  assign n7242 = ~n6878 & n7241;
  assign n7243 = n7242 ^ n6877;
  assign n7528 = n7240 & n7243;
  assign n7231 = ~n6835 & ~n6875;
  assign n7232 = ~n5850 & n6851;
  assign n7233 = ~n6839 & ~n7232;
  assign n7234 = ~n7231 & n7233;
  assign n7228 = n6875 ^ n6830;
  assign n7229 = ~n6876 & n7228;
  assign n7230 = n7229 ^ n6833;
  assign n7235 = n7234 ^ n7230;
  assign n7224 = ~n5886 & n5893;
  assign n7225 = n6830 & ~n7224;
  assign n7226 = ~n5890 & n6827;
  assign n7227 = ~n7225 & ~n7226;
  assign n7236 = n7235 ^ n7227;
  assign n7216 = ~n6740 & n6747;
  assign n7217 = ~n6726 & n6730;
  assign n7218 = ~n7216 & ~n7217;
  assign n7219 = ~n6759 & n6797;
  assign n7220 = ~n6758 & ~n6774;
  assign n7221 = ~n7219 & n7220;
  assign n7222 = ~n6794 & n7221;
  assign n7534 = n7218 & n7222;
  assign n7536 = ~n7236 & ~n7534;
  assign n7537 = n7528 & n7536;
  assign n7529 = n7236 & ~n7528;
  assign n7535 = n7529 & n7534;
  assign n7530 = ~n7240 & ~n7243;
  assign n7531 = ~n7529 & ~n7530;
  assign n7532 = ~n7218 & ~n7222;
  assign n7533 = n7531 & n7532;
  assign n7525 = n7234 ^ n7227;
  assign n7526 = n7235 & ~n7525;
  assign n7527 = n7526 ^ n7230;
  assign n7538 = n7236 & ~n7532;
  assign n7539 = n7530 & n7538;
  assign n7692 = ~n7527 & ~n7539;
  assign n7693 = ~n7533 & ~n7692;
  assign n7694 = ~n7535 & ~n7693;
  assign n7695 = ~n7537 & ~n7694;
  assign n7741 = ~n7688 & n7695;
  assign n7742 = ~n7690 & ~n7741;
  assign n7523 = n7522 ^ n7515;
  assign n7328 = n7327 ^ n7266;
  assign n6719 = n6718 ^ n6675;
  assign n5907 = n5906 ^ n5844;
  assign n2796 = n2795 ^ n2170;
  assign n1231 = n1230 ^ n1143;
  assign n1232 = n1095 ^ n1048;
  assign n1233 = n1231 & n1232;
  assign n5776 = n2796 ^ n1233;
  assign n1808 = n1807 ^ n1545;
  assign n1234 = ~n1096 & ~n1233;
  assign n1809 = n1808 ^ n1234;
  assign n5777 = n1809 ^ n1808;
  assign n5778 = n1808 ^ n1233;
  assign n5779 = n5778 ^ n1808;
  assign n5780 = n5777 & ~n5779;
  assign n5781 = n5780 ^ n1808;
  assign n5782 = n5776 & ~n5781;
  assign n5783 = n5782 ^ n2796;
  assign n5908 = n5907 ^ n5783;
  assign n6090 = n6089 ^ n5977;
  assign n6608 = n6090 ^ n5783;
  assign n6609 = ~n5908 & n6608;
  assign n6610 = n6609 ^ n5907;
  assign n6720 = n6719 ^ n6610;
  assign n6879 = n6878 ^ n6799;
  assign n7246 = n6879 ^ n6610;
  assign n7247 = ~n6720 & n7246;
  assign n7248 = n7247 ^ n6719;
  assign n7329 = n7328 ^ n7248;
  assign n7244 = n7243 ^ n7240;
  assign n7223 = n7222 ^ n7218;
  assign n7237 = n7236 ^ n7223;
  assign n7245 = n7244 ^ n7237;
  assign n7504 = n7248 ^ n7245;
  assign n7505 = n7329 & ~n7504;
  assign n7506 = n7505 ^ n7328;
  assign n7524 = n7523 ^ n7506;
  assign n7540 = ~n7537 & ~n7539;
  assign n7541 = ~n7535 & n7540;
  assign n7542 = ~n7533 & n7541;
  assign n7543 = n7542 ^ n7527;
  assign n7680 = n7543 ^ n7523;
  assign n7681 = ~n7524 & n7680;
  assign n7682 = n7681 ^ n7543;
  assign n7743 = n7688 & ~n7695;
  assign n7744 = n7682 & ~n7743;
  assign n7745 = n7742 & ~n7744;
  assign n7691 = ~n7688 & ~n7690;
  assign n7696 = n7695 ^ n7691;
  assign n7697 = n7696 ^ n7682;
  assign n7544 = n7543 ^ n7524;
  assign n7330 = n7329 ^ n7245;
  assign n6880 = n6879 ^ n6720;
  assign n6091 = n6090 ^ n5908;
  assign n2797 = n2796 ^ n1809;
  assign n3181 = n3180 ^ n2797;
  assign n3182 = n1232 ^ n1231;
  assign n3183 = n3182 ^ n2797;
  assign n5758 = n5757 ^ n4527;
  assign n5759 = n5758 ^ n2797;
  assign n5760 = ~n2797 & ~n5759;
  assign n5761 = n5760 ^ n2797;
  assign n5762 = n3183 & ~n5761;
  assign n5763 = n5762 ^ n5760;
  assign n5764 = n5763 ^ n2797;
  assign n5765 = n5764 ^ n5758;
  assign n5766 = ~n3181 & ~n5765;
  assign n5767 = n5766 ^ n2797;
  assign n5768 = ~n3182 & ~n5758;
  assign n5769 = n5768 ^ n3179;
  assign n5770 = n2797 & n5758;
  assign n5771 = ~n2988 & ~n5770;
  assign n5772 = n5771 ^ n3179;
  assign n5773 = ~n5769 & ~n5772;
  assign n5774 = n5773 ^ n3179;
  assign n5775 = n5767 & n5774;
  assign n6092 = n6091 ^ n5775;
  assign n6604 = n6603 ^ n6339;
  assign n6605 = n6604 ^ n6091;
  assign n6606 = n6092 & n6605;
  assign n6607 = n6606 ^ n5775;
  assign n6881 = n6880 ^ n6607;
  assign n7212 = n7211 ^ n7041;
  assign n7213 = n7212 ^ n6607;
  assign n7214 = ~n6881 & n7213;
  assign n7215 = n7214 ^ n6880;
  assign n7331 = n7330 ^ n7215;
  assign n7500 = n7499 ^ n7334;
  assign n7501 = n7500 ^ n7330;
  assign n7502 = n7331 & ~n7501;
  assign n7503 = n7502 ^ n7500;
  assign n7545 = n7544 ^ n7503;
  assign n7676 = n7675 ^ n7612;
  assign n7677 = n7676 ^ n7503;
  assign n7678 = n7545 & n7677;
  assign n7679 = n7678 ^ n7676;
  assign n7698 = n7697 ^ n7679;
  assign n7736 = n7735 ^ n7711;
  assign n7707 = n7706 ^ n7703;
  assign n7708 = n7707 ^ n7700;
  assign n7737 = n7736 ^ n7708;
  assign n7738 = n7737 ^ n7697;
  assign n7739 = ~n7698 & n7738;
  assign n7740 = n7739 ^ n7679;
  assign n7746 = n7745 ^ n7740;
  assign n7752 = n7711 ^ n7703;
  assign n7753 = n7752 ^ n7711;
  assign n7755 = n7754 ^ n7711;
  assign n7756 = n7755 ^ n7711;
  assign n7757 = n7753 & ~n7756;
  assign n7758 = n7757 ^ n7711;
  assign n7759 = n7707 & n7758;
  assign n7760 = n7759 ^ n7711;
  assign n7761 = n7700 & n7760;
  assign n7762 = ~n7560 & ~n7700;
  assign n7763 = n7552 & n7558;
  assign n7764 = ~n7762 & ~n7763;
  assign n7765 = n7560 & n7590;
  assign n7766 = n6941 & n7765;
  assign n7767 = ~n7764 & ~n7766;
  assign n7768 = ~n7560 & ~n7609;
  assign n7769 = n7700 & ~n7768;
  assign n7770 = ~n7552 & ~n7558;
  assign n7771 = ~n7769 & ~n7770;
  assign n7772 = ~n7767 & ~n7771;
  assign n7773 = n7555 & ~n7772;
  assign n7774 = n7735 & ~n7773;
  assign n7775 = ~n7566 & n7604;
  assign n7776 = ~n7764 & n7771;
  assign n7777 = ~n7775 & ~n7776;
  assign n7778 = n7774 & n7777;
  assign n7779 = ~n7761 & ~n7778;
  assign n7782 = n7780 & ~n7781;
  assign n7783 = n7736 ^ n7735;
  assign n7785 = n7784 ^ n7735;
  assign n7786 = ~n7783 & n7785;
  assign n7787 = n7786 ^ n7735;
  assign n7788 = ~n7700 & ~n7787;
  assign n7789 = ~n7782 & n7788;
  assign n7790 = n7779 & ~n7789;
  assign n7791 = n7790 ^ n7751;
  assign n7792 = n7791 ^ n7740;
  assign n7793 = ~n7746 & n7792;
  assign n7794 = n7793 ^ n7791;
  assign n7811 = n7810 ^ n7794;
  assign n11861 = n7791 ^ n7746;
  assign n8286 = x659 & x660;
  assign n8287 = x657 & x658;
  assign n8288 = ~n8286 & ~n8287;
  assign n8289 = ~x659 & ~x660;
  assign n8290 = ~x657 & ~x658;
  assign n8291 = ~n8289 & ~n8290;
  assign n8292 = ~n8288 & n8291;
  assign n8293 = x656 & n8292;
  assign n8294 = n8286 & n8287;
  assign n8295 = ~n8293 & ~n8294;
  assign n8296 = n8288 & ~n8291;
  assign n8297 = ~x656 & n8296;
  assign n8298 = n8295 & ~n8297;
  assign n8299 = ~x655 & ~n8298;
  assign n7914 = x656 ^ x655;
  assign n8300 = n8289 & n8290;
  assign n8301 = n7914 & n8300;
  assign n8302 = n8292 ^ x656;
  assign n8303 = n8302 ^ n8292;
  assign n8304 = ~n8294 & ~n8296;
  assign n8305 = n8304 ^ n8292;
  assign n8306 = n8303 & n8305;
  assign n8307 = n8306 ^ n8292;
  assign n8308 = x655 & n8307;
  assign n8309 = ~n8301 & ~n8308;
  assign n8310 = ~n8299 & n8309;
  assign n8261 = x665 & x666;
  assign n8262 = ~x663 & ~x664;
  assign n8263 = ~n8261 & n8262;
  assign n8264 = ~x665 & ~x666;
  assign n8265 = x662 & ~n8264;
  assign n8266 = n8263 & ~n8265;
  assign n8267 = x663 & x664;
  assign n8268 = n8261 & n8267;
  assign n8269 = ~n8266 & ~n8268;
  assign n8270 = n8264 & ~n8267;
  assign n8271 = ~x662 & n8270;
  assign n8272 = n8269 & ~n8271;
  assign n8273 = ~x661 & ~n8272;
  assign n8274 = ~n8263 & ~n8268;
  assign n8275 = x661 & x662;
  assign n8276 = ~n8270 & n8275;
  assign n8277 = n8274 & n8276;
  assign n7909 = x662 ^ x661;
  assign n8278 = n8261 & ~n8262;
  assign n8279 = ~n8264 & n8267;
  assign n8280 = ~n8278 & ~n8279;
  assign n8281 = n7909 & ~n8280;
  assign n8282 = ~n8277 & ~n8281;
  assign n8283 = n8262 & n8271;
  assign n8284 = n8282 & ~n8283;
  assign n8285 = ~n8273 & n8284;
  assign n8311 = n8310 ^ n8285;
  assign n7908 = x664 ^ x663;
  assign n7910 = n7909 ^ n7908;
  assign n7907 = x666 ^ x665;
  assign n7911 = n7910 ^ n7907;
  assign n7913 = x658 ^ x657;
  assign n7915 = n7914 ^ n7913;
  assign n7912 = x660 ^ x659;
  assign n7916 = n7915 ^ n7912;
  assign n8253 = n7911 & n7916;
  assign n10792 = n8285 ^ n8253;
  assign n10793 = n8311 & ~n10792;
  assign n10794 = n10793 ^ n8310;
  assign n10795 = ~n8268 & n8282;
  assign n11417 = n10794 & ~n10795;
  assign n8213 = ~x671 & ~x672;
  assign n8214 = x668 & ~n8213;
  assign n8215 = x671 & x672;
  assign n8216 = ~x669 & ~x670;
  assign n8217 = ~n8215 & n8216;
  assign n8218 = ~n8214 & n8217;
  assign n8219 = x669 & x670;
  assign n8220 = n8219 ^ n8215;
  assign n8221 = n8219 ^ n8214;
  assign n8222 = n8220 & n8221;
  assign n8223 = n8222 ^ n8219;
  assign n8224 = ~n8216 & n8223;
  assign n8225 = ~n8218 & ~n8224;
  assign n8226 = ~x667 & ~n8225;
  assign n8227 = ~n8215 & ~n8219;
  assign n8228 = ~n8216 & ~n8227;
  assign n8229 = x667 & ~n8213;
  assign n8230 = n8228 & n8229;
  assign n8231 = x667 & x668;
  assign n8232 = ~n8230 & ~n8231;
  assign n8233 = ~n8213 & ~n8219;
  assign n8234 = ~n8217 & n8233;
  assign n8235 = ~x672 & n8219;
  assign n8236 = x668 & ~n8235;
  assign n8237 = ~n8234 & n8236;
  assign n8238 = ~n8232 & ~n8237;
  assign n8239 = ~n8226 & ~n8238;
  assign n8240 = ~x668 & ~x672;
  assign n8241 = n8240 ^ n8231;
  assign n8242 = n8241 ^ n8231;
  assign n8243 = x667 & ~n8216;
  assign n8244 = n8243 ^ n8231;
  assign n8245 = n8244 ^ n8231;
  assign n8246 = n8242 & ~n8245;
  assign n8247 = n8246 ^ n8231;
  assign n8248 = ~n8219 & n8247;
  assign n8249 = n8248 ^ n8231;
  assign n8250 = ~x671 & n8249;
  assign n8251 = n8239 & ~n8250;
  assign n8176 = ~x677 & ~x678;
  assign n8177 = x673 & ~n8176;
  assign n7919 = x676 ^ x675;
  assign n8178 = x677 & x678;
  assign n8179 = n8178 ^ x676;
  assign n8180 = n7919 & ~n8179;
  assign n8181 = n8180 ^ x675;
  assign n8182 = n8177 & n8181;
  assign n8183 = x673 & x674;
  assign n8184 = ~n8182 & ~n8183;
  assign n8185 = ~x675 & ~x676;
  assign n8186 = ~n8178 & n8185;
  assign n8187 = x675 & x676;
  assign n8188 = ~n8176 & ~n8187;
  assign n8189 = ~n8186 & n8188;
  assign n8190 = ~x678 & n8187;
  assign n8191 = x674 & ~n8190;
  assign n8192 = ~n8189 & n8191;
  assign n8193 = ~n8184 & ~n8192;
  assign n8194 = x674 & ~n8176;
  assign n8195 = n8178 & n8187;
  assign n8196 = ~n8194 & ~n8195;
  assign n8197 = n8181 & ~n8196;
  assign n8198 = n8186 & ~n8194;
  assign n8199 = ~n8197 & ~n8198;
  assign n8200 = ~x673 & ~n8199;
  assign n8201 = ~n8193 & ~n8200;
  assign n8202 = ~x674 & ~x678;
  assign n8203 = n8202 ^ n8183;
  assign n8204 = n8203 ^ n8183;
  assign n7920 = x674 ^ x673;
  assign n7921 = n7920 ^ n7919;
  assign n8205 = n8183 ^ n7921;
  assign n8206 = n8205 ^ n8183;
  assign n8207 = n8204 & n8206;
  assign n8208 = n8207 ^ n8183;
  assign n8209 = ~n8187 & n8208;
  assign n8210 = n8209 ^ n8183;
  assign n8211 = ~x677 & n8210;
  assign n8212 = n8201 & ~n8211;
  assign n8252 = n8251 ^ n8212;
  assign n7918 = x678 ^ x677;
  assign n7922 = n7921 ^ n7918;
  assign n7925 = x672 ^ x671;
  assign n7924 = x670 ^ x669;
  assign n7926 = n7925 ^ n7924;
  assign n7923 = x668 ^ x667;
  assign n7927 = n7926 ^ n7923;
  assign n8254 = n7922 & n7927;
  assign n10810 = n8252 & n8254;
  assign n10811 = n8212 & n8251;
  assign n10812 = ~n10810 & ~n10811;
  assign n10808 = ~n8193 & ~n8197;
  assign n10807 = ~n8224 & ~n8238;
  assign n10809 = n10808 ^ n10807;
  assign n10813 = n10812 ^ n10809;
  assign n10799 = n8253 & n8311;
  assign n7928 = n7927 ^ n7922;
  assign n7917 = n7916 ^ n7911;
  assign n8256 = n7922 ^ n7917;
  assign n8257 = n7928 & n8256;
  assign n8258 = n8257 ^ n7922;
  assign n8259 = ~n8253 & ~n8258;
  assign n10800 = n8259 & ~n8311;
  assign n10801 = ~n10799 & ~n10800;
  assign n8255 = n8253 & n8254;
  assign n8260 = ~n8255 & ~n8259;
  assign n8312 = n8311 ^ n8260;
  assign n8313 = n8312 ^ n8252;
  assign n10802 = n8313 ^ n8312;
  assign n10803 = n8312 ^ n8254;
  assign n10804 = n10802 & n10803;
  assign n10805 = n10804 ^ n8312;
  assign n10806 = n10801 & ~n10805;
  assign n10814 = n10813 ^ n10806;
  assign n10797 = n8295 & ~n8308;
  assign n11418 = n10813 ^ n10797;
  assign n11419 = ~n10814 & ~n11418;
  assign n11420 = n11419 ^ n10806;
  assign n11421 = n11417 & ~n11420;
  assign n11422 = ~n10806 & n10813;
  assign n10796 = n10795 ^ n10794;
  assign n11423 = ~n10796 & n10797;
  assign n11424 = ~n11422 & n11423;
  assign n11425 = ~n11421 & ~n11424;
  assign n11426 = ~n10794 & n10795;
  assign n11427 = n11420 & n11426;
  assign n11428 = n10806 & ~n10813;
  assign n11429 = ~n10796 & ~n10797;
  assign n11430 = ~n11428 & n11429;
  assign n11431 = ~n11427 & ~n11430;
  assign n11432 = n11425 & n11431;
  assign n11414 = n10812 ^ n10808;
  assign n11415 = ~n10809 & n11414;
  assign n11416 = n11415 ^ n10812;
  assign n11433 = n11432 ^ n11416;
  assign n11662 = ~n11417 & n11433;
  assign n11663 = n11416 & ~n11420;
  assign n11664 = ~n11662 & ~n11663;
  assign n8125 = x693 & x694;
  assign n8123 = ~x695 & ~x696;
  assign n8124 = x692 & ~n8123;
  assign n8126 = n8125 ^ n8124;
  assign n8127 = x695 & x696;
  assign n8128 = ~x693 & ~x694;
  assign n8129 = n8127 & ~n8128;
  assign n8130 = n8129 ^ n8124;
  assign n8131 = n8130 ^ n8129;
  assign n8132 = n8129 ^ n8127;
  assign n8133 = ~n8131 & ~n8132;
  assign n8134 = n8133 ^ n8129;
  assign n8135 = n8126 & n8134;
  assign n8136 = n8135 ^ n8125;
  assign n8152 = ~n8125 & ~n8129;
  assign n8153 = x691 & ~n8123;
  assign n8154 = ~n8152 & n8153;
  assign n8155 = x691 & x692;
  assign n8156 = ~n8154 & ~n8155;
  assign n8137 = ~n8127 & n8128;
  assign n8157 = ~n8123 & ~n8125;
  assign n8158 = ~n8137 & n8157;
  assign n8159 = ~x696 & n8125;
  assign n8160 = x692 & ~n8159;
  assign n8161 = ~n8158 & n8160;
  assign n8162 = ~n8156 & ~n8161;
  assign n10832 = ~n8136 & ~n8162;
  assign n8082 = x699 & x700;
  assign n8081 = x701 & x702;
  assign n8083 = n8082 ^ n8081;
  assign n8084 = ~x699 & ~x700;
  assign n8085 = ~x701 & ~x702;
  assign n8086 = ~n8084 & ~n8085;
  assign n8087 = n8086 ^ n8081;
  assign n8088 = n8087 ^ n8081;
  assign n8089 = n8081 ^ x698;
  assign n8090 = n8089 ^ n8081;
  assign n8091 = n8088 & n8090;
  assign n8092 = n8091 ^ n8081;
  assign n8093 = n8083 & ~n8092;
  assign n8094 = n8093 ^ n8082;
  assign n8096 = ~n8081 & ~n8082;
  assign n8109 = n8086 & ~n8096;
  assign n8108 = x702 & n8082;
  assign n8110 = n8109 ^ n8108;
  assign n8111 = n8110 ^ n8109;
  assign n8112 = ~n8086 & n8096;
  assign n8113 = n8112 ^ n8109;
  assign n8114 = n8113 ^ n8109;
  assign n8115 = ~n8111 & ~n8114;
  assign n8116 = n8115 ^ n8109;
  assign n8117 = x698 & n8116;
  assign n8118 = n8117 ^ n8109;
  assign n10830 = x697 & n8118;
  assign n10831 = ~n8094 & ~n10830;
  assign n10833 = n10832 ^ n10831;
  assign n8138 = n8137 ^ n8123;
  assign n8139 = n8137 ^ n8125;
  assign n8140 = n8123 ^ x692;
  assign n8141 = n8140 ^ n8137;
  assign n8142 = ~n8137 & ~n8141;
  assign n8143 = n8142 ^ n8137;
  assign n8144 = ~n8139 & ~n8143;
  assign n8145 = n8144 ^ n8142;
  assign n8146 = n8145 ^ n8137;
  assign n8147 = n8146 ^ n8140;
  assign n8148 = n8138 & ~n8147;
  assign n8149 = n8148 ^ n8137;
  assign n8150 = ~n8136 & ~n8149;
  assign n8151 = ~x691 & ~n8150;
  assign n8163 = ~n8151 & ~n8162;
  assign n7948 = x694 ^ x693;
  assign n8164 = n8155 ^ x694;
  assign n8165 = n8164 ^ n8155;
  assign n8166 = ~x692 & ~x696;
  assign n8167 = n8166 ^ n8155;
  assign n8168 = ~n8165 & n8167;
  assign n8169 = n8168 ^ n8155;
  assign n8170 = ~n7948 & n8169;
  assign n8171 = ~x695 & n8170;
  assign n8172 = n8163 & ~n8171;
  assign n7943 = x700 ^ x699;
  assign n8072 = x697 & x698;
  assign n8073 = n8072 ^ x700;
  assign n8074 = n8073 ^ n8072;
  assign n8075 = ~x698 & ~x702;
  assign n8076 = n8075 ^ n8072;
  assign n8077 = ~n8074 & n8076;
  assign n8078 = n8077 ^ n8072;
  assign n8079 = ~n7943 & n8078;
  assign n8080 = ~x701 & n8079;
  assign n8095 = n8085 ^ n8084;
  assign n8097 = n8096 ^ n8085;
  assign n8098 = n8097 ^ n8085;
  assign n8099 = n8085 ^ x698;
  assign n8100 = n8099 ^ n8085;
  assign n8101 = n8098 & ~n8100;
  assign n8102 = n8101 ^ n8085;
  assign n8103 = n8095 & ~n8102;
  assign n8104 = n8103 ^ n8084;
  assign n8105 = ~n8094 & ~n8104;
  assign n8106 = n8105 ^ x697;
  assign n8107 = n8106 ^ n8105;
  assign n8119 = n8118 ^ n8105;
  assign n8120 = n8107 & ~n8119;
  assign n8121 = n8120 ^ n8105;
  assign n8122 = ~n8080 & n8121;
  assign n8173 = n8172 ^ n8122;
  assign n7942 = x702 ^ x701;
  assign n7944 = n7943 ^ n7942;
  assign n7941 = x698 ^ x697;
  assign n7945 = n7944 ^ n7941;
  assign n7947 = x696 ^ x695;
  assign n7949 = n7948 ^ n7947;
  assign n7946 = x692 ^ x691;
  assign n7950 = n7949 ^ n7946;
  assign n8071 = n7945 & n7950;
  assign n10827 = n8122 ^ n8071;
  assign n10828 = n8173 & ~n10827;
  assign n10829 = n10828 ^ n8172;
  assign n10834 = n10833 ^ n10829;
  assign n8010 = ~x689 & ~x690;
  assign n7936 = x688 ^ x687;
  assign n8011 = x689 & x690;
  assign n8012 = n8011 ^ x688;
  assign n8013 = n7936 & ~n8012;
  assign n8014 = n8013 ^ x687;
  assign n8015 = ~n8010 & n8014;
  assign n8016 = ~x686 & ~n8015;
  assign n8019 = x687 & x688;
  assign n8022 = n8010 & ~n8019;
  assign n8017 = ~x687 & ~x688;
  assign n8018 = ~n8011 & n8017;
  assign n8020 = n8011 & n8019;
  assign n8021 = ~n8018 & ~n8020;
  assign n8023 = n8022 ^ n8021;
  assign n8024 = n8021 ^ x685;
  assign n8025 = n8021 & n8024;
  assign n8026 = n8025 ^ n8021;
  assign n8027 = ~n8023 & n8026;
  assign n8028 = n8027 ^ n8025;
  assign n8029 = n8028 ^ n8021;
  assign n8030 = n8029 ^ x685;
  assign n8031 = x686 & n8030;
  assign n8032 = n8031 ^ x685;
  assign n8033 = ~n8016 & n8032;
  assign n8034 = x686 & ~n8010;
  assign n8035 = ~n8020 & ~n8034;
  assign n8036 = n8014 & ~n8035;
  assign n8037 = n8018 & ~n8034;
  assign n8038 = ~n8036 & ~n8037;
  assign n8039 = ~x685 & ~n8038;
  assign n8040 = ~n8033 & ~n8039;
  assign n7937 = x690 ^ x689;
  assign n7938 = n7937 ^ n7936;
  assign n7935 = x686 ^ x685;
  assign n7939 = n7938 ^ n7935;
  assign n8041 = ~x686 & n8022;
  assign n8042 = n7939 & n8041;
  assign n8043 = n8040 & ~n8042;
  assign n8044 = x681 & x682;
  assign n8045 = x683 & x684;
  assign n8046 = ~n8044 & ~n8045;
  assign n8047 = ~x681 & ~x682;
  assign n8048 = ~x683 & ~x684;
  assign n8049 = ~n8047 & ~n8048;
  assign n8050 = ~n8046 & n8049;
  assign n8051 = x680 & n8050;
  assign n8052 = n8044 & n8045;
  assign n8053 = ~n8051 & ~n8052;
  assign n8054 = n8046 & ~n8049;
  assign n8055 = ~x680 & n8054;
  assign n8056 = n8053 & ~n8055;
  assign n8057 = ~x679 & ~n8056;
  assign n7932 = x680 ^ x679;
  assign n8058 = n8047 & n8048;
  assign n8059 = n7932 & n8058;
  assign n8060 = n8050 ^ x680;
  assign n8061 = n8060 ^ n8050;
  assign n8062 = ~n8052 & ~n8054;
  assign n8063 = n8062 ^ n8050;
  assign n8064 = n8061 & n8063;
  assign n8065 = n8064 ^ n8050;
  assign n8066 = x679 & n8065;
  assign n8067 = ~n8059 & ~n8066;
  assign n8068 = ~n8057 & n8067;
  assign n10825 = n8043 & n8068;
  assign n10823 = ~n8033 & ~n8036;
  assign n10822 = n8053 & ~n8066;
  assign n10824 = n10823 ^ n10822;
  assign n10826 = n10825 ^ n10824;
  assign n10835 = n10834 ^ n10826;
  assign n8069 = n8068 ^ n8043;
  assign n7951 = n7950 ^ n7945;
  assign n8006 = n7951 ^ n7939;
  assign n7931 = x684 ^ x683;
  assign n7933 = n7932 ^ n7931;
  assign n7930 = x682 ^ x681;
  assign n7934 = n7933 ^ n7930;
  assign n8007 = n7951 ^ n7934;
  assign n8008 = n8006 & ~n8007;
  assign n8009 = n8008 ^ n7939;
  assign n8070 = n8069 ^ n8009;
  assign n8174 = n8173 ^ n8071;
  assign n10819 = n8174 ^ n8069;
  assign n10820 = ~n8070 & n10819;
  assign n10821 = n10820 ^ n8174;
  assign n10836 = n10835 ^ n10821;
  assign n11397 = ~n10822 & ~n10823;
  assign n11398 = ~n10836 & n11397;
  assign n11399 = n10824 & n10825;
  assign n11400 = n10821 & n11399;
  assign n11401 = ~n11398 & ~n11400;
  assign n11402 = n10834 & ~n11401;
  assign n11394 = n10832 ^ n10829;
  assign n11395 = ~n10833 & ~n11394;
  assign n11396 = n11395 ^ n10829;
  assign n11403 = ~n10821 & n10835;
  assign n11404 = n10823 & ~n11399;
  assign n11405 = n11403 & n11404;
  assign n11406 = n10822 & ~n10825;
  assign n11407 = ~n10834 & n11406;
  assign n11408 = ~n11405 & ~n11407;
  assign n11409 = n10821 & ~n10823;
  assign n11410 = ~n11408 & ~n11409;
  assign n11411 = ~n11402 & ~n11410;
  assign n11660 = n11396 & n11411;
  assign n11661 = ~n11402 & ~n11660;
  assign n11665 = n11664 ^ n11661;
  assign n11412 = n11411 ^ n11396;
  assign n7929 = n7928 ^ n7917;
  assign n7940 = n7939 ^ n7934;
  assign n7952 = n7951 ^ n7940;
  assign n8003 = n7929 & n7952;
  assign n8175 = n8174 ^ n8070;
  assign n8314 = n8313 ^ n8175;
  assign n10816 = n8003 & n8314;
  assign n10817 = n8175 & n8313;
  assign n10818 = ~n10816 & ~n10817;
  assign n10837 = n10836 ^ n10818;
  assign n10798 = n10797 ^ n10796;
  assign n10815 = n10814 ^ n10798;
  assign n11391 = n10818 ^ n10815;
  assign n11392 = ~n10837 & ~n11391;
  assign n11393 = n11392 ^ n10836;
  assign n11413 = n11412 ^ n11393;
  assign n11657 = n11433 ^ n11412;
  assign n11658 = ~n11413 & n11657;
  assign n11659 = n11658 ^ n11433;
  assign n11666 = n11665 ^ n11659;
  assign n7984 = x746 ^ x745;
  assign n7983 = x748 ^ x747;
  assign n8636 = x749 & x750;
  assign n8637 = n8636 ^ x748;
  assign n8638 = n7983 & ~n8637;
  assign n8639 = n8638 ^ x747;
  assign n8640 = n7984 & n8639;
  assign n8641 = ~x747 & ~x748;
  assign n8642 = ~n8636 & n8641;
  assign n8643 = x747 & x748;
  assign n8644 = x745 & x746;
  assign n8645 = ~n8643 & n8644;
  assign n8646 = ~n8642 & n8645;
  assign n8647 = ~n8640 & ~n8646;
  assign n8648 = ~x749 & ~x750;
  assign n8649 = ~n8647 & ~n8648;
  assign n8650 = n8643 & n8644;
  assign n8651 = ~x750 & n8650;
  assign n8652 = ~n8649 & ~n8651;
  assign n8653 = x746 & ~n8648;
  assign n8654 = n8636 & n8643;
  assign n8655 = ~n8653 & ~n8654;
  assign n8656 = n8639 & ~n8655;
  assign n10885 = n8652 & ~n8656;
  assign n8595 = x741 & x742;
  assign n8594 = x743 & x744;
  assign n8596 = n8595 ^ n8594;
  assign n8597 = ~x741 & ~x742;
  assign n8598 = ~x743 & ~x744;
  assign n8599 = ~n8597 & ~n8598;
  assign n8600 = n8599 ^ n8594;
  assign n8601 = n8600 ^ n8594;
  assign n8602 = n8594 ^ x740;
  assign n8603 = n8602 ^ n8594;
  assign n8604 = n8601 & n8603;
  assign n8605 = n8604 ^ n8594;
  assign n8606 = n8596 & ~n8605;
  assign n8607 = n8606 ^ n8595;
  assign n8609 = ~n8594 & ~n8595;
  assign n8622 = n8599 & ~n8609;
  assign n8621 = x744 & n8595;
  assign n8623 = n8622 ^ n8621;
  assign n8624 = n8623 ^ n8622;
  assign n8625 = ~n8599 & n8609;
  assign n8626 = n8625 ^ n8622;
  assign n8627 = n8626 ^ n8622;
  assign n8628 = ~n8624 & ~n8627;
  assign n8629 = n8628 ^ n8622;
  assign n8630 = x740 & n8629;
  assign n8631 = n8630 ^ n8622;
  assign n10883 = x739 & n8631;
  assign n10884 = ~n8607 & ~n10883;
  assign n10886 = n10885 ^ n10884;
  assign n8657 = n8648 ^ n8642;
  assign n8658 = n8648 ^ n8643;
  assign n8659 = n8642 ^ x746;
  assign n8660 = n8659 ^ n8648;
  assign n8661 = n8648 & ~n8660;
  assign n8662 = n8661 ^ n8648;
  assign n8663 = n8658 & n8662;
  assign n8664 = n8663 ^ n8661;
  assign n8665 = n8664 ^ n8648;
  assign n8666 = n8665 ^ n8659;
  assign n8667 = n8657 & ~n8666;
  assign n8668 = n8667 ^ n8642;
  assign n8669 = ~n8656 & ~n8668;
  assign n8670 = ~x745 & ~n8669;
  assign n8671 = n8652 & ~n8670;
  assign n8672 = ~x746 & ~x750;
  assign n8673 = n8641 & n8672;
  assign n8674 = ~n8650 & ~n8673;
  assign n8675 = ~x749 & ~n8674;
  assign n8676 = n8671 & ~n8675;
  assign n7979 = x742 ^ x741;
  assign n8585 = x739 & x740;
  assign n8586 = n8585 ^ x742;
  assign n8587 = n8586 ^ n8585;
  assign n8588 = ~x740 & ~x744;
  assign n8589 = n8588 ^ n8585;
  assign n8590 = ~n8587 & n8589;
  assign n8591 = n8590 ^ n8585;
  assign n8592 = ~n7979 & n8591;
  assign n8593 = ~x743 & n8592;
  assign n8608 = n8598 ^ n8597;
  assign n8610 = n8609 ^ n8598;
  assign n8611 = n8610 ^ n8598;
  assign n8612 = n8598 ^ x740;
  assign n8613 = n8612 ^ n8598;
  assign n8614 = n8611 & ~n8613;
  assign n8615 = n8614 ^ n8598;
  assign n8616 = n8608 & ~n8615;
  assign n8617 = n8616 ^ n8597;
  assign n8618 = ~n8607 & ~n8617;
  assign n8619 = n8618 ^ x739;
  assign n8620 = n8619 ^ n8618;
  assign n8632 = n8631 ^ n8618;
  assign n8633 = n8620 & ~n8632;
  assign n8634 = n8633 ^ n8618;
  assign n8635 = ~n8593 & n8634;
  assign n8677 = n8676 ^ n8635;
  assign n7978 = x744 ^ x743;
  assign n7980 = n7979 ^ n7978;
  assign n7977 = x740 ^ x739;
  assign n7981 = n7980 ^ n7977;
  assign n7985 = n7984 ^ n7983;
  assign n7982 = x750 ^ x749;
  assign n7986 = n7985 ^ n7982;
  assign n8498 = n7981 & n7986;
  assign n10880 = n8635 ^ n8498;
  assign n10881 = n8677 & ~n10880;
  assign n10882 = n10881 ^ n8676;
  assign n10887 = n10886 ^ n10882;
  assign n8508 = x731 & x732;
  assign n8507 = x729 & x730;
  assign n8509 = n8508 ^ n8507;
  assign n8510 = ~x731 & ~x732;
  assign n8511 = ~x729 & ~x730;
  assign n8512 = ~n8510 & ~n8511;
  assign n8513 = n8512 ^ n8507;
  assign n8514 = n8513 ^ n8507;
  assign n8515 = n8507 ^ x728;
  assign n8516 = n8515 ^ n8507;
  assign n8517 = n8514 & n8516;
  assign n8518 = n8517 ^ n8507;
  assign n8519 = n8509 & ~n8518;
  assign n8520 = n8519 ^ n8508;
  assign n7995 = x732 ^ x731;
  assign n7994 = x730 ^ x729;
  assign n7996 = n7995 ^ n7994;
  assign n7993 = x728 ^ x727;
  assign n7997 = n7996 ^ n7993;
  assign n8506 = x727 & ~n7997;
  assign n8522 = ~n8507 & ~n8508;
  assign n8535 = ~n8512 & n8522;
  assign n10878 = n8506 & ~n8535;
  assign n10879 = ~n8520 & ~n10878;
  assign n10888 = n10887 ^ n10879;
  assign n8543 = x737 & x738;
  assign n8542 = x735 & x736;
  assign n8544 = n8543 ^ n8542;
  assign n8545 = ~x737 & ~x738;
  assign n8546 = ~x735 & ~x736;
  assign n8547 = ~n8545 & ~n8546;
  assign n8548 = n8547 ^ n8542;
  assign n8549 = n8548 ^ n8542;
  assign n8550 = n8542 ^ x734;
  assign n8551 = n8550 ^ n8542;
  assign n8552 = n8549 & n8551;
  assign n8553 = n8552 ^ n8542;
  assign n8554 = n8544 & ~n8553;
  assign n8555 = n8554 ^ n8543;
  assign n7988 = x738 ^ x737;
  assign n8556 = x737 ^ x734;
  assign n8557 = n7988 & n8556;
  assign n8558 = n8557 ^ x737;
  assign n8559 = n8546 & ~n8558;
  assign n8560 = ~n8555 & ~n8559;
  assign n8561 = ~x733 & ~n8560;
  assign n7990 = x734 ^ x733;
  assign n8562 = ~n8542 & ~n8543;
  assign n8563 = n8547 & ~n8562;
  assign n8564 = n7990 & n8563;
  assign n8565 = ~n8547 & n8562;
  assign n8566 = x733 & x734;
  assign n8567 = x738 & n8542;
  assign n8568 = n8566 & ~n8567;
  assign n8569 = ~n8565 & n8568;
  assign n8570 = ~n8564 & ~n8569;
  assign n8571 = ~x737 & n8566;
  assign n7989 = x736 ^ x735;
  assign n7991 = n7990 ^ n7989;
  assign n8572 = n8571 ^ n7991;
  assign n8573 = n8572 ^ n8571;
  assign n8574 = ~x734 & n8545;
  assign n8575 = n8574 ^ n8571;
  assign n8576 = n8575 ^ n8571;
  assign n8577 = n8573 & n8576;
  assign n8578 = n8577 ^ n8571;
  assign n8579 = ~n8542 & n8578;
  assign n8580 = n8579 ^ n8571;
  assign n8581 = n8570 & ~n8580;
  assign n8582 = ~n8561 & n8581;
  assign n8532 = n8507 & n8508;
  assign n8521 = n8511 ^ n8510;
  assign n8523 = n8522 ^ n8511;
  assign n8524 = n8523 ^ n8511;
  assign n8525 = n8511 ^ x728;
  assign n8526 = n8525 ^ n8511;
  assign n8527 = n8524 & ~n8526;
  assign n8528 = n8527 ^ n8511;
  assign n8529 = n8521 & ~n8528;
  assign n8530 = n8529 ^ n8510;
  assign n8531 = ~n8520 & ~n8530;
  assign n8533 = n8532 ^ n8531;
  assign n8534 = n8533 ^ n8531;
  assign n8536 = n8535 ^ n8531;
  assign n8537 = n8536 ^ n8531;
  assign n8538 = ~n8534 & ~n8537;
  assign n8539 = n8538 ^ n8531;
  assign n8540 = n8506 & ~n8539;
  assign n8541 = n8540 ^ n8531;
  assign n8583 = n8582 ^ n8541;
  assign n7992 = n7991 ^ n7988;
  assign n8502 = n7992 & n7997;
  assign n7998 = n7997 ^ n7992;
  assign n7987 = n7986 ^ n7981;
  assign n8499 = n7992 ^ n7987;
  assign n8500 = n7998 & ~n8499;
  assign n8501 = n8500 ^ n7997;
  assign n8503 = n8502 ^ n8501;
  assign n8504 = ~n8498 & ~n8503;
  assign n8505 = n8504 ^ n8502;
  assign n8584 = n8583 ^ n8505;
  assign n8678 = n8677 ^ n8584;
  assign n10872 = ~n8498 & n8677;
  assign n10873 = ~n8678 & ~n10872;
  assign n10874 = ~n8503 & ~n8583;
  assign n10875 = n10874 ^ n8502;
  assign n10876 = ~n10873 & ~n10875;
  assign n10867 = ~n8555 & n8570;
  assign n10868 = ~n8502 & n8583;
  assign n10869 = ~n8541 & ~n8582;
  assign n10870 = ~n10868 & ~n10869;
  assign n11446 = n10867 & ~n10870;
  assign n11447 = ~n10876 & n11446;
  assign n11448 = n11447 ^ n10879;
  assign n11449 = n11448 ^ n11447;
  assign n10871 = n10870 ^ n10867;
  assign n11441 = n10876 ^ n10870;
  assign n11442 = n10871 & n11441;
  assign n11443 = n11442 ^ n10876;
  assign n11450 = n11447 ^ n11443;
  assign n11451 = n11450 ^ n11447;
  assign n11452 = n11449 & ~n11451;
  assign n11453 = n11452 ^ n11447;
  assign n11454 = n10888 & n11453;
  assign n11455 = n11454 ^ n11447;
  assign n11438 = n10885 ^ n10882;
  assign n11439 = ~n10886 & ~n11438;
  assign n11440 = n11439 ^ n10882;
  assign n10877 = n10876 ^ n10871;
  assign n10889 = n10888 ^ n10877;
  assign n11444 = n10887 & n11443;
  assign n11445 = ~n10889 & n11444;
  assign n11653 = ~n11440 & ~n11445;
  assign n11654 = ~n11455 & ~n11653;
  assign n8360 = x705 & x706;
  assign n8359 = x707 & x708;
  assign n8361 = n8360 ^ n8359;
  assign n8362 = ~x705 & ~x706;
  assign n8363 = ~x707 & ~x708;
  assign n8364 = ~n8362 & ~n8363;
  assign n8365 = n8364 ^ n8359;
  assign n8366 = n8365 ^ n8359;
  assign n8367 = n8359 ^ x704;
  assign n8368 = n8367 ^ n8359;
  assign n8369 = n8366 & n8368;
  assign n8370 = n8369 ^ n8359;
  assign n8371 = n8361 & ~n8370;
  assign n8372 = n8371 ^ n8360;
  assign n8390 = ~n8359 & ~n8360;
  assign n8391 = ~n8364 & n8390;
  assign n8379 = x703 & x704;
  assign n8392 = n8360 & n8379;
  assign n8393 = x708 & n8392;
  assign n8394 = n8393 ^ n8379;
  assign n8395 = ~n8391 & n8394;
  assign n7972 = x704 ^ x703;
  assign n8396 = n8364 & ~n8390;
  assign n8397 = n7972 & n8396;
  assign n8398 = ~n8395 & ~n8397;
  assign n10843 = ~n8372 & n8398;
  assign n8318 = x711 & x712;
  assign n8317 = x713 & x714;
  assign n8319 = n8318 ^ n8317;
  assign n8320 = ~x711 & ~x712;
  assign n8321 = ~x713 & ~x714;
  assign n8322 = ~n8320 & ~n8321;
  assign n8323 = n8322 ^ n8317;
  assign n8324 = n8323 ^ n8317;
  assign n8325 = n8317 ^ x710;
  assign n8326 = n8325 ^ n8317;
  assign n8327 = n8324 & n8326;
  assign n8328 = n8327 ^ n8317;
  assign n8329 = n8319 & ~n8328;
  assign n8330 = n8329 ^ n8318;
  assign n8348 = ~n8317 & ~n8318;
  assign n8349 = ~n8322 & n8348;
  assign n8337 = x709 & x710;
  assign n8350 = n8318 & n8337;
  assign n8351 = x714 & n8350;
  assign n8352 = n8351 ^ n8337;
  assign n8353 = ~n8349 & n8352;
  assign n7967 = x710 ^ x709;
  assign n8354 = n8322 & ~n8348;
  assign n8355 = n7967 & n8354;
  assign n8356 = ~n8353 & ~n8355;
  assign n10842 = ~n8330 & n8356;
  assign n10844 = n10843 ^ n10842;
  assign n7970 = x708 ^ x707;
  assign n8373 = x707 ^ x704;
  assign n8374 = n7970 & n8373;
  assign n8375 = n8374 ^ x707;
  assign n8376 = n8362 & ~n8375;
  assign n8377 = ~n8372 & ~n8376;
  assign n8378 = ~x703 & ~n8377;
  assign n7971 = x706 ^ x705;
  assign n7973 = n7972 ^ n7971;
  assign n8380 = n8379 ^ n7973;
  assign n8381 = n8380 ^ n8379;
  assign n8382 = ~x704 & ~x708;
  assign n8383 = n8382 ^ n8379;
  assign n8384 = n8383 ^ n8379;
  assign n8385 = n8381 & n8384;
  assign n8386 = n8385 ^ n8379;
  assign n8387 = ~n8360 & n8386;
  assign n8388 = n8387 ^ n8379;
  assign n8389 = ~x707 & n8388;
  assign n8399 = ~n8389 & n8398;
  assign n8400 = ~n8378 & n8399;
  assign n7965 = x714 ^ x713;
  assign n8331 = x713 ^ x710;
  assign n8332 = n7965 & n8331;
  assign n8333 = n8332 ^ x713;
  assign n8334 = n8320 & ~n8333;
  assign n8335 = ~n8330 & ~n8334;
  assign n8336 = ~x709 & ~n8335;
  assign n7966 = x712 ^ x711;
  assign n7968 = n7967 ^ n7966;
  assign n8338 = n8337 ^ n7968;
  assign n8339 = n8338 ^ n8337;
  assign n8340 = ~x710 & ~x714;
  assign n8341 = n8340 ^ n8337;
  assign n8342 = n8341 ^ n8337;
  assign n8343 = n8339 & n8342;
  assign n8344 = n8343 ^ n8337;
  assign n8345 = ~n8318 & n8344;
  assign n8346 = n8345 ^ n8337;
  assign n8347 = ~x713 & n8346;
  assign n8357 = ~n8347 & n8356;
  assign n8358 = ~n8336 & n8357;
  assign n8401 = n8400 ^ n8358;
  assign n7969 = n7968 ^ n7965;
  assign n7974 = n7973 ^ n7970;
  assign n8402 = n7969 & n7974;
  assign n10845 = n8401 & n8402;
  assign n10846 = n8358 & n8400;
  assign n10847 = ~n10845 & ~n10846;
  assign n11464 = n10847 ^ n10843;
  assign n11465 = ~n10844 & n11464;
  assign n11466 = n11465 ^ n10847;
  assign n7956 = x716 ^ x715;
  assign n7955 = x718 ^ x717;
  assign n7957 = n7956 ^ n7955;
  assign n7954 = x720 ^ x719;
  assign n7958 = n7957 ^ n7954;
  assign n7961 = x722 ^ x721;
  assign n7960 = x724 ^ x723;
  assign n7962 = n7961 ^ n7960;
  assign n7959 = x726 ^ x725;
  assign n7963 = n7962 ^ n7959;
  assign n8403 = n7958 & n7963;
  assign n8453 = x723 & x724;
  assign n8452 = x725 & x726;
  assign n8454 = n8453 ^ n8452;
  assign n8455 = ~x723 & ~x724;
  assign n8456 = ~x725 & ~x726;
  assign n8457 = ~n8455 & ~n8456;
  assign n8458 = n8457 ^ n8452;
  assign n8459 = n8458 ^ n8452;
  assign n8460 = n8452 ^ x722;
  assign n8461 = n8460 ^ n8452;
  assign n8462 = n8459 & n8461;
  assign n8463 = n8462 ^ n8452;
  assign n8464 = n8454 & ~n8463;
  assign n8465 = n8464 ^ n8453;
  assign n8466 = x725 ^ x722;
  assign n8467 = n7959 & n8466;
  assign n8468 = n8467 ^ x725;
  assign n8469 = n8455 & ~n8468;
  assign n8470 = ~n8465 & ~n8469;
  assign n8471 = ~x721 & ~n8470;
  assign n8472 = x721 & x722;
  assign n8473 = n8472 ^ n7962;
  assign n8474 = n8473 ^ n8472;
  assign n8475 = ~x722 & ~x726;
  assign n8476 = n8475 ^ n8472;
  assign n8477 = n8476 ^ n8472;
  assign n8478 = n8474 & n8477;
  assign n8479 = n8478 ^ n8472;
  assign n8480 = ~n8453 & n8479;
  assign n8481 = n8480 ^ n8472;
  assign n8482 = ~x725 & n8481;
  assign n8483 = ~n8452 & ~n8453;
  assign n8484 = ~n8457 & n8483;
  assign n8485 = n8453 & n8472;
  assign n8486 = x726 & n8485;
  assign n8487 = n8486 ^ n8472;
  assign n8488 = ~n8484 & n8487;
  assign n8489 = n8457 & ~n8483;
  assign n8490 = n7961 & n8489;
  assign n8491 = ~n8488 & ~n8490;
  assign n8492 = ~n8482 & n8491;
  assign n8493 = ~n8471 & n8492;
  assign n8411 = x717 & x718;
  assign n8410 = x719 & x720;
  assign n8412 = n8411 ^ n8410;
  assign n8413 = ~x717 & ~x718;
  assign n8414 = ~x719 & ~x720;
  assign n8415 = ~n8413 & ~n8414;
  assign n8416 = n8415 ^ n8410;
  assign n8417 = n8416 ^ n8410;
  assign n8418 = n8410 ^ x716;
  assign n8419 = n8418 ^ n8410;
  assign n8420 = n8417 & n8419;
  assign n8421 = n8420 ^ n8410;
  assign n8422 = n8412 & ~n8421;
  assign n8423 = n8422 ^ n8411;
  assign n8424 = x719 ^ x716;
  assign n8425 = n7954 & n8424;
  assign n8426 = n8425 ^ x719;
  assign n8427 = n8413 & ~n8426;
  assign n8428 = ~n8423 & ~n8427;
  assign n8429 = ~x715 & ~n8428;
  assign n8430 = x715 & x716;
  assign n8431 = n8430 ^ n7957;
  assign n8432 = n8431 ^ n8430;
  assign n8433 = ~x716 & ~x720;
  assign n8434 = n8433 ^ n8430;
  assign n8435 = n8434 ^ n8430;
  assign n8436 = n8432 & n8435;
  assign n8437 = n8436 ^ n8430;
  assign n8438 = ~n8411 & n8437;
  assign n8439 = n8438 ^ n8430;
  assign n8440 = ~x719 & n8439;
  assign n8441 = ~n8410 & ~n8411;
  assign n8442 = ~n8415 & n8441;
  assign n8443 = n8411 & n8430;
  assign n8444 = x720 & n8443;
  assign n8445 = n8444 ^ n8430;
  assign n8446 = ~n8442 & n8445;
  assign n8447 = n8415 & ~n8441;
  assign n8448 = n7956 & n8447;
  assign n8449 = ~n8446 & ~n8448;
  assign n8450 = ~n8440 & n8449;
  assign n8451 = ~n8429 & n8450;
  assign n8494 = n8493 ^ n8451;
  assign n10860 = n8403 & n8494;
  assign n10861 = n8451 & n8493;
  assign n10862 = ~n10860 & ~n10861;
  assign n10858 = ~n8465 & n8491;
  assign n10857 = ~n8423 & n8449;
  assign n10859 = n10858 ^ n10857;
  assign n10863 = n10862 ^ n10859;
  assign n7975 = n7974 ^ n7969;
  assign n7964 = n7963 ^ n7958;
  assign n8405 = n7969 ^ n7964;
  assign n8406 = n7975 & n8405;
  assign n8407 = n8406 ^ n7969;
  assign n8408 = ~n8403 & ~n8407;
  assign n10849 = n8408 ^ n8403;
  assign n10850 = ~n8494 & n10849;
  assign n10851 = n10850 ^ n8403;
  assign n8404 = n8402 & n8403;
  assign n8409 = ~n8404 & ~n8408;
  assign n8495 = n8494 ^ n8409;
  assign n8496 = n8495 ^ n8401;
  assign n10852 = n8496 ^ n8495;
  assign n10853 = n8495 ^ n8402;
  assign n10854 = n10852 & n10853;
  assign n10855 = n10854 ^ n8495;
  assign n10856 = ~n10851 & ~n10855;
  assign n10864 = n10863 ^ n10856;
  assign n10848 = n10847 ^ n10844;
  assign n11469 = n10863 ^ n10848;
  assign n11470 = ~n10864 & n11469;
  assign n11471 = n11470 ^ n10863;
  assign n11472 = n11466 & n11471;
  assign n11461 = n10862 ^ n10858;
  assign n11462 = ~n10859 & n11461;
  assign n11463 = n11462 ^ n10862;
  assign n10865 = n10864 ^ n10848;
  assign n11467 = ~n10863 & ~n11466;
  assign n11468 = ~n10865 & n11467;
  assign n11473 = ~n11468 & ~n11472;
  assign n11651 = n11463 & n11473;
  assign n11652 = ~n11472 & ~n11651;
  assign n11655 = n11654 ^ n11652;
  assign n11474 = n11473 ^ n11463;
  assign n7976 = n7975 ^ n7964;
  assign n7999 = n7998 ^ n7987;
  assign n8316 = n7976 & n7999;
  assign n8497 = n8496 ^ n8316;
  assign n10839 = n8678 ^ n8316;
  assign n10840 = n8497 & n10839;
  assign n10841 = n10840 ^ n8496;
  assign n10866 = n10865 ^ n10841;
  assign n11458 = n10889 ^ n10841;
  assign n11459 = n10866 & ~n11458;
  assign n11460 = n11459 ^ n10865;
  assign n11475 = n11474 ^ n11460;
  assign n11456 = ~n11445 & ~n11455;
  assign n11457 = n11456 ^ n11440;
  assign n11648 = n11460 ^ n11457;
  assign n11649 = ~n11475 & ~n11648;
  assign n11650 = n11649 ^ n11474;
  assign n11656 = n11655 ^ n11650;
  assign n11667 = n11666 ^ n11656;
  assign n11476 = n11475 ^ n11457;
  assign n10890 = n10889 ^ n10866;
  assign n10838 = n10837 ^ n10815;
  assign n10891 = n10890 ^ n10838;
  assign n10782 = n8314 ^ n8003;
  assign n8679 = n8678 ^ n8497;
  assign n10783 = n10782 ^ n8679;
  assign n10784 = n8679 ^ n8003;
  assign n10785 = n10784 ^ n8679;
  assign n7953 = n7952 ^ n7929;
  assign n8000 = n7999 ^ n7976;
  assign n8004 = n7953 & n8000;
  assign n10786 = n8679 ^ n8004;
  assign n10787 = n10786 ^ n8679;
  assign n10788 = ~n10785 & n10787;
  assign n10789 = n10788 ^ n8679;
  assign n10790 = ~n10783 & ~n10789;
  assign n10791 = n10790 ^ n8679;
  assign n11435 = n10838 ^ n10791;
  assign n11436 = n10891 & n11435;
  assign n11437 = n11436 ^ n10890;
  assign n11477 = n11476 ^ n11437;
  assign n11434 = n11433 ^ n11413;
  assign n11645 = n11437 ^ n11434;
  assign n11646 = ~n11477 & ~n11645;
  assign n11647 = n11646 ^ n11476;
  assign n11701 = n11656 ^ n11647;
  assign n11702 = n11667 & ~n11701;
  assign n11703 = n11702 ^ n11666;
  assign n11707 = n11654 ^ n11650;
  assign n11708 = ~n11655 & ~n11707;
  assign n11709 = n11708 ^ n11650;
  assign n11806 = n11703 & n11709;
  assign n8737 = x789 & x790;
  assign n8736 = x791 & x792;
  assign n8738 = n8737 ^ n8736;
  assign n8739 = ~x789 & ~x790;
  assign n8740 = ~x791 & ~x792;
  assign n8741 = ~n8739 & ~n8740;
  assign n8742 = n8741 ^ n8736;
  assign n8743 = n8742 ^ n8736;
  assign n8744 = n8736 ^ x788;
  assign n8745 = n8744 ^ n8736;
  assign n8746 = n8743 & n8745;
  assign n8747 = n8746 ^ n8736;
  assign n8748 = n8738 & ~n8747;
  assign n8749 = n8748 ^ n8737;
  assign n7884 = x788 ^ x787;
  assign n8751 = ~n8736 & ~n8737;
  assign n8762 = n8741 & ~n8751;
  assign n8763 = n7884 & n8762;
  assign n8764 = ~n8741 & n8751;
  assign n8765 = x787 & x788;
  assign n8766 = n8737 & n8765;
  assign n8767 = x792 & n8766;
  assign n8768 = n8767 ^ n8765;
  assign n8769 = ~n8764 & n8768;
  assign n8770 = ~n8763 & ~n8769;
  assign n10694 = ~n8749 & n8770;
  assign n8692 = x795 & x796;
  assign n8691 = x797 & x798;
  assign n8693 = n8692 ^ n8691;
  assign n8694 = ~x795 & ~x796;
  assign n8695 = ~x797 & ~x798;
  assign n8696 = ~n8694 & ~n8695;
  assign n8697 = n8696 ^ n8691;
  assign n8698 = n8697 ^ n8691;
  assign n8699 = n8691 ^ x794;
  assign n8700 = n8699 ^ n8691;
  assign n8701 = n8698 & n8700;
  assign n8702 = n8701 ^ n8691;
  assign n8703 = n8693 & ~n8702;
  assign n8704 = n8703 ^ n8692;
  assign n7889 = x794 ^ x793;
  assign n8706 = ~n8691 & ~n8692;
  assign n8717 = n8696 & ~n8706;
  assign n8718 = n7889 & n8717;
  assign n8719 = ~n8696 & n8706;
  assign n8720 = x793 & x794;
  assign n8721 = n8692 & n8720;
  assign n8722 = x798 & n8721;
  assign n8723 = n8722 ^ n8720;
  assign n8724 = ~n8719 & n8723;
  assign n8725 = ~n8718 & ~n8724;
  assign n10693 = ~n8704 & n8725;
  assign n10695 = n10694 ^ n10693;
  assign n7883 = x790 ^ x789;
  assign n7885 = n7884 ^ n7883;
  assign n7882 = x792 ^ x791;
  assign n7886 = n7885 ^ n7882;
  assign n7888 = x796 ^ x795;
  assign n7890 = n7889 ^ n7888;
  assign n7887 = x798 ^ x797;
  assign n7891 = n7890 ^ n7887;
  assign n8690 = n7886 & n7891;
  assign n8750 = n8740 ^ n8739;
  assign n8752 = n8751 ^ n8740;
  assign n8753 = n8752 ^ n8740;
  assign n8754 = n8740 ^ x788;
  assign n8755 = n8754 ^ n8740;
  assign n8756 = n8753 & ~n8755;
  assign n8757 = n8756 ^ n8740;
  assign n8758 = n8750 & ~n8757;
  assign n8759 = n8758 ^ n8739;
  assign n8760 = ~n8749 & ~n8759;
  assign n8761 = ~x787 & ~n8760;
  assign n8771 = n8765 ^ x790;
  assign n8772 = n8771 ^ n8765;
  assign n8773 = ~x788 & ~x792;
  assign n8774 = n8773 ^ n8765;
  assign n8775 = ~n8772 & n8774;
  assign n8776 = n8775 ^ n8765;
  assign n8777 = ~n7883 & n8776;
  assign n8778 = ~x791 & n8777;
  assign n8779 = n8770 & ~n8778;
  assign n8780 = ~n8761 & n8779;
  assign n8705 = n8695 ^ n8694;
  assign n8707 = n8706 ^ n8695;
  assign n8708 = n8707 ^ n8695;
  assign n8709 = n8695 ^ x794;
  assign n8710 = n8709 ^ n8695;
  assign n8711 = n8708 & ~n8710;
  assign n8712 = n8711 ^ n8695;
  assign n8713 = n8705 & ~n8712;
  assign n8714 = n8713 ^ n8694;
  assign n8715 = ~n8704 & ~n8714;
  assign n8716 = ~x793 & ~n8715;
  assign n8726 = n8720 ^ x796;
  assign n8727 = n8726 ^ n8720;
  assign n8728 = ~x794 & ~x798;
  assign n8729 = n8728 ^ n8720;
  assign n8730 = ~n8727 & n8729;
  assign n8731 = n8730 ^ n8720;
  assign n8732 = ~n7888 & n8731;
  assign n8733 = ~x797 & n8732;
  assign n8734 = n8725 & ~n8733;
  assign n8735 = ~n8716 & n8734;
  assign n8781 = n8780 ^ n8735;
  assign n10696 = ~n8690 & n8781;
  assign n10697 = ~n8735 & ~n8780;
  assign n10698 = ~n10696 & ~n10697;
  assign n11549 = n10698 ^ n10694;
  assign n11550 = ~n10695 & ~n11549;
  assign n11551 = n11550 ^ n10698;
  assign n10699 = n10698 ^ n10695;
  assign n8828 = x779 & x780;
  assign n8829 = x777 & x778;
  assign n8830 = ~n8828 & ~n8829;
  assign n8831 = ~x779 & ~x780;
  assign n8832 = ~x777 & ~x778;
  assign n8833 = ~n8831 & ~n8832;
  assign n8834 = ~n8830 & n8833;
  assign n8835 = x776 & n8834;
  assign n8836 = n8828 & n8829;
  assign n8837 = ~n8835 & ~n8836;
  assign n8838 = n8830 & ~n8833;
  assign n8839 = ~x776 & n8838;
  assign n8840 = n8837 & ~n8839;
  assign n8841 = ~x775 & ~n8840;
  assign n7895 = x776 ^ x775;
  assign n8842 = n8831 & n8832;
  assign n8843 = n7895 & n8842;
  assign n8844 = n8834 ^ x776;
  assign n8845 = n8844 ^ n8834;
  assign n8846 = ~n8836 & ~n8838;
  assign n8847 = n8846 ^ n8834;
  assign n8848 = n8845 & n8847;
  assign n8849 = n8848 ^ n8834;
  assign n8850 = x775 & n8849;
  assign n8851 = ~n8843 & ~n8850;
  assign n8852 = ~n8841 & n8851;
  assign n8784 = x785 & x786;
  assign n8783 = x783 & x784;
  assign n8785 = n8784 ^ n8783;
  assign n8786 = ~x785 & ~x786;
  assign n8787 = ~x783 & ~x784;
  assign n8788 = ~n8786 & ~n8787;
  assign n8789 = n8788 ^ n8783;
  assign n8790 = n8789 ^ n8783;
  assign n8791 = n8783 ^ x782;
  assign n8792 = n8791 ^ n8783;
  assign n8793 = n8790 & n8792;
  assign n8794 = n8793 ^ n8783;
  assign n8795 = n8785 & ~n8794;
  assign n8796 = n8795 ^ n8784;
  assign n8797 = n8787 ^ n8786;
  assign n8798 = ~n8783 & ~n8784;
  assign n8799 = n8798 ^ n8787;
  assign n8800 = n8799 ^ n8787;
  assign n8801 = n8787 ^ x782;
  assign n8802 = n8801 ^ n8787;
  assign n8803 = n8800 & ~n8802;
  assign n8804 = n8803 ^ n8787;
  assign n8805 = n8797 & ~n8804;
  assign n8806 = n8805 ^ n8786;
  assign n8807 = ~n8796 & ~n8806;
  assign n8808 = ~x781 & ~n8807;
  assign n7900 = x782 ^ x781;
  assign n8809 = n8788 & ~n8798;
  assign n8810 = n7900 & n8809;
  assign n8811 = ~n8788 & n8798;
  assign n8812 = x781 & x782;
  assign n8813 = n8783 & n8812;
  assign n8814 = x786 & n8813;
  assign n8815 = n8814 ^ n8812;
  assign n8816 = ~n8811 & n8815;
  assign n8817 = ~n8810 & ~n8816;
  assign n7899 = x784 ^ x783;
  assign n8818 = n8812 ^ x784;
  assign n8819 = n8818 ^ n8812;
  assign n8820 = ~x782 & ~x786;
  assign n8821 = n8820 ^ n8812;
  assign n8822 = ~n8819 & n8821;
  assign n8823 = n8822 ^ n8812;
  assign n8824 = ~n7899 & n8823;
  assign n8825 = ~x785 & n8824;
  assign n8826 = n8817 & ~n8825;
  assign n8827 = ~n8808 & n8826;
  assign n8853 = n8852 ^ n8827;
  assign n7894 = x778 ^ x777;
  assign n7896 = n7895 ^ n7894;
  assign n7893 = x780 ^ x779;
  assign n7897 = n7896 ^ n7893;
  assign n7901 = n7900 ^ n7899;
  assign n7898 = x786 ^ x785;
  assign n7902 = n7901 ^ n7898;
  assign n10701 = ~n7897 & ~n7902;
  assign n8686 = n7897 & n7902;
  assign n10702 = n10701 ^ n8686;
  assign n10703 = n8853 & n10702;
  assign n10704 = n10703 ^ n10701;
  assign n10709 = ~n8686 & ~n8853;
  assign n10710 = n8781 & ~n10709;
  assign n7903 = n7902 ^ n7897;
  assign n7892 = n7891 ^ n7886;
  assign n7904 = n7903 ^ n7892;
  assign n10711 = ~n7886 & n7904;
  assign n10712 = ~n10710 & n10711;
  assign n10713 = n10709 ^ n8690;
  assign n10714 = n10713 ^ n8690;
  assign n10715 = ~n7891 & ~n7903;
  assign n10716 = n10715 ^ n8690;
  assign n10717 = n10716 ^ n8690;
  assign n10718 = ~n10714 & ~n10717;
  assign n10719 = n10718 ^ n8690;
  assign n10720 = ~n8781 & ~n10719;
  assign n10721 = n10720 ^ n8690;
  assign n10722 = ~n10712 & ~n10721;
  assign n10723 = ~n10704 & n10722;
  assign n10705 = ~n8852 & ~n10704;
  assign n10706 = ~n8686 & ~n8827;
  assign n10707 = ~n10705 & ~n10706;
  assign n10690 = ~n8796 & n8817;
  assign n10691 = n8837 & ~n8850;
  assign n11552 = ~n10690 & ~n10691;
  assign n11553 = n10707 & n11552;
  assign n11554 = ~n10723 & ~n11553;
  assign n11555 = n10699 & ~n11554;
  assign n11556 = ~n10707 & ~n11552;
  assign n11557 = n11555 & ~n11556;
  assign n11558 = ~n11551 & ~n11557;
  assign n10692 = n10691 ^ n10690;
  assign n10700 = n10699 ^ n10692;
  assign n10708 = n10707 ^ n10700;
  assign n10724 = n10723 ^ n10708;
  assign n11559 = n10690 & n10691;
  assign n11560 = n10724 & n11559;
  assign n11561 = ~n11558 & ~n11560;
  assign n11563 = ~n10699 & n11556;
  assign n11564 = ~n11560 & ~n11563;
  assign n11565 = ~n10723 & ~n11564;
  assign n11692 = n11561 & ~n11565;
  assign n8953 = x767 & x768;
  assign n8954 = x765 & x766;
  assign n8955 = ~n8953 & ~n8954;
  assign n8956 = ~x767 & ~x768;
  assign n8957 = ~x765 & ~x766;
  assign n8958 = ~n8956 & ~n8957;
  assign n8959 = n8955 & ~n8958;
  assign n8960 = x763 & x764;
  assign n8961 = n8954 & n8960;
  assign n8962 = x768 & n8961;
  assign n8963 = n8962 ^ n8960;
  assign n8964 = ~n8959 & n8963;
  assign n8965 = ~n8955 & n8958;
  assign n8966 = ~x764 & n8965;
  assign n8967 = ~x763 & n8966;
  assign n8968 = n8967 ^ n8965;
  assign n8969 = ~n8964 & ~n8968;
  assign n8970 = n8953 & n8954;
  assign n8971 = n8969 & ~n8970;
  assign n7859 = x768 ^ x767;
  assign n8972 = x767 ^ x764;
  assign n8973 = n7859 & n8972;
  assign n8974 = n8973 ^ x767;
  assign n8975 = n8957 & ~n8974;
  assign n8976 = n8971 & ~n8975;
  assign n8977 = x763 & ~n8964;
  assign n8978 = ~n8966 & n8977;
  assign n8979 = ~n8976 & ~n8978;
  assign n8980 = ~x764 & ~x768;
  assign n8981 = n8980 ^ n8960;
  assign n8982 = n8981 ^ n8960;
  assign n7861 = x764 ^ x763;
  assign n7860 = x766 ^ x765;
  assign n7862 = n7861 ^ n7860;
  assign n8983 = n8960 ^ n7862;
  assign n8984 = n8983 ^ n8960;
  assign n8985 = n8982 & n8984;
  assign n8986 = n8985 ^ n8960;
  assign n8987 = ~n8954 & n8986;
  assign n8988 = n8987 ^ n8960;
  assign n8989 = ~x767 & n8988;
  assign n8990 = ~n8979 & ~n8989;
  assign n8928 = x773 & x774;
  assign n8929 = x771 & x772;
  assign n8930 = ~n8928 & ~n8929;
  assign n8931 = ~x773 & ~x774;
  assign n8932 = ~x771 & ~x772;
  assign n8933 = ~n8931 & ~n8932;
  assign n8934 = ~n8930 & n8933;
  assign n8935 = x770 & n8934;
  assign n8936 = n8928 & n8929;
  assign n8937 = ~n8935 & ~n8936;
  assign n8938 = n8930 & ~n8933;
  assign n8939 = ~x770 & n8938;
  assign n8940 = n8937 & ~n8939;
  assign n8941 = ~x769 & ~n8940;
  assign n7866 = x770 ^ x769;
  assign n8942 = n8931 & n8932;
  assign n8943 = n7866 & n8942;
  assign n8944 = n8934 ^ x770;
  assign n8945 = n8944 ^ n8934;
  assign n8946 = ~n8936 & ~n8938;
  assign n8947 = n8946 ^ n8934;
  assign n8948 = n8945 & n8947;
  assign n8949 = n8948 ^ n8934;
  assign n8950 = x769 & n8949;
  assign n8951 = ~n8943 & ~n8950;
  assign n8952 = ~n8941 & n8951;
  assign n8991 = n8990 ^ n8952;
  assign n7863 = n7862 ^ n7859;
  assign n7865 = x772 ^ x771;
  assign n7867 = n7866 ^ n7865;
  assign n7864 = x774 ^ x773;
  assign n7868 = n7867 ^ n7864;
  assign n8856 = n7863 & n7868;
  assign n10664 = n8952 ^ n8856;
  assign n10665 = n8991 & ~n10664;
  assign n10666 = n10665 ^ n8990;
  assign n11531 = n10666 ^ n8971;
  assign n10667 = n8937 & ~n8950;
  assign n11532 = n10667 ^ n10666;
  assign n11533 = ~n11531 & n11532;
  assign n11534 = n11533 ^ n8971;
  assign n10668 = n10667 ^ n8971;
  assign n10669 = n10668 ^ n10666;
  assign n8864 = x761 & x762;
  assign n8865 = x759 & x760;
  assign n8866 = ~n8864 & ~n8865;
  assign n8867 = ~x761 & ~x762;
  assign n8868 = ~x759 & ~x760;
  assign n8869 = ~n8867 & ~n8868;
  assign n8870 = ~n8866 & n8869;
  assign n8871 = x758 & n8870;
  assign n8872 = n8864 & n8865;
  assign n8873 = ~n8871 & ~n8872;
  assign n8880 = n8870 ^ x758;
  assign n8881 = n8880 ^ n8870;
  assign n8874 = n8866 & ~n8869;
  assign n8882 = ~n8872 & ~n8874;
  assign n8883 = n8882 ^ n8870;
  assign n8884 = n8881 & n8883;
  assign n8885 = n8884 ^ n8870;
  assign n8886 = x757 & n8885;
  assign n10671 = n8873 & ~n8886;
  assign n8889 = x755 & x756;
  assign n8890 = x753 & x754;
  assign n8891 = n8889 & n8890;
  assign n8892 = ~n8889 & ~n8890;
  assign n8893 = ~x755 & ~x756;
  assign n8894 = ~x753 & ~x754;
  assign n8895 = ~n8893 & ~n8894;
  assign n8896 = ~n8892 & n8895;
  assign n8897 = ~x752 & n8896;
  assign n8898 = ~x751 & n8897;
  assign n8899 = n8898 ^ n8896;
  assign n8900 = ~n8891 & ~n8899;
  assign n8919 = n8892 & ~n8895;
  assign n8908 = x751 & x752;
  assign n8920 = n8890 & n8908;
  assign n8921 = x756 & n8920;
  assign n8922 = n8921 ^ n8908;
  assign n8923 = ~n8919 & n8922;
  assign n10670 = n8900 & ~n8923;
  assign n10672 = n10671 ^ n10670;
  assign n7870 = x756 ^ x755;
  assign n8901 = x755 ^ x752;
  assign n8902 = n7870 & n8901;
  assign n8903 = n8902 ^ x755;
  assign n8904 = n8894 & ~n8903;
  assign n8905 = n8900 & ~n8904;
  assign n8906 = x751 & ~n8897;
  assign n8907 = ~n8905 & ~n8906;
  assign n7872 = x752 ^ x751;
  assign n7871 = x754 ^ x753;
  assign n7873 = n7872 ^ n7871;
  assign n8909 = n8908 ^ n7873;
  assign n8910 = n8909 ^ n8908;
  assign n8911 = ~x752 & ~x756;
  assign n8912 = n8911 ^ n8908;
  assign n8913 = n8912 ^ n8908;
  assign n8914 = n8910 & n8913;
  assign n8915 = n8914 ^ n8908;
  assign n8916 = ~n8890 & n8915;
  assign n8917 = n8916 ^ n8908;
  assign n8918 = ~x755 & n8917;
  assign n8924 = ~n8918 & ~n8923;
  assign n8925 = ~n8907 & n8924;
  assign n8875 = ~x758 & n8874;
  assign n8876 = n8873 & ~n8875;
  assign n8877 = ~x757 & ~n8876;
  assign n7877 = x758 ^ x757;
  assign n8878 = n8867 & n8868;
  assign n8879 = n7877 & n8878;
  assign n8887 = ~n8879 & ~n8886;
  assign n8888 = ~n8877 & n8887;
  assign n8926 = n8925 ^ n8888;
  assign n7874 = n7873 ^ n7870;
  assign n7876 = x760 ^ x759;
  assign n7878 = n7877 ^ n7876;
  assign n7875 = x762 ^ x761;
  assign n7879 = n7878 ^ n7875;
  assign n8860 = n7874 & n7879;
  assign n7880 = n7879 ^ n7874;
  assign n7869 = n7868 ^ n7863;
  assign n8857 = n7874 ^ n7869;
  assign n8858 = n7880 & ~n8857;
  assign n8859 = n8858 ^ n7879;
  assign n8861 = n8860 ^ n8859;
  assign n8862 = ~n8856 & ~n8861;
  assign n8863 = n8862 ^ n8860;
  assign n8927 = n8926 ^ n8863;
  assign n8992 = n8991 ^ n8927;
  assign n10677 = ~n8856 & n8991;
  assign n10678 = ~n8992 & ~n10677;
  assign n10679 = ~n8861 & ~n8926;
  assign n10680 = n10679 ^ n8860;
  assign n10681 = ~n10678 & ~n10680;
  assign n10674 = ~n8860 & n8926;
  assign n10675 = ~n8888 & ~n8925;
  assign n10676 = ~n10674 & ~n10675;
  assign n10682 = n10681 ^ n10676;
  assign n11535 = n10672 & n10682;
  assign n11536 = n10669 & ~n11535;
  assign n11538 = ~n10676 & ~n10681;
  assign n11537 = n10670 & n10671;
  assign n11539 = n11538 ^ n11537;
  assign n11540 = n11536 & ~n11539;
  assign n11541 = ~n10670 & ~n10671;
  assign n11542 = ~n10669 & ~n11541;
  assign n11543 = n11537 ^ n10676;
  assign n11544 = n10682 & ~n11543;
  assign n11545 = n11544 ^ n10676;
  assign n11546 = n11542 & ~n11545;
  assign n11547 = ~n11540 & ~n11546;
  assign n11688 = ~n11534 & n11547;
  assign n11689 = ~n11537 & ~n11538;
  assign n11690 = n11536 & n11689;
  assign n11691 = ~n11688 & ~n11690;
  assign n11693 = n11692 ^ n11691;
  assign n9194 = x813 & x814;
  assign n9193 = x815 & x816;
  assign n9195 = n9194 ^ n9193;
  assign n9196 = ~x813 & ~x814;
  assign n9197 = ~x815 & ~x816;
  assign n9198 = ~n9196 & ~n9197;
  assign n9199 = n9198 ^ n9193;
  assign n9200 = n9199 ^ n9193;
  assign n9201 = n9193 ^ x812;
  assign n9202 = n9201 ^ n9193;
  assign n9203 = n9200 & n9202;
  assign n9204 = n9203 ^ n9193;
  assign n9205 = n9195 & ~n9204;
  assign n9206 = n9205 ^ n9194;
  assign n7829 = x816 ^ x815;
  assign n9207 = x815 ^ x812;
  assign n9208 = n7829 & n9207;
  assign n9209 = n9208 ^ x815;
  assign n9210 = n9196 & ~n9209;
  assign n9211 = ~n9206 & ~n9210;
  assign n9212 = ~x811 & ~n9211;
  assign n9214 = x811 & ~n9196;
  assign n9213 = x811 & x812;
  assign n9215 = n9214 ^ n9213;
  assign n9216 = n9215 ^ n9213;
  assign n9217 = ~x812 & ~x816;
  assign n9218 = n9217 ^ n9213;
  assign n9219 = n9218 ^ n9213;
  assign n9220 = ~n9216 & n9219;
  assign n9221 = n9220 ^ n9213;
  assign n9222 = ~n9194 & n9221;
  assign n9223 = n9222 ^ n9213;
  assign n9224 = ~x815 & n9223;
  assign n7830 = x812 ^ x811;
  assign n9225 = ~n9193 & ~n9194;
  assign n9226 = n9198 & ~n9225;
  assign n9227 = n7830 & n9226;
  assign n9228 = ~n9198 & n9225;
  assign n9229 = n9194 & n9213;
  assign n9230 = x816 & n9229;
  assign n9231 = n9230 ^ n9213;
  assign n9232 = ~n9228 & n9231;
  assign n9233 = ~n9227 & ~n9232;
  assign n9234 = ~n9224 & n9233;
  assign n9235 = ~n9212 & n9234;
  assign n9151 = x819 & x820;
  assign n9150 = x821 & x822;
  assign n9152 = n9151 ^ n9150;
  assign n9153 = ~x819 & ~x820;
  assign n9154 = ~x821 & ~x822;
  assign n9155 = ~n9153 & ~n9154;
  assign n9156 = n9155 ^ n9150;
  assign n9157 = n9156 ^ n9150;
  assign n9158 = n9150 ^ x818;
  assign n9159 = n9158 ^ n9150;
  assign n9160 = n9157 & n9159;
  assign n9161 = n9160 ^ n9150;
  assign n9162 = n9152 & ~n9161;
  assign n9163 = n9162 ^ n9151;
  assign n7824 = x822 ^ x821;
  assign n9164 = x821 ^ x818;
  assign n9165 = n7824 & n9164;
  assign n9166 = n9165 ^ x821;
  assign n9167 = n9153 & ~n9166;
  assign n9168 = ~n9163 & ~n9167;
  assign n9169 = ~x817 & ~n9168;
  assign n9171 = x817 & ~n9153;
  assign n9170 = x817 & x818;
  assign n9172 = n9171 ^ n9170;
  assign n9173 = n9172 ^ n9170;
  assign n9174 = ~x818 & ~x822;
  assign n9175 = n9174 ^ n9170;
  assign n9176 = n9175 ^ n9170;
  assign n9177 = ~n9173 & n9176;
  assign n9178 = n9177 ^ n9170;
  assign n9179 = ~n9151 & n9178;
  assign n9180 = n9179 ^ n9170;
  assign n9181 = ~x821 & n9180;
  assign n7825 = x818 ^ x817;
  assign n9182 = ~n9150 & ~n9151;
  assign n9183 = n9155 & ~n9182;
  assign n9184 = n7825 & n9183;
  assign n9185 = ~n9155 & n9182;
  assign n9186 = n9151 & n9170;
  assign n9187 = x822 & n9186;
  assign n9188 = n9187 ^ n9170;
  assign n9189 = ~n9185 & n9188;
  assign n9190 = ~n9184 & ~n9189;
  assign n9191 = ~n9181 & n9190;
  assign n9192 = ~n9169 & n9191;
  assign n9236 = n9235 ^ n9192;
  assign n7826 = n7825 ^ n7824;
  assign n7823 = x820 ^ x819;
  assign n7827 = n7826 ^ n7823;
  assign n7831 = n7830 ^ n7829;
  assign n7828 = x814 ^ x813;
  assign n7832 = n7831 ^ n7828;
  assign n9239 = n7827 & n7832;
  assign n10760 = n9236 & n9239;
  assign n10761 = n9192 & n9235;
  assign n10762 = ~n10760 & ~n10761;
  assign n10758 = ~n9163 & n9190;
  assign n10757 = ~n9206 & n9233;
  assign n10759 = n10758 ^ n10757;
  assign n10763 = n10762 ^ n10759;
  assign n9242 = x803 & x804;
  assign n9243 = x801 & x802;
  assign n9244 = ~n9242 & ~n9243;
  assign n9245 = ~x803 & ~x804;
  assign n9246 = ~x801 & ~x802;
  assign n9247 = ~n9245 & ~n9246;
  assign n9248 = ~n9244 & n9247;
  assign n9249 = x800 & n9248;
  assign n9250 = n9242 & n9243;
  assign n9251 = ~n9249 & ~n9250;
  assign n9258 = n9248 ^ x800;
  assign n9259 = n9258 ^ n9248;
  assign n9252 = n9244 & ~n9247;
  assign n9260 = ~n9250 & ~n9252;
  assign n9261 = n9260 ^ n9248;
  assign n9262 = n9259 & n9261;
  assign n9263 = n9262 ^ n9248;
  assign n9264 = x799 & n9263;
  assign n10765 = n9251 & ~n9264;
  assign n9268 = x809 & x810;
  assign n9267 = x807 & x808;
  assign n9269 = n9268 ^ n9267;
  assign n9270 = ~x809 & ~x810;
  assign n9271 = ~x807 & ~x808;
  assign n9272 = ~n9270 & ~n9271;
  assign n9273 = n9272 ^ n9267;
  assign n9274 = n9273 ^ n9267;
  assign n9275 = n9267 ^ x806;
  assign n9276 = n9275 ^ n9267;
  assign n9277 = n9274 & n9276;
  assign n9278 = n9277 ^ n9267;
  assign n9279 = n9269 & ~n9278;
  assign n9280 = n9279 ^ n9268;
  assign n7819 = x806 ^ x805;
  assign n9281 = ~n9267 & ~n9268;
  assign n9289 = n9272 & ~n9281;
  assign n9290 = n7819 & n9289;
  assign n9291 = ~n9272 & n9281;
  assign n9292 = x805 & x806;
  assign n9293 = n9267 & n9292;
  assign n9294 = x810 & n9293;
  assign n9295 = n9294 ^ n9292;
  assign n9296 = ~n9291 & n9295;
  assign n9297 = ~n9290 & ~n9296;
  assign n10764 = ~n9280 & n9297;
  assign n10766 = n10765 ^ n10764;
  assign n9282 = n9270 ^ x806;
  assign n9283 = n9271 ^ n9270;
  assign n9284 = ~n9282 & n9283;
  assign n9285 = n9284 ^ n9270;
  assign n9286 = n9281 & n9285;
  assign n9287 = ~n9280 & ~n9286;
  assign n9288 = ~x805 & ~n9287;
  assign n7818 = x808 ^ x807;
  assign n9298 = n9292 ^ x808;
  assign n9299 = n9298 ^ n9292;
  assign n9300 = ~x806 & ~x810;
  assign n9301 = n9300 ^ n9292;
  assign n9302 = ~n9299 & n9301;
  assign n9303 = n9302 ^ n9292;
  assign n9304 = ~n7818 & n9303;
  assign n9305 = ~x809 & n9304;
  assign n9306 = n9297 & ~n9305;
  assign n9307 = ~n9288 & n9306;
  assign n9253 = ~x800 & n9252;
  assign n9254 = n9251 & ~n9253;
  assign n9255 = ~x799 & ~n9254;
  assign n7814 = x800 ^ x799;
  assign n9256 = n9245 & n9246;
  assign n9257 = n7814 & n9256;
  assign n9265 = ~n9257 & ~n9264;
  assign n9266 = ~n9255 & n9265;
  assign n9308 = n9307 ^ n9266;
  assign n7820 = n7819 ^ n7818;
  assign n7817 = x810 ^ x809;
  assign n7821 = n7820 ^ n7817;
  assign n7813 = x802 ^ x801;
  assign n7815 = n7814 ^ n7813;
  assign n7812 = x804 ^ x803;
  assign n7816 = n7815 ^ n7812;
  assign n7822 = n7821 ^ n7816;
  assign n7833 = n7832 ^ n7827;
  assign n9237 = n7822 & n7833;
  assign n9238 = n7816 & n7821;
  assign n9240 = n9239 ^ n9238;
  assign n9241 = ~n9237 & ~n9240;
  assign n9309 = n9308 ^ n9241;
  assign n9310 = n9309 ^ n9236;
  assign n10769 = ~n9237 & ~n9238;
  assign n10771 = n9266 & n9307;
  assign n10776 = ~n10769 & n10771;
  assign n10777 = n9310 & n10776;
  assign n10768 = ~n9266 & ~n9307;
  assign n10770 = n10768 & n10769;
  assign n10772 = n9239 ^ n9236;
  assign n10773 = ~n9310 & ~n10772;
  assign n10774 = ~n10771 & n10773;
  assign n10775 = ~n10770 & ~n10774;
  assign n11506 = n10777 ^ n10775;
  assign n11507 = n11506 ^ n10777;
  assign n11508 = n10777 ^ n10764;
  assign n11509 = n11508 ^ n10777;
  assign n11510 = n11507 & n11509;
  assign n11511 = n11510 ^ n10777;
  assign n11512 = ~n10766 & ~n11511;
  assign n11513 = n11512 ^ n10777;
  assign n11514 = ~n10763 & ~n11513;
  assign n11515 = n10765 ^ n10763;
  assign n11516 = n10775 & ~n11515;
  assign n11517 = n11516 ^ n10765;
  assign n11518 = ~n10764 & ~n11517;
  assign n11519 = ~n11514 & ~n11518;
  assign n11520 = n10763 & n10775;
  assign n11521 = n10765 & ~n10777;
  assign n11522 = n11520 & ~n11521;
  assign n11523 = n11519 & ~n11522;
  assign n11503 = n10762 ^ n10758;
  assign n11504 = ~n10759 & n11503;
  assign n11505 = n11504 ^ n10762;
  assign n11524 = n11523 ^ n11505;
  assign n9041 = x839 & x840;
  assign n9040 = x837 & x838;
  assign n9042 = n9041 ^ n9040;
  assign n9043 = ~x839 & ~x840;
  assign n9044 = ~x837 & ~x838;
  assign n9045 = ~n9043 & ~n9044;
  assign n9046 = n9045 ^ n9040;
  assign n9047 = n9046 ^ n9040;
  assign n9048 = n9040 ^ x836;
  assign n9049 = n9048 ^ n9040;
  assign n9050 = n9047 & n9049;
  assign n9051 = n9050 ^ n9040;
  assign n9052 = n9042 & ~n9051;
  assign n9053 = n9052 ^ n9041;
  assign n9071 = ~n9040 & ~n9041;
  assign n9072 = ~n9045 & n9071;
  assign n9060 = x835 & x836;
  assign n9073 = n9040 & n9060;
  assign n9074 = x840 & n9073;
  assign n9075 = n9074 ^ n9060;
  assign n9076 = ~n9072 & n9075;
  assign n7841 = x836 ^ x835;
  assign n9077 = n9045 & ~n9071;
  assign n9078 = n7841 & n9077;
  assign n9079 = ~n9076 & ~n9078;
  assign n10751 = ~n9053 & n9079;
  assign n8999 = x845 & x846;
  assign n8998 = x843 & x844;
  assign n9000 = n8999 ^ n8998;
  assign n9001 = ~x845 & ~x846;
  assign n9002 = ~x843 & ~x844;
  assign n9003 = ~n9001 & ~n9002;
  assign n9004 = n9003 ^ n8998;
  assign n9005 = n9004 ^ n8998;
  assign n9006 = n8998 ^ x842;
  assign n9007 = n9006 ^ n8998;
  assign n9008 = n9005 & n9007;
  assign n9009 = n9008 ^ n8998;
  assign n9010 = n9000 & ~n9009;
  assign n9011 = n9010 ^ n8999;
  assign n9029 = ~n8998 & ~n8999;
  assign n9030 = ~n9003 & n9029;
  assign n9018 = x841 & x842;
  assign n9031 = n8998 & n9018;
  assign n9032 = x846 & n9031;
  assign n9033 = n9032 ^ n9018;
  assign n9034 = ~n9030 & n9033;
  assign n7836 = x842 ^ x841;
  assign n9035 = n9003 & ~n9029;
  assign n9036 = n7836 & n9035;
  assign n9037 = ~n9034 & ~n9036;
  assign n10750 = ~n9011 & n9037;
  assign n10752 = n10751 ^ n10750;
  assign n7840 = x840 ^ x839;
  assign n9054 = x839 ^ x836;
  assign n9055 = n7840 & n9054;
  assign n9056 = n9055 ^ x839;
  assign n9057 = n9044 & ~n9056;
  assign n9058 = ~n9053 & ~n9057;
  assign n9059 = ~x835 & ~n9058;
  assign n7842 = x838 ^ x837;
  assign n7843 = n7842 ^ n7841;
  assign n9061 = n9060 ^ n7843;
  assign n9062 = n9061 ^ n9060;
  assign n9063 = ~x836 & ~x840;
  assign n9064 = n9063 ^ n9060;
  assign n9065 = n9064 ^ n9060;
  assign n9066 = n9062 & n9065;
  assign n9067 = n9066 ^ n9060;
  assign n9068 = ~n9040 & n9067;
  assign n9069 = n9068 ^ n9060;
  assign n9070 = ~x839 & n9069;
  assign n9080 = ~n9070 & n9079;
  assign n9081 = ~n9059 & n9080;
  assign n7835 = x846 ^ x845;
  assign n9012 = x845 ^ x842;
  assign n9013 = n7835 & n9012;
  assign n9014 = n9013 ^ x845;
  assign n9015 = n9002 & ~n9014;
  assign n9016 = ~n9011 & ~n9015;
  assign n9017 = ~x841 & ~n9016;
  assign n7837 = x844 ^ x843;
  assign n7838 = n7837 ^ n7836;
  assign n9019 = n9018 ^ n7838;
  assign n9020 = n9019 ^ n9018;
  assign n9021 = ~x842 & ~x846;
  assign n9022 = n9021 ^ n9018;
  assign n9023 = n9022 ^ n9018;
  assign n9024 = n9020 & n9023;
  assign n9025 = n9024 ^ n9018;
  assign n9026 = ~n8998 & n9025;
  assign n9027 = n9026 ^ n9018;
  assign n9028 = ~x845 & n9027;
  assign n9038 = ~n9028 & n9037;
  assign n9039 = ~n9017 & n9038;
  assign n9082 = n9081 ^ n9039;
  assign n7839 = n7838 ^ n7835;
  assign n7844 = n7843 ^ n7840;
  assign n8996 = n7839 & n7844;
  assign n10747 = n9039 ^ n8996;
  assign n10748 = n9082 & ~n10747;
  assign n10749 = n10748 ^ n9081;
  assign n10753 = n10752 ^ n10749;
  assign n7853 = x824 ^ x823;
  assign n7852 = x826 ^ x825;
  assign n9110 = x827 & x828;
  assign n9111 = n9110 ^ x826;
  assign n9112 = n7852 & ~n9111;
  assign n9113 = n9112 ^ x825;
  assign n9114 = n7853 & n9113;
  assign n9115 = ~x825 & ~x826;
  assign n9116 = ~n9110 & n9115;
  assign n9117 = x825 & x826;
  assign n9118 = x823 & x824;
  assign n9119 = ~n9117 & n9118;
  assign n9120 = ~n9116 & n9119;
  assign n9121 = ~n9114 & ~n9120;
  assign n9122 = ~x827 & ~x828;
  assign n9123 = ~n9121 & ~n9122;
  assign n9124 = n9117 & n9118;
  assign n9125 = ~x828 & n9124;
  assign n9126 = ~n9123 & ~n9125;
  assign n9127 = n9110 & n9117;
  assign n9128 = x824 & ~n9122;
  assign n9129 = ~n9127 & ~n9128;
  assign n9130 = n9113 & ~n9129;
  assign n9131 = n9116 & ~n9128;
  assign n9132 = ~n9130 & ~n9131;
  assign n9133 = ~x823 & ~n9132;
  assign n9134 = ~x824 & ~x828;
  assign n9135 = n9134 ^ n9118;
  assign n9136 = n9135 ^ n9118;
  assign n7854 = n7853 ^ n7852;
  assign n9137 = n9118 ^ n7854;
  assign n9138 = n9137 ^ n9118;
  assign n9139 = n9136 & n9138;
  assign n9140 = n9139 ^ n9118;
  assign n9141 = ~n9117 & n9140;
  assign n9142 = n9141 ^ n9118;
  assign n9143 = ~x827 & n9142;
  assign n9144 = ~n9133 & ~n9143;
  assign n9145 = n9126 & n9144;
  assign n7848 = x830 ^ x829;
  assign n7847 = x832 ^ x831;
  assign n7849 = n7848 ^ n7847;
  assign n7846 = x834 ^ x833;
  assign n7850 = n7849 ^ n7846;
  assign n7851 = x828 ^ x827;
  assign n7855 = n7854 ^ n7851;
  assign n9109 = n7850 & n7855;
  assign n9146 = n9145 ^ n9109;
  assign n9084 = x831 & x832;
  assign n9085 = x833 & x834;
  assign n9086 = n9084 & n9085;
  assign n9087 = ~x833 & ~x834;
  assign n9088 = ~n9084 & n9087;
  assign n9089 = ~n9086 & ~n9088;
  assign n9090 = ~x831 & ~x832;
  assign n9091 = ~n9085 & n9090;
  assign n9092 = x829 & x830;
  assign n9093 = ~n9091 & n9092;
  assign n9094 = n9089 & n9093;
  assign n9095 = n7848 & ~n9087;
  assign n9096 = n9085 ^ x832;
  assign n9097 = n7847 & ~n9096;
  assign n9098 = n9097 ^ x831;
  assign n9099 = n9095 & n9098;
  assign n9100 = ~n9094 & ~n9099;
  assign n9101 = x830 & ~n9087;
  assign n9102 = n9091 & ~n9101;
  assign n9103 = ~n9086 & ~n9102;
  assign n9104 = ~x829 & ~n9103;
  assign n9105 = n9100 & ~n9104;
  assign n9106 = ~x830 & n9088;
  assign n9107 = n7849 & n9106;
  assign n9108 = n9105 & ~n9107;
  assign n9147 = n9146 ^ n9108;
  assign n7845 = n7844 ^ n7839;
  assign n7856 = n7855 ^ n7850;
  assign n8995 = n7845 & n7856;
  assign n10738 = n9147 ^ n8995;
  assign n10739 = n9082 ^ n8996;
  assign n10740 = n10739 ^ n9082;
  assign n10741 = n9082 ^ n8995;
  assign n10742 = n10741 ^ n9082;
  assign n10743 = ~n10740 & ~n10742;
  assign n10744 = n10743 ^ n9082;
  assign n10745 = n10738 & n10744;
  assign n10746 = n10745 ^ n9147;
  assign n10754 = n10753 ^ n10746;
  assign n10735 = n9126 & ~n9130;
  assign n10734 = ~n9086 & n9100;
  assign n10736 = n10735 ^ n10734;
  assign n10731 = n9109 ^ n9108;
  assign n10732 = n9146 & ~n10731;
  assign n10733 = n10732 ^ n9145;
  assign n10737 = n10736 ^ n10733;
  assign n10755 = n10754 ^ n10737;
  assign n8997 = ~n8995 & ~n8996;
  assign n9083 = n9082 ^ n8997;
  assign n9148 = n9147 ^ n9083;
  assign n7834 = n7833 ^ n7822;
  assign n7857 = n7856 ^ n7845;
  assign n8994 = n7834 & n7857;
  assign n9149 = n9148 ^ n8994;
  assign n10728 = n9310 ^ n9148;
  assign n10729 = n9149 & n10728;
  assign n10730 = n10729 ^ n9310;
  assign n10756 = n10755 ^ n10730;
  assign n10778 = n10775 & ~n10777;
  assign n10767 = n10766 ^ n10763;
  assign n10779 = n10778 ^ n10767;
  assign n11500 = n10779 ^ n10755;
  assign n11501 = n10756 & ~n11500;
  assign n11502 = n11501 ^ n10779;
  assign n11525 = n11524 ^ n11502;
  assign n11486 = ~n10746 & ~n10753;
  assign n11487 = n10733 & ~n11486;
  assign n11488 = ~n10734 & ~n10735;
  assign n11489 = ~n11487 & ~n11488;
  assign n11490 = n10734 & n10735;
  assign n11491 = ~n10755 & ~n11490;
  assign n11492 = n11489 & ~n11491;
  assign n11493 = n10746 & n10753;
  assign n11494 = ~n11487 & ~n11493;
  assign n11495 = n11491 & ~n11494;
  assign n11496 = ~n11492 & ~n11495;
  assign n11483 = n10751 ^ n10749;
  assign n11484 = ~n10752 & ~n11483;
  assign n11485 = n11484 ^ n10749;
  assign n11497 = n11496 ^ n11485;
  assign n11498 = n11489 & n11493;
  assign n11499 = ~n11497 & ~n11498;
  assign n11526 = n11525 ^ n11499;
  assign n8782 = n8781 ^ n8690;
  assign n8854 = n8853 ^ n8782;
  assign n7881 = n7880 ^ n7869;
  assign n8681 = n7881 & n7904;
  assign n8682 = n7897 ^ n7892;
  assign n8683 = n7903 & ~n8682;
  assign n8684 = n8683 ^ n7902;
  assign n8685 = ~n8681 & ~n8684;
  assign n8687 = n7892 & n8686;
  assign n8688 = n7881 & n8687;
  assign n8689 = ~n8685 & ~n8688;
  assign n8855 = n8854 ^ n8689;
  assign n10684 = n8855 & n8992;
  assign n10685 = n8684 & ~n8688;
  assign n10686 = n10685 ^ n8685;
  assign n10687 = n8854 & n10686;
  assign n10688 = n10687 ^ n8685;
  assign n10689 = ~n10684 & ~n10688;
  assign n10725 = n10724 ^ n10689;
  assign n10673 = n10672 ^ n10669;
  assign n10683 = n10682 ^ n10673;
  assign n10726 = n10725 ^ n10683;
  assign n7858 = n7857 ^ n7834;
  assign n7905 = n7904 ^ n7881;
  assign n9314 = n7858 & n7905;
  assign n9311 = n9310 ^ n9149;
  assign n10660 = n9314 ^ n9311;
  assign n8993 = n8992 ^ n8855;
  assign n10661 = n9314 ^ n8993;
  assign n10662 = n10660 & n10661;
  assign n10663 = n10662 ^ n9311;
  assign n10727 = n10726 ^ n10663;
  assign n10780 = n10779 ^ n10756;
  assign n11480 = n10780 ^ n10663;
  assign n11481 = n10727 & ~n11480;
  assign n11482 = n11481 ^ n10726;
  assign n11527 = n11526 ^ n11482;
  assign n11562 = n11555 & n11561;
  assign n11566 = ~n10707 & n11560;
  assign n11567 = ~n11565 & ~n11566;
  assign n11568 = ~n11562 & n11567;
  assign n11569 = n11568 ^ n11551;
  assign n11548 = n11547 ^ n11534;
  assign n11570 = n11569 ^ n11548;
  assign n11528 = n10689 ^ n10683;
  assign n11529 = n10725 & ~n11528;
  assign n11530 = n11529 ^ n10724;
  assign n11571 = n11570 ^ n11530;
  assign n11685 = n11571 ^ n11526;
  assign n11686 = ~n11527 & ~n11685;
  assign n11687 = n11686 ^ n11571;
  assign n11694 = n11693 ^ n11687;
  assign n11677 = ~n10764 & ~n10765;
  assign n11678 = n11524 & ~n11677;
  assign n11679 = n11517 & ~n11521;
  assign n11680 = n11505 & ~n11679;
  assign n11681 = ~n11678 & ~n11680;
  assign n11675 = ~n11485 & ~n11495;
  assign n11676 = ~n11492 & ~n11675;
  assign n11682 = n11681 ^ n11676;
  assign n11672 = n11502 ^ n11499;
  assign n11673 = ~n11525 & ~n11672;
  assign n11674 = n11673 ^ n11524;
  assign n11683 = n11682 ^ n11674;
  assign n11669 = n11548 ^ n11530;
  assign n11670 = ~n11570 & n11669;
  assign n11671 = n11670 ^ n11569;
  assign n11684 = n11683 ^ n11671;
  assign n11695 = n11694 ^ n11684;
  assign n11718 = n11671 & n11683;
  assign n11719 = n11691 & ~n11692;
  assign n11720 = n11718 & ~n11719;
  assign n11721 = ~n11687 & n11720;
  assign n11726 = ~n11691 & n11692;
  assign n11786 = ~n11721 & ~n11726;
  assign n11787 = ~n11671 & n11786;
  assign n11788 = n11695 & n11787;
  assign n11722 = ~n11683 & n11719;
  assign n11789 = n11687 & n11722;
  assign n11790 = ~n11676 & ~n11681;
  assign n11791 = ~n11674 & n11790;
  assign n11792 = ~n11789 & ~n11791;
  assign n11793 = ~n11788 & n11792;
  assign n11715 = n11681 ^ n11674;
  assign n11716 = ~n11682 & n11715;
  assign n11717 = n11716 ^ n11674;
  assign n11725 = ~n11671 & n11687;
  assign n11794 = ~n11725 & ~n11786;
  assign n11795 = ~n11717 & ~n11794;
  assign n11796 = n11793 & ~n11795;
  assign n11704 = n11661 ^ n11659;
  assign n11705 = ~n11665 & n11704;
  assign n11706 = n11705 ^ n11664;
  assign n11723 = ~n11671 & n11722;
  assign n11724 = ~n11721 & ~n11723;
  assign n11727 = n11683 & n11726;
  assign n11728 = ~n11725 & n11727;
  assign n11729 = n11724 & ~n11728;
  assign n11730 = n11693 ^ n11671;
  assign n11731 = n11730 ^ n11684;
  assign n11732 = n11692 ^ n11683;
  assign n11733 = n11732 ^ n11671;
  assign n11734 = n11733 ^ n11671;
  assign n11735 = n11693 & n11734;
  assign n11736 = n11735 ^ n11693;
  assign n11737 = n11733 & n11736;
  assign n11738 = n11737 ^ n11671;
  assign n11739 = ~n11731 & n11738;
  assign n11740 = n11739 ^ n11735;
  assign n11741 = n11740 ^ n11671;
  assign n11742 = n11741 ^ n11684;
  assign n11743 = n11687 & ~n11742;
  assign n11744 = n11729 & ~n11743;
  assign n11745 = n11744 ^ n11717;
  assign n11668 = n11667 ^ n11647;
  assign n11696 = n11695 ^ n11668;
  assign n11478 = n11477 ^ n11434;
  assign n10892 = n10891 ^ n10791;
  assign n10781 = n10780 ^ n10727;
  assign n10893 = n10892 ^ n10781;
  assign n7906 = n7905 ^ n7858;
  assign n8001 = n8000 ^ n7953;
  assign n8002 = n7906 & n8001;
  assign n9312 = n9311 ^ n8993;
  assign n8005 = ~n8003 & ~n8004;
  assign n8315 = n8314 ^ n8005;
  assign n8680 = n8679 ^ n8315;
  assign n9313 = n9312 ^ n8680;
  assign n9315 = n9314 ^ n9313;
  assign n10894 = ~n8002 & ~n9315;
  assign n10895 = n8002 & ~n9312;
  assign n10896 = ~n8680 & ~n10895;
  assign n10897 = ~n10894 & ~n10896;
  assign n11388 = n10897 ^ n10781;
  assign n11389 = ~n10893 & ~n11388;
  assign n11390 = n11389 ^ n10892;
  assign n11479 = n11478 ^ n11390;
  assign n11572 = n11571 ^ n11527;
  assign n11642 = n11572 ^ n11478;
  assign n11643 = ~n11479 & n11642;
  assign n11644 = n11643 ^ n11572;
  assign n11712 = n11668 ^ n11644;
  assign n11713 = ~n11696 & ~n11712;
  assign n11714 = n11713 ^ n11695;
  assign n11746 = n11745 ^ n11714;
  assign n11847 = n11706 & n11746;
  assign n11848 = n11796 & n11847;
  assign n11849 = n11806 & ~n11848;
  assign n11803 = n11706 & n11745;
  assign n11850 = n11714 & n11745;
  assign n11851 = ~n11796 & ~n11850;
  assign n11852 = ~n11803 & n11851;
  assign n11853 = ~n11849 & ~n11852;
  assign n11802 = ~n11703 & ~n11709;
  assign n11854 = ~n11706 & ~n11746;
  assign n11855 = ~n11714 & ~n11796;
  assign n11856 = ~n11854 & ~n11855;
  assign n11857 = ~n11802 & ~n11856;
  assign n11858 = n11853 & ~n11857;
  assign n10088 = x615 & x616;
  assign n10087 = x617 & x618;
  assign n10089 = n10088 ^ n10087;
  assign n10090 = ~x615 & ~x616;
  assign n10091 = ~x617 & ~x618;
  assign n10092 = ~n10090 & ~n10091;
  assign n10093 = n10092 ^ n10087;
  assign n10094 = n10093 ^ n10087;
  assign n10095 = n10087 ^ x614;
  assign n10096 = n10095 ^ n10087;
  assign n10097 = n10094 & n10096;
  assign n10098 = n10097 ^ n10087;
  assign n10099 = n10089 & ~n10098;
  assign n10100 = n10099 ^ n10088;
  assign n10101 = ~n10087 & ~n10088;
  assign n10102 = n10090 ^ x614;
  assign n10103 = n10091 ^ n10090;
  assign n10104 = ~n10102 & n10103;
  assign n10105 = n10104 ^ n10090;
  assign n10106 = n10101 & n10105;
  assign n10107 = ~n10100 & ~n10106;
  assign n10108 = ~x613 & ~n10107;
  assign n9453 = x614 ^ x613;
  assign n10109 = n10092 & ~n10101;
  assign n10110 = n9453 & n10109;
  assign n10111 = ~n10092 & n10101;
  assign n10112 = x613 & x614;
  assign n10113 = n10088 & n10112;
  assign n10114 = x618 & n10113;
  assign n10115 = n10114 ^ n10112;
  assign n10116 = ~n10111 & n10115;
  assign n10117 = ~n10110 & ~n10116;
  assign n9452 = x616 ^ x615;
  assign n10118 = n10112 ^ x616;
  assign n10119 = n10118 ^ n10112;
  assign n10120 = ~x614 & ~x618;
  assign n10121 = n10120 ^ n10112;
  assign n10122 = ~n10119 & n10121;
  assign n10123 = n10122 ^ n10112;
  assign n10124 = ~n9452 & n10123;
  assign n10125 = ~x617 & n10124;
  assign n10126 = n10117 & ~n10125;
  assign n10127 = ~n10108 & n10126;
  assign n10051 = x609 & x610;
  assign n10050 = x611 & x612;
  assign n10052 = n10051 ^ n10050;
  assign n10053 = ~x609 & ~x610;
  assign n10054 = ~x611 & ~x612;
  assign n10055 = ~n10053 & ~n10054;
  assign n10056 = n10055 ^ n10050;
  assign n10057 = n10056 ^ n10050;
  assign n10058 = n10050 ^ x608;
  assign n10059 = n10058 ^ n10050;
  assign n10060 = n10057 & n10059;
  assign n10061 = n10060 ^ n10050;
  assign n10062 = n10052 & ~n10061;
  assign n10063 = n10062 ^ n10051;
  assign n9446 = x612 ^ x611;
  assign n10064 = x611 ^ x608;
  assign n10065 = n9446 & n10064;
  assign n10066 = n10065 ^ x611;
  assign n10067 = n10053 & ~n10066;
  assign n10068 = ~n10063 & ~n10067;
  assign n10069 = ~x607 & ~n10068;
  assign n9448 = x608 ^ x607;
  assign n10070 = ~n10050 & ~n10051;
  assign n10071 = n10055 & ~n10070;
  assign n10072 = n9448 & n10071;
  assign n10073 = ~n10055 & n10070;
  assign n10074 = x612 & n10051;
  assign n10075 = x607 & x608;
  assign n10076 = ~n10074 & n10075;
  assign n10077 = ~n10073 & n10076;
  assign n10078 = ~n10072 & ~n10077;
  assign n9447 = x610 ^ x609;
  assign n9449 = n9448 ^ n9447;
  assign n10079 = ~x608 & ~n10051;
  assign n10080 = n10054 & n10079;
  assign n10081 = n9449 & n10080;
  assign n10082 = ~x611 & n10051;
  assign n10083 = n10075 & n10082;
  assign n10084 = ~n10081 & ~n10083;
  assign n10085 = n10078 & n10084;
  assign n10086 = ~n10069 & n10085;
  assign n10128 = n10127 ^ n10086;
  assign n9435 = x628 ^ x627;
  assign n10025 = x629 & x630;
  assign n10026 = n10025 ^ x628;
  assign n10027 = ~n9435 & ~n10026;
  assign n10028 = ~x625 & n10027;
  assign n10029 = x627 & x628;
  assign n10030 = ~x629 & ~x630;
  assign n10031 = ~n10029 & n10030;
  assign n10032 = ~x626 & n10031;
  assign n10033 = ~n10028 & ~n10032;
  assign n10034 = ~x627 & ~x628;
  assign n10035 = x625 & ~n10034;
  assign n10036 = x626 & ~n10030;
  assign n10037 = ~n10035 & ~n10036;
  assign n10038 = ~n10033 & n10037;
  assign n9437 = x626 ^ x625;
  assign n10039 = n10025 & ~n10034;
  assign n10040 = n10029 & ~n10030;
  assign n10041 = ~n10039 & ~n10040;
  assign n10042 = n9437 & ~n10041;
  assign n10043 = x625 & x626;
  assign n10044 = ~n10031 & n10043;
  assign n10045 = ~n10027 & n10044;
  assign n10046 = ~n10042 & ~n10045;
  assign n10047 = ~n10038 & n10046;
  assign n9440 = x622 ^ x621;
  assign n10002 = x623 & x624;
  assign n10003 = n10002 ^ x622;
  assign n10004 = ~n9440 & ~n10003;
  assign n10005 = ~x619 & n10004;
  assign n10006 = x621 & x622;
  assign n10007 = ~x623 & ~x624;
  assign n10008 = ~n10006 & n10007;
  assign n10009 = ~x620 & n10008;
  assign n10010 = ~n10005 & ~n10009;
  assign n10011 = ~x621 & ~x622;
  assign n10012 = x619 & ~n10011;
  assign n10013 = x620 & ~n10007;
  assign n10014 = ~n10012 & ~n10013;
  assign n10015 = ~n10010 & n10014;
  assign n9442 = x620 ^ x619;
  assign n10016 = n10002 & ~n10011;
  assign n10017 = n10006 & ~n10007;
  assign n10018 = ~n10016 & ~n10017;
  assign n10019 = n9442 & ~n10018;
  assign n10020 = x619 & x620;
  assign n10021 = ~n10008 & n10020;
  assign n10022 = ~n10004 & n10021;
  assign n10023 = ~n10019 & ~n10022;
  assign n10024 = ~n10015 & n10023;
  assign n10048 = n10047 ^ n10024;
  assign n9441 = x624 ^ x623;
  assign n9443 = n9442 ^ n9441;
  assign n9444 = n9443 ^ n9440;
  assign n9436 = x630 ^ x629;
  assign n9438 = n9437 ^ n9436;
  assign n9439 = n9438 ^ n9435;
  assign n9445 = n9444 ^ n9439;
  assign n9454 = n9453 ^ n9452;
  assign n9451 = x618 ^ x617;
  assign n9455 = n9454 ^ n9451;
  assign n9450 = n9449 ^ n9446;
  assign n9456 = n9455 ^ n9450;
  assign n9997 = n9445 & n9456;
  assign n9999 = n9450 & n9455;
  assign n9998 = n9439 & n9444;
  assign n10000 = n9999 ^ n9998;
  assign n10001 = ~n9997 & ~n10000;
  assign n10049 = n10048 ^ n10001;
  assign n10129 = n10128 ^ n10049;
  assign n11155 = ~n9998 & n10048;
  assign n11156 = ~n10129 & ~n11155;
  assign n11157 = n10128 ^ n9999;
  assign n11158 = ~n9997 & ~n11157;
  assign n11159 = ~n11156 & ~n11158;
  assign n11154 = ~n10100 & n10117;
  assign n11160 = n11159 ^ n11154;
  assign n11151 = ~n10063 & n10078;
  assign n11148 = n10086 ^ n9999;
  assign n11149 = n10128 & ~n11148;
  assign n11150 = n11149 ^ n10127;
  assign n11152 = n11151 ^ n11150;
  assign n11144 = n10025 & n10029;
  assign n11145 = n10046 & ~n11144;
  assign n11142 = n10002 & n10006;
  assign n11143 = n10023 & ~n11142;
  assign n11146 = n11145 ^ n11143;
  assign n11139 = n10024 ^ n9998;
  assign n11140 = n10048 & ~n11139;
  assign n11141 = n11140 ^ n10047;
  assign n11147 = n11146 ^ n11141;
  assign n11153 = n11152 ^ n11147;
  assign n11161 = n11160 ^ n11153;
  assign n11204 = n11154 & ~n11159;
  assign n11205 = ~n11150 & n11151;
  assign n11206 = ~n11204 & ~n11205;
  assign n11207 = n11147 & n11206;
  assign n11208 = ~n11161 & n11207;
  assign n11209 = ~n11147 & n11161;
  assign n11210 = n11209 ^ n11204;
  assign n11211 = n11205 ^ n11204;
  assign n11212 = n11210 & ~n11211;
  assign n11213 = n11212 ^ n11209;
  assign n11214 = ~n11208 & ~n11213;
  assign n11201 = n11145 ^ n11141;
  assign n11202 = ~n11146 & ~n11201;
  assign n11203 = n11202 ^ n11141;
  assign n11215 = n11214 ^ n11203;
  assign n9414 = x638 ^ x637;
  assign n9413 = x640 ^ x639;
  assign n9959 = x641 & x642;
  assign n9960 = n9959 ^ x640;
  assign n9961 = n9413 & ~n9960;
  assign n9962 = n9961 ^ x639;
  assign n9963 = n9414 & n9962;
  assign n9964 = ~x639 & ~x640;
  assign n9965 = ~n9959 & n9964;
  assign n9966 = x639 & x640;
  assign n9967 = x637 & x638;
  assign n9968 = ~n9966 & n9967;
  assign n9969 = ~n9965 & n9968;
  assign n9970 = ~n9963 & ~n9969;
  assign n9971 = ~x641 & ~x642;
  assign n9972 = ~n9970 & ~n9971;
  assign n9973 = n9966 & n9967;
  assign n9974 = ~x642 & n9973;
  assign n9975 = ~n9972 & ~n9974;
  assign n9976 = x638 & ~n9971;
  assign n9977 = n9959 & n9966;
  assign n9978 = ~n9976 & ~n9977;
  assign n9979 = n9962 & ~n9978;
  assign n9980 = n9965 & ~n9976;
  assign n9981 = ~n9979 & ~n9980;
  assign n9982 = ~x637 & ~n9981;
  assign n9983 = n9975 & ~n9982;
  assign n9984 = ~x638 & ~x642;
  assign n9985 = n9984 ^ n9967;
  assign n9986 = n9985 ^ n9967;
  assign n9415 = n9414 ^ n9413;
  assign n9987 = n9967 ^ n9415;
  assign n9988 = n9987 ^ n9967;
  assign n9989 = n9986 & n9988;
  assign n9990 = n9989 ^ n9967;
  assign n9991 = ~n9966 & n9990;
  assign n9992 = n9991 ^ n9967;
  assign n9993 = ~x641 & n9992;
  assign n9994 = n9983 & ~n9993;
  assign n9915 = x633 & x634;
  assign n9914 = x635 & x636;
  assign n9916 = n9915 ^ n9914;
  assign n9917 = ~x633 & ~x634;
  assign n9918 = ~x635 & ~x636;
  assign n9919 = ~n9917 & ~n9918;
  assign n9920 = n9919 ^ n9914;
  assign n9921 = n9920 ^ n9914;
  assign n9922 = n9914 ^ x632;
  assign n9923 = n9922 ^ n9914;
  assign n9924 = n9921 & n9923;
  assign n9925 = n9924 ^ n9914;
  assign n9926 = n9916 & ~n9925;
  assign n9927 = n9926 ^ n9915;
  assign n9928 = n9918 ^ n9917;
  assign n9929 = ~n9914 & ~n9915;
  assign n9930 = n9929 ^ n9918;
  assign n9931 = n9930 ^ n9918;
  assign n9932 = n9918 ^ x632;
  assign n9933 = n9932 ^ n9918;
  assign n9934 = n9931 & ~n9933;
  assign n9935 = n9934 ^ n9918;
  assign n9936 = n9928 & ~n9935;
  assign n9937 = n9936 ^ n9917;
  assign n9938 = ~n9927 & ~n9937;
  assign n9939 = ~x631 & ~n9938;
  assign n9419 = x632 ^ x631;
  assign n9940 = n9919 & ~n9929;
  assign n9941 = n9419 & n9940;
  assign n9942 = ~n9919 & n9929;
  assign n9943 = x631 & x632;
  assign n9944 = n9915 & n9943;
  assign n9945 = x636 & n9944;
  assign n9946 = n9945 ^ n9943;
  assign n9947 = ~n9942 & n9946;
  assign n9948 = ~n9941 & ~n9947;
  assign n9418 = x634 ^ x633;
  assign n9949 = n9943 ^ x634;
  assign n9950 = n9949 ^ n9943;
  assign n9951 = ~x632 & ~x636;
  assign n9952 = n9951 ^ n9943;
  assign n9953 = ~n9950 & n9952;
  assign n9954 = n9953 ^ n9943;
  assign n9955 = ~n9418 & n9954;
  assign n9956 = ~x635 & n9955;
  assign n9957 = n9948 & ~n9956;
  assign n9958 = ~n9939 & n9957;
  assign n9995 = n9994 ^ n9958;
  assign n9876 = x651 & x652;
  assign n9875 = x653 & x654;
  assign n9877 = n9876 ^ n9875;
  assign n9878 = ~x653 & ~x654;
  assign n9879 = ~x651 & ~x652;
  assign n9880 = ~n9878 & ~n9879;
  assign n9881 = n9880 ^ n9875;
  assign n9882 = n9881 ^ n9875;
  assign n9883 = n9875 ^ x650;
  assign n9884 = n9883 ^ n9875;
  assign n9885 = n9882 & n9884;
  assign n9886 = n9885 ^ n9875;
  assign n9887 = n9877 & ~n9886;
  assign n9888 = n9887 ^ n9876;
  assign n9423 = x654 ^ x653;
  assign n9889 = x653 ^ x650;
  assign n9890 = n9423 & n9889;
  assign n9891 = n9890 ^ x653;
  assign n9892 = n9879 & ~n9891;
  assign n9893 = ~n9888 & ~n9892;
  assign n9894 = ~x649 & ~n9893;
  assign n9425 = x650 ^ x649;
  assign n9895 = ~n9875 & ~n9876;
  assign n9896 = n9880 & ~n9895;
  assign n9897 = n9425 & n9896;
  assign n9898 = ~n9880 & n9895;
  assign n9899 = x654 & n9876;
  assign n9900 = x649 & x650;
  assign n9901 = ~n9899 & n9900;
  assign n9902 = ~n9898 & n9901;
  assign n9903 = ~n9897 & ~n9902;
  assign n9424 = x652 ^ x651;
  assign n9426 = n9425 ^ n9424;
  assign n9904 = ~x650 & ~n9876;
  assign n9905 = n9878 & n9904;
  assign n9906 = n9426 & n9905;
  assign n9907 = ~x653 & n9876;
  assign n9908 = n9900 & n9907;
  assign n9909 = ~n9906 & ~n9908;
  assign n9910 = n9903 & n9909;
  assign n9911 = ~n9894 & n9910;
  assign n9430 = x644 ^ x643;
  assign n9847 = x645 & x646;
  assign n9848 = x647 & x648;
  assign n9849 = ~n9847 & ~n9848;
  assign n9850 = ~x645 & ~x646;
  assign n9851 = ~x647 & ~x648;
  assign n9852 = ~n9850 & ~n9851;
  assign n9853 = n9849 & ~n9852;
  assign n9854 = ~n9430 & n9853;
  assign n9855 = n9847 & n9848;
  assign n9856 = n9850 & n9851;
  assign n9857 = ~n9855 & ~n9856;
  assign n9858 = ~n9854 & n9857;
  assign n9859 = x643 & x644;
  assign n9860 = ~n9858 & ~n9859;
  assign n9861 = ~n9855 & n9859;
  assign n9862 = n9861 ^ n9852;
  assign n9863 = n9861 ^ n9430;
  assign n9864 = n9852 ^ n9849;
  assign n9865 = n9864 ^ n9861;
  assign n9866 = ~n9861 & ~n9865;
  assign n9867 = n9866 ^ n9861;
  assign n9868 = n9863 & ~n9867;
  assign n9869 = n9868 ^ n9866;
  assign n9870 = n9869 ^ n9861;
  assign n9871 = n9870 ^ n9864;
  assign n9872 = n9862 & ~n9871;
  assign n9873 = n9872 ^ n9861;
  assign n9874 = ~n9860 & ~n9873;
  assign n9912 = n9911 ^ n9874;
  assign n9420 = n9419 ^ n9418;
  assign n9417 = x636 ^ x635;
  assign n9421 = n9420 ^ n9417;
  assign n9429 = x648 ^ x647;
  assign n9431 = n9430 ^ n9429;
  assign n9428 = x646 ^ x645;
  assign n9432 = n9431 ^ n9428;
  assign n9412 = x642 ^ x641;
  assign n9416 = n9415 ^ n9412;
  assign n9842 = n9432 ^ n9416;
  assign n9427 = n9426 ^ n9423;
  assign n9844 = n9842 ^ n9427;
  assign n9845 = ~n9421 & n9844;
  assign n9433 = n9432 ^ n9427;
  assign n9843 = ~n9433 & ~n9842;
  assign n9846 = n9845 ^ n9843;
  assign n9913 = n9912 ^ n9846;
  assign n9996 = n9995 ^ n9913;
  assign n10130 = n10129 ^ n9996;
  assign n9422 = n9421 ^ n9416;
  assign n9434 = n9433 ^ n9422;
  assign n9457 = n9456 ^ n9445;
  assign n9513 = n9434 & n9457;
  assign n11136 = n9996 ^ n9513;
  assign n11137 = n10130 & n11136;
  assign n11138 = n11137 ^ n10129;
  assign n11162 = n11161 ^ n11138;
  assign n11120 = ~n9416 & ~n9421;
  assign n11121 = n9913 & ~n11120;
  assign n11106 = n9416 & n9421;
  assign n11122 = n11121 ^ n11106;
  assign n11123 = ~n9995 & ~n11122;
  assign n11124 = n11123 ^ n11106;
  assign n11125 = ~n9427 & ~n9432;
  assign n11113 = n9427 & n9432;
  assign n11126 = n11125 ^ n11113;
  assign n11127 = n11126 ^ n11113;
  assign n11128 = n11113 ^ n9996;
  assign n11129 = n11128 ^ n11113;
  assign n11130 = ~n11127 & n11129;
  assign n11131 = n11130 ^ n11113;
  assign n11132 = ~n9912 & ~n11131;
  assign n11133 = n11132 ^ n11113;
  assign n11134 = ~n11124 & ~n11133;
  assign n11114 = n9912 & ~n11113;
  assign n11115 = ~n9874 & ~n9911;
  assign n11116 = ~n11114 & ~n11115;
  assign n11111 = ~n9855 & ~n9873;
  assign n11110 = ~n9888 & n9903;
  assign n11112 = n11111 ^ n11110;
  assign n11117 = n11116 ^ n11112;
  assign n11107 = n9995 & n11106;
  assign n11108 = n9958 & n9994;
  assign n11109 = ~n11107 & ~n11108;
  assign n11118 = n11117 ^ n11109;
  assign n11104 = n9975 & ~n9979;
  assign n11103 = ~n9927 & n9948;
  assign n11105 = n11104 ^ n11103;
  assign n11119 = n11118 ^ n11105;
  assign n11135 = n11134 ^ n11119;
  assign n11198 = n11138 ^ n11135;
  assign n11199 = ~n11162 & ~n11198;
  assign n11200 = n11199 ^ n11161;
  assign n11216 = n11215 ^ n11200;
  assign n11179 = n11109 & ~n11117;
  assign n11180 = n11179 ^ n11109;
  assign n11181 = ~n11134 & ~n11180;
  assign n11182 = n11181 ^ n11109;
  assign n11183 = n11105 & n11182;
  assign n11184 = n11103 & n11104;
  assign n11185 = ~n11117 & ~n11184;
  assign n11186 = n11119 & n11185;
  assign n11187 = ~n11183 & ~n11186;
  assign n11188 = ~n11118 & ~n11134;
  assign n11189 = n11188 ^ n11103;
  assign n11190 = n11189 ^ n11188;
  assign n11191 = ~n11179 & ~n11188;
  assign n11192 = n11191 ^ n11188;
  assign n11193 = n11190 & n11192;
  assign n11194 = n11193 ^ n11188;
  assign n11195 = ~n11105 & n11194;
  assign n11196 = n11187 & ~n11195;
  assign n11176 = n11116 ^ n11111;
  assign n11177 = ~n11112 & ~n11176;
  assign n11178 = n11177 ^ n11116;
  assign n11197 = n11196 ^ n11178;
  assign n11621 = n11200 ^ n11197;
  assign n11622 = n11216 & n11621;
  assign n11623 = n11622 ^ n11215;
  assign n9749 = x561 & x562;
  assign n9750 = x563 & x564;
  assign n9751 = ~n9749 & ~n9750;
  assign n9752 = ~x561 & ~x562;
  assign n9753 = ~x563 & ~x564;
  assign n9754 = ~n9752 & ~n9753;
  assign n9755 = n9751 & ~n9754;
  assign n9756 = n9749 & n9750;
  assign n9757 = x559 & x560;
  assign n9758 = ~n9756 & n9757;
  assign n9759 = ~n9755 & n9758;
  assign n9760 = n9750 ^ n9749;
  assign n9761 = n9754 ^ n9750;
  assign n9762 = n9761 ^ n9750;
  assign n9495 = x560 ^ x559;
  assign n9763 = n9750 ^ n9495;
  assign n9764 = n9763 ^ n9750;
  assign n9765 = n9762 & n9764;
  assign n9766 = n9765 ^ n9750;
  assign n9767 = n9760 & ~n9766;
  assign n9768 = n9767 ^ n9749;
  assign n9769 = ~n9759 & ~n9768;
  assign n9724 = x569 & x570;
  assign n9730 = x567 & x568;
  assign n9731 = n9724 & n9730;
  assign n9725 = ~x567 & ~x568;
  assign n9726 = ~n9724 & n9725;
  assign n9727 = ~x569 & ~x570;
  assign n9733 = n9727 & ~n9730;
  assign n9737 = ~n9726 & ~n9733;
  assign n9738 = x565 & x566;
  assign n9739 = ~n9731 & n9738;
  assign n9740 = n9737 & n9739;
  assign n9500 = x566 ^ x565;
  assign n9741 = n9724 & ~n9725;
  assign n9742 = ~n9727 & n9730;
  assign n9743 = ~n9741 & ~n9742;
  assign n9744 = n9500 & ~n9743;
  assign n9745 = ~n9740 & ~n9744;
  assign n11071 = ~n9731 & n9745;
  assign n11260 = ~n9769 & ~n11071;
  assign n9728 = x566 & ~n9727;
  assign n9729 = n9726 & ~n9728;
  assign n9732 = ~n9729 & ~n9731;
  assign n9734 = ~x566 & n9733;
  assign n9735 = n9732 & ~n9734;
  assign n9736 = ~x565 & ~n9735;
  assign n9746 = n9725 & n9734;
  assign n9747 = n9745 & ~n9746;
  assign n9748 = ~n9736 & n9747;
  assign n9770 = n9753 ^ n9752;
  assign n9771 = n9753 ^ n9751;
  assign n9772 = n9771 ^ n9753;
  assign n9773 = n9753 ^ n9495;
  assign n9774 = n9773 ^ n9753;
  assign n9775 = n9772 & ~n9774;
  assign n9776 = n9775 ^ n9753;
  assign n9777 = n9770 & ~n9776;
  assign n9778 = n9777 ^ n9752;
  assign n9779 = n9769 & ~n9778;
  assign n9780 = n9757 & ~n9759;
  assign n9781 = ~n9779 & ~n9780;
  assign n11082 = n9748 & ~n9781;
  assign n9494 = x564 ^ x563;
  assign n9496 = n9495 ^ n9494;
  assign n9493 = x562 ^ x561;
  assign n9497 = n9496 ^ n9493;
  assign n9499 = x568 ^ x567;
  assign n9501 = n9500 ^ n9499;
  assign n9498 = x570 ^ x569;
  assign n9502 = n9501 ^ n9498;
  assign n11083 = n9497 & n9502;
  assign n11084 = ~n11082 & ~n11083;
  assign n9813 = x579 & x580;
  assign n9814 = x581 & x582;
  assign n9815 = ~n9813 & ~n9814;
  assign n9816 = ~x579 & ~x580;
  assign n9817 = ~x581 & ~x582;
  assign n9818 = ~n9816 & ~n9817;
  assign n9819 = ~n9815 & n9818;
  assign n9820 = x578 & n9819;
  assign n9821 = n9813 & n9814;
  assign n9822 = ~n9820 & ~n9821;
  assign n9823 = n9815 & ~n9818;
  assign n9824 = ~x578 & n9823;
  assign n9825 = n9822 & ~n9824;
  assign n9826 = ~x577 & ~n9825;
  assign n9489 = x578 ^ x577;
  assign n9827 = n9816 & n9817;
  assign n9828 = n9489 & n9827;
  assign n9829 = n9819 ^ x578;
  assign n9830 = n9829 ^ n9819;
  assign n9831 = ~n9821 & ~n9823;
  assign n9832 = n9831 ^ n9819;
  assign n9833 = n9830 & n9832;
  assign n9834 = n9833 ^ n9819;
  assign n9835 = x577 & n9834;
  assign n9836 = ~n9828 & ~n9835;
  assign n9837 = ~n9826 & n9836;
  assign n9788 = x573 & x574;
  assign n9789 = x575 & x576;
  assign n9790 = ~n9788 & ~n9789;
  assign n9791 = ~x573 & ~x574;
  assign n9792 = ~x575 & ~x576;
  assign n9793 = ~n9791 & ~n9792;
  assign n9794 = ~n9790 & n9793;
  assign n9795 = x572 & n9794;
  assign n9796 = n9788 & n9789;
  assign n9797 = ~n9795 & ~n9796;
  assign n9798 = n9790 & ~n9793;
  assign n9799 = ~x572 & n9798;
  assign n9800 = n9797 & ~n9799;
  assign n9801 = ~x571 & ~n9800;
  assign n9484 = x572 ^ x571;
  assign n9802 = n9791 & n9792;
  assign n9803 = n9484 & n9802;
  assign n9804 = n9794 ^ x572;
  assign n9805 = n9804 ^ n9794;
  assign n9806 = ~n9796 & ~n9798;
  assign n9807 = n9806 ^ n9794;
  assign n9808 = n9805 & n9807;
  assign n9809 = n9808 ^ n9794;
  assign n9810 = x571 & n9809;
  assign n9811 = ~n9803 & ~n9810;
  assign n9812 = ~n9801 & n9811;
  assign n9838 = n9837 ^ n9812;
  assign n9503 = n9502 ^ n9497;
  assign n9488 = x580 ^ x579;
  assign n9490 = n9489 ^ n9488;
  assign n9487 = x582 ^ x581;
  assign n9491 = n9490 ^ n9487;
  assign n9483 = x574 ^ x573;
  assign n9485 = n9484 ^ n9483;
  assign n9482 = x576 ^ x575;
  assign n9486 = n9485 ^ n9482;
  assign n9492 = n9491 ^ n9486;
  assign n9504 = n9503 ^ n9492;
  assign n11076 = n9486 & n9491;
  assign n11085 = ~n9497 & ~n11076;
  assign n11086 = n9504 & n11085;
  assign n11087 = ~n9486 & ~n9491;
  assign n11088 = ~n11086 & ~n11087;
  assign n11089 = n11088 ^ n11076;
  assign n11090 = ~n9838 & ~n11089;
  assign n11091 = n11090 ^ n11076;
  assign n11092 = n11084 & n11091;
  assign n9783 = n9502 ^ n9486;
  assign n9785 = n9783 ^ n9497;
  assign n9786 = ~n9491 & n9785;
  assign n9784 = ~n9503 & ~n9783;
  assign n9787 = n9786 ^ n9784;
  assign n9839 = n9838 ^ n9787;
  assign n11093 = ~n9748 & n9781;
  assign n11094 = ~n9839 & n11093;
  assign n11095 = ~n11092 & ~n11094;
  assign n11077 = n9838 & n11076;
  assign n11078 = n9812 & n9837;
  assign n11079 = ~n11077 & ~n11078;
  assign n11074 = n9797 & ~n9810;
  assign n11073 = n9822 & ~n9835;
  assign n11075 = n11074 ^ n11073;
  assign n11080 = n11079 ^ n11075;
  assign n11242 = n11095 ^ n11080;
  assign n11096 = n9839 & n11082;
  assign n11097 = ~n11091 & n11096;
  assign n11243 = n9769 & ~n11097;
  assign n11244 = n11243 ^ n11080;
  assign n11245 = ~n11242 & ~n11244;
  assign n11246 = n11245 ^ n11095;
  assign n11239 = n11079 ^ n11074;
  assign n11240 = ~n11075 & n11239;
  assign n11241 = n11240 ^ n11079;
  assign n11247 = n11246 ^ n11241;
  assign n11248 = n9756 & n11075;
  assign n11249 = n11097 & n11248;
  assign n11250 = n11071 & ~n11249;
  assign n11251 = ~n11247 & n11250;
  assign n11098 = n11095 & ~n11097;
  assign n11252 = ~n11071 & n11241;
  assign n11253 = n11098 & n11252;
  assign n11254 = n11080 & ~n11095;
  assign n11255 = ~n11241 & n11254;
  assign n11256 = ~n11253 & ~n11255;
  assign n11257 = n9769 & ~n11256;
  assign n11258 = ~n11080 & n11095;
  assign n11259 = ~n11241 & ~n11258;
  assign n11261 = ~n11253 & n11260;
  assign n11262 = ~n11259 & n11261;
  assign n11263 = ~n11242 & n11252;
  assign n11264 = ~n11262 & ~n11263;
  assign n11265 = ~n11257 & n11264;
  assign n11266 = ~n11251 & n11265;
  assign n11626 = ~n11260 & ~n11266;
  assign n11627 = n11241 & ~n11258;
  assign n11628 = ~n11626 & ~n11627;
  assign n9538 = x605 & x606;
  assign n9537 = x603 & x604;
  assign n9539 = n9538 ^ n9537;
  assign n9540 = ~x605 & ~x606;
  assign n9541 = ~x603 & ~x604;
  assign n9542 = ~n9540 & ~n9541;
  assign n9543 = n9542 ^ n9537;
  assign n9544 = n9543 ^ n9537;
  assign n9545 = n9537 ^ x602;
  assign n9546 = n9545 ^ n9537;
  assign n9547 = n9544 & n9546;
  assign n9548 = n9547 ^ n9537;
  assign n9549 = n9539 & ~n9548;
  assign n9550 = n9549 ^ n9538;
  assign n9466 = x602 ^ x601;
  assign n9552 = ~n9537 & ~n9538;
  assign n9563 = n9542 & ~n9552;
  assign n9564 = n9466 & n9563;
  assign n9565 = ~n9542 & n9552;
  assign n9566 = x601 & x602;
  assign n9567 = n9537 & n9566;
  assign n9568 = x606 & n9567;
  assign n9569 = n9568 ^ n9566;
  assign n9570 = ~n9565 & n9569;
  assign n9571 = ~n9564 & ~n9570;
  assign n11046 = ~n9550 & n9571;
  assign n9583 = x599 & x600;
  assign n9582 = x597 & x598;
  assign n9584 = n9583 ^ n9582;
  assign n9585 = ~x599 & ~x600;
  assign n9586 = ~x597 & ~x598;
  assign n9587 = ~n9585 & ~n9586;
  assign n9588 = n9587 ^ n9582;
  assign n9589 = n9588 ^ n9582;
  assign n9590 = n9582 ^ x596;
  assign n9591 = n9590 ^ n9582;
  assign n9592 = n9589 & n9591;
  assign n9593 = n9592 ^ n9582;
  assign n9594 = n9584 & ~n9593;
  assign n9595 = n9594 ^ n9583;
  assign n9461 = x596 ^ x595;
  assign n9597 = ~n9582 & ~n9583;
  assign n9608 = n9587 & ~n9597;
  assign n9609 = n9461 & n9608;
  assign n9610 = ~n9587 & n9597;
  assign n9611 = x595 & x596;
  assign n9612 = n9582 & n9611;
  assign n9613 = x600 & n9612;
  assign n9614 = n9613 ^ n9611;
  assign n9615 = ~n9610 & n9614;
  assign n9616 = ~n9609 & ~n9615;
  assign n11045 = ~n9595 & n9616;
  assign n11047 = n11046 ^ n11045;
  assign n9596 = n9586 ^ n9585;
  assign n9598 = n9597 ^ n9586;
  assign n9599 = n9598 ^ n9586;
  assign n9600 = n9586 ^ x596;
  assign n9601 = n9600 ^ n9586;
  assign n9602 = n9599 & ~n9601;
  assign n9603 = n9602 ^ n9586;
  assign n9604 = n9596 & ~n9603;
  assign n9605 = n9604 ^ n9585;
  assign n9606 = ~n9595 & ~n9605;
  assign n9607 = ~x595 & ~n9606;
  assign n9460 = x598 ^ x597;
  assign n9617 = n9611 ^ x598;
  assign n9618 = n9617 ^ n9611;
  assign n9619 = ~x596 & ~x600;
  assign n9620 = n9619 ^ n9611;
  assign n9621 = ~n9618 & n9620;
  assign n9622 = n9621 ^ n9611;
  assign n9623 = ~n9460 & n9622;
  assign n9624 = ~x599 & n9623;
  assign n9625 = n9616 & ~n9624;
  assign n9626 = ~n9607 & n9625;
  assign n9551 = n9541 ^ n9540;
  assign n9553 = n9552 ^ n9541;
  assign n9554 = n9553 ^ n9541;
  assign n9555 = n9541 ^ x602;
  assign n9556 = n9555 ^ n9541;
  assign n9557 = n9554 & ~n9556;
  assign n9558 = n9557 ^ n9541;
  assign n9559 = n9551 & ~n9558;
  assign n9560 = n9559 ^ n9540;
  assign n9561 = ~n9550 & ~n9560;
  assign n9562 = ~x601 & ~n9561;
  assign n9465 = x604 ^ x603;
  assign n9572 = n9566 ^ x604;
  assign n9573 = n9572 ^ n9566;
  assign n9574 = ~x602 & ~x606;
  assign n9575 = n9574 ^ n9566;
  assign n9576 = ~n9573 & n9575;
  assign n9577 = n9576 ^ n9566;
  assign n9578 = ~n9465 & n9577;
  assign n9579 = ~x605 & n9578;
  assign n9580 = n9571 & ~n9579;
  assign n9581 = ~n9562 & n9580;
  assign n9627 = n9626 ^ n9581;
  assign n9462 = n9461 ^ n9460;
  assign n9459 = x600 ^ x599;
  assign n9463 = n9462 ^ n9459;
  assign n9467 = n9466 ^ n9465;
  assign n9464 = x606 ^ x605;
  assign n9468 = n9467 ^ n9464;
  assign n9517 = n9463 & n9468;
  assign n11042 = n9581 ^ n9517;
  assign n11043 = n9627 & ~n11042;
  assign n11044 = n11043 ^ n9626;
  assign n11048 = n11047 ^ n11044;
  assign n9472 = x586 ^ x585;
  assign n9471 = x588 ^ x587;
  assign n9473 = n9472 ^ n9471;
  assign n9470 = x584 ^ x583;
  assign n9474 = n9473 ^ n9470;
  assign n9477 = x590 ^ x589;
  assign n9476 = x592 ^ x591;
  assign n9478 = n9477 ^ n9476;
  assign n9475 = x594 ^ x593;
  assign n9479 = n9478 ^ n9475;
  assign n9527 = n9474 & n9479;
  assign n9681 = x591 & x592;
  assign n9680 = x593 & x594;
  assign n9682 = n9681 ^ n9680;
  assign n9683 = ~x591 & ~x592;
  assign n9684 = ~x593 & ~x594;
  assign n9685 = ~n9683 & ~n9684;
  assign n9686 = n9685 ^ n9680;
  assign n9687 = n9686 ^ n9680;
  assign n9688 = n9680 ^ x590;
  assign n9689 = n9688 ^ n9680;
  assign n9690 = n9687 & n9689;
  assign n9691 = n9690 ^ n9680;
  assign n9692 = n9682 & ~n9691;
  assign n9693 = n9692 ^ n9681;
  assign n9694 = x593 ^ x590;
  assign n9695 = n9475 & n9694;
  assign n9696 = n9695 ^ x593;
  assign n9697 = n9683 & ~n9696;
  assign n9698 = ~n9693 & ~n9697;
  assign n9699 = ~x589 & ~n9698;
  assign n9700 = x589 & x590;
  assign n9701 = n9700 ^ n9478;
  assign n9702 = n9701 ^ n9700;
  assign n9703 = ~x590 & ~x594;
  assign n9704 = n9703 ^ n9700;
  assign n9705 = n9704 ^ n9700;
  assign n9706 = n9702 & n9705;
  assign n9707 = n9706 ^ n9700;
  assign n9708 = ~n9681 & n9707;
  assign n9709 = n9708 ^ n9700;
  assign n9710 = ~x593 & n9709;
  assign n9711 = ~n9680 & ~n9681;
  assign n9712 = ~n9685 & n9711;
  assign n9713 = n9681 & n9700;
  assign n9714 = x594 & n9713;
  assign n9715 = n9714 ^ n9700;
  assign n9716 = ~n9712 & n9715;
  assign n9717 = n9685 & ~n9711;
  assign n9718 = n9477 & n9717;
  assign n9719 = ~n9716 & ~n9718;
  assign n9720 = ~n9710 & n9719;
  assign n9721 = ~n9699 & n9720;
  assign n9629 = x583 & x584;
  assign n9630 = n9629 ^ x586;
  assign n9631 = n9630 ^ n9629;
  assign n9632 = ~x584 & ~x588;
  assign n9633 = n9632 ^ n9629;
  assign n9634 = ~n9631 & n9633;
  assign n9635 = n9634 ^ n9629;
  assign n9636 = ~n9472 & n9635;
  assign n9637 = ~x587 & n9636;
  assign n9639 = x585 & x586;
  assign n9638 = x587 & x588;
  assign n9640 = n9639 ^ n9638;
  assign n9641 = ~x585 & ~x586;
  assign n9642 = ~x587 & ~x588;
  assign n9643 = ~n9641 & ~n9642;
  assign n9644 = n9643 ^ n9638;
  assign n9645 = n9644 ^ n9638;
  assign n9646 = n9638 ^ x584;
  assign n9647 = n9646 ^ n9638;
  assign n9648 = n9645 & n9647;
  assign n9649 = n9648 ^ n9638;
  assign n9650 = n9640 & ~n9649;
  assign n9651 = n9650 ^ n9639;
  assign n9652 = n9642 ^ n9641;
  assign n9653 = ~n9638 & ~n9639;
  assign n9654 = n9653 ^ n9642;
  assign n9655 = n9654 ^ n9642;
  assign n9656 = n9642 ^ x584;
  assign n9657 = n9656 ^ n9642;
  assign n9658 = n9655 & ~n9657;
  assign n9659 = n9658 ^ n9642;
  assign n9660 = n9652 & ~n9659;
  assign n9661 = n9660 ^ n9641;
  assign n9662 = ~n9651 & ~n9661;
  assign n9663 = n9662 ^ x583;
  assign n9664 = n9663 ^ n9662;
  assign n9666 = n9643 & ~n9653;
  assign n9665 = x588 & n9639;
  assign n9667 = n9666 ^ n9665;
  assign n9668 = n9667 ^ n9666;
  assign n9669 = ~n9643 & n9653;
  assign n9670 = n9669 ^ n9666;
  assign n9671 = n9670 ^ n9666;
  assign n9672 = ~n9668 & ~n9671;
  assign n9673 = n9672 ^ n9666;
  assign n9674 = x584 & n9673;
  assign n9675 = n9674 ^ n9666;
  assign n9676 = n9675 ^ n9662;
  assign n9677 = n9664 & ~n9676;
  assign n9678 = n9677 ^ n9662;
  assign n9679 = ~n9637 & n9678;
  assign n9722 = n9721 ^ n9679;
  assign n11058 = ~n9527 & ~n9722;
  assign n9469 = n9468 ^ n9463;
  assign n9480 = n9479 ^ n9474;
  assign n11059 = n9480 ^ n9463;
  assign n11060 = n9469 & ~n11059;
  assign n11061 = n11060 ^ n9468;
  assign n11062 = ~n9627 & n11061;
  assign n11063 = ~n11058 & n11062;
  assign n11064 = ~n9517 & n9627;
  assign n11065 = ~n11063 & ~n11064;
  assign n9525 = ~n9474 & ~n9479;
  assign n9526 = ~n9517 & n9525;
  assign n9518 = ~n9463 & ~n9468;
  assign n9528 = n9518 & ~n9527;
  assign n9529 = ~n9526 & ~n9528;
  assign n11066 = n9529 ^ n9527;
  assign n11067 = ~n9722 & ~n11066;
  assign n11068 = n11067 ^ n9527;
  assign n11069 = ~n11065 & ~n11068;
  assign n11225 = ~n11048 & ~n11069;
  assign n11050 = x583 & n9675;
  assign n11051 = ~n9651 & ~n11050;
  assign n11049 = ~n9693 & n9719;
  assign n11052 = n11051 ^ n11049;
  assign n11053 = ~n9527 & n9722;
  assign n11054 = ~n9679 & ~n9721;
  assign n11055 = ~n11053 & ~n11054;
  assign n11226 = n11055 ^ n11051;
  assign n11227 = ~n11052 & ~n11226;
  assign n11228 = n11227 ^ n11055;
  assign n11229 = n11225 & ~n11228;
  assign n11056 = n11055 ^ n11052;
  assign n11057 = n11056 ^ n11048;
  assign n11070 = n11069 ^ n11057;
  assign n11230 = n11049 & n11051;
  assign n11231 = ~n11055 & n11230;
  assign n11232 = n11070 & n11231;
  assign n11233 = ~n11229 & ~n11232;
  assign n11234 = n11048 & n11228;
  assign n11235 = ~n11070 & n11234;
  assign n11236 = n11233 & ~n11235;
  assign n11222 = n11046 ^ n11044;
  assign n11223 = ~n11047 & ~n11222;
  assign n11224 = n11223 ^ n11044;
  assign n11237 = n11236 ^ n11224;
  assign n11072 = n11071 ^ n9769;
  assign n11081 = n11080 ^ n11072;
  assign n11099 = n11098 ^ n11081;
  assign n11100 = n11099 ^ n11070;
  assign n9519 = n9518 ^ n9517;
  assign n9520 = n9517 ^ n9474;
  assign n9521 = n9480 & ~n9520;
  assign n9522 = n9521 ^ n9474;
  assign n9523 = n9519 & n9522;
  assign n9524 = n9523 ^ n9518;
  assign n9530 = n9529 ^ n9504;
  assign n9531 = n9530 ^ n9504;
  assign n9481 = n9480 ^ n9469;
  assign n9532 = n9481 & n9504;
  assign n9533 = n9532 ^ n9504;
  assign n9534 = n9531 & ~n9533;
  assign n9535 = n9534 ^ n9504;
  assign n9536 = ~n9524 & n9535;
  assign n9628 = n9627 ^ n9536;
  assign n9723 = n9722 ^ n9628;
  assign n9782 = n9781 ^ n9748;
  assign n9840 = n9839 ^ n9782;
  assign n11039 = n9840 ^ n9532;
  assign n11040 = ~n9723 & n11039;
  assign n11041 = n11040 ^ n9840;
  assign n11219 = n11070 ^ n11041;
  assign n11220 = ~n11100 & ~n11219;
  assign n11221 = n11220 ^ n11099;
  assign n11238 = n11237 ^ n11221;
  assign n11629 = n11266 ^ n11221;
  assign n11630 = n11238 & n11629;
  assign n11631 = n11630 ^ n11266;
  assign n11632 = ~n11628 & n11631;
  assign n11633 = n11221 & n11266;
  assign n11634 = n11237 & ~n11633;
  assign n11635 = n11628 & n11634;
  assign n11636 = ~n11632 & ~n11635;
  assign n11624 = ~n11224 & ~n11235;
  assign n11625 = n11233 & ~n11624;
  assign n11637 = n11636 ^ n11625;
  assign n11767 = ~n11623 & ~n11637;
  assign n11615 = ~n11103 & ~n11104;
  assign n11616 = ~n11197 & ~n11615;
  assign n11617 = ~n11178 & ~n11191;
  assign n11618 = ~n11616 & ~n11617;
  assign n11613 = ~n11203 & ~n11208;
  assign n11614 = ~n11213 & ~n11613;
  assign n11619 = n11618 ^ n11614;
  assign n11217 = n11216 ^ n11197;
  assign n11163 = n11162 ^ n11135;
  assign n11101 = n11100 ^ n11041;
  assign n11172 = n11163 ^ n11101;
  assign n11034 = n9513 & n10130;
  assign n9841 = n9840 ^ n9723;
  assign n10131 = n10130 ^ n9841;
  assign n9458 = n9457 ^ n9434;
  assign n9505 = n9504 ^ n9481;
  assign n9506 = n9505 ^ n9434;
  assign n9507 = n9458 & ~n9506;
  assign n9508 = n9507 ^ n9457;
  assign n11035 = n10130 ^ n9508;
  assign n11036 = n10131 & n11035;
  assign n11037 = n11036 ^ n10130;
  assign n11038 = ~n11034 & n11037;
  assign n11173 = n11163 ^ n11038;
  assign n11174 = ~n11172 & ~n11173;
  assign n11175 = n11174 ^ n11101;
  assign n11218 = n11217 ^ n11175;
  assign n11267 = n11266 ^ n11238;
  assign n11610 = n11267 ^ n11175;
  assign n11611 = n11218 & n11610;
  assign n11612 = n11611 ^ n11217;
  assign n11768 = n11618 ^ n11612;
  assign n11769 = ~n11619 & ~n11768;
  assign n11770 = n11769 ^ n11612;
  assign n11771 = n11767 & n11770;
  assign n11772 = ~n11614 & ~n11618;
  assign n11773 = n11612 & n11772;
  assign n11638 = n11637 ^ n11623;
  assign n11620 = n11619 ^ n11612;
  assign n11639 = n11638 ^ n11620;
  assign n11774 = n11612 & ~n11623;
  assign n11775 = n11639 & ~n11774;
  assign n11776 = n11773 & ~n11775;
  assign n11777 = ~n11771 & ~n11776;
  assign n11778 = n11637 & ~n11770;
  assign n11779 = n11639 & n11778;
  assign n11780 = n11777 & ~n11779;
  assign n11765 = ~n11625 & ~n11635;
  assign n11766 = ~n11632 & ~n11765;
  assign n11781 = n11780 ^ n11766;
  assign n10616 = x515 & x516;
  assign n10617 = x513 & x514;
  assign n10618 = ~n10616 & ~n10617;
  assign n10619 = ~x515 & ~x516;
  assign n10620 = ~x513 & ~x514;
  assign n10621 = ~n10619 & ~n10620;
  assign n10622 = ~n10618 & n10621;
  assign n10623 = x512 & n10622;
  assign n10624 = n10616 & n10617;
  assign n10625 = ~n10623 & ~n10624;
  assign n10632 = n10622 ^ x512;
  assign n10633 = n10632 ^ n10622;
  assign n10626 = n10618 & ~n10621;
  assign n10634 = ~n10624 & ~n10626;
  assign n10635 = n10634 ^ n10622;
  assign n10636 = n10633 & n10635;
  assign n10637 = n10636 ^ n10622;
  assign n10638 = x511 & n10637;
  assign n10984 = n10625 & ~n10638;
  assign n10591 = x521 & x522;
  assign n10592 = x519 & x520;
  assign n10593 = ~n10591 & ~n10592;
  assign n10594 = ~x521 & ~x522;
  assign n10595 = ~x519 & ~x520;
  assign n10596 = ~n10594 & ~n10595;
  assign n10597 = ~n10593 & n10596;
  assign n10598 = x518 & n10597;
  assign n10599 = n10591 & n10592;
  assign n10600 = ~n10598 & ~n10599;
  assign n10607 = n10597 ^ x518;
  assign n10608 = n10607 ^ n10597;
  assign n10601 = n10593 & ~n10596;
  assign n10609 = ~n10599 & ~n10601;
  assign n10610 = n10609 ^ n10597;
  assign n10611 = n10608 & n10610;
  assign n10612 = n10611 ^ n10597;
  assign n10613 = x517 & n10612;
  assign n10985 = n10600 & ~n10613;
  assign n11348 = ~n10984 & ~n10985;
  assign n10627 = ~x512 & n10626;
  assign n10628 = n10625 & ~n10627;
  assign n10629 = ~x511 & ~n10628;
  assign n9389 = x512 ^ x511;
  assign n10630 = n10619 & n10620;
  assign n10631 = n9389 & n10630;
  assign n10639 = ~n10631 & ~n10638;
  assign n10640 = ~n10629 & n10639;
  assign n10602 = ~x518 & n10601;
  assign n10603 = n10600 & ~n10602;
  assign n10604 = ~x517 & ~n10603;
  assign n9394 = x518 ^ x517;
  assign n10605 = n10594 & n10595;
  assign n10606 = n9394 & n10605;
  assign n10614 = ~n10606 & ~n10613;
  assign n10615 = ~n10604 & n10614;
  assign n10641 = n10640 ^ n10615;
  assign n9388 = x514 ^ x513;
  assign n9390 = n9389 ^ n9388;
  assign n9387 = x516 ^ x515;
  assign n9391 = n9390 ^ n9387;
  assign n9393 = x520 ^ x519;
  assign n9395 = n9394 ^ n9393;
  assign n9392 = x522 ^ x521;
  assign n9396 = n9395 ^ n9392;
  assign n10587 = n9391 & n9396;
  assign n10981 = n10615 ^ n10587;
  assign n10982 = n10641 & ~n10981;
  assign n10983 = n10982 ^ n10640;
  assign n9397 = n9396 ^ n9391;
  assign n9405 = x530 ^ x529;
  assign n9404 = x532 ^ x531;
  assign n9406 = n9405 ^ n9404;
  assign n9403 = x534 ^ x533;
  assign n9407 = n9406 ^ n9403;
  assign n9400 = x524 ^ x523;
  assign n9399 = x526 ^ x525;
  assign n9401 = n9400 ^ n9399;
  assign n9398 = x528 ^ x527;
  assign n9402 = n9401 ^ n9398;
  assign n9408 = n9407 ^ n9402;
  assign n10584 = n9408 ^ n9396;
  assign n10585 = ~n9397 & n10584;
  assign n10586 = n10585 ^ n9408;
  assign n10996 = ~n10586 & ~n10641;
  assign n10997 = n10587 & n10641;
  assign n10583 = n9402 & n9407;
  assign n10588 = n10587 ^ n10586;
  assign n10589 = ~n10583 & ~n10588;
  assign n10590 = n10589 ^ n10587;
  assign n10642 = n10641 ^ n10590;
  assign n10557 = x527 & x528;
  assign n10558 = x525 & x526;
  assign n10559 = ~n10557 & ~n10558;
  assign n10560 = ~x527 & ~x528;
  assign n10561 = ~x525 & ~x526;
  assign n10562 = ~n10560 & ~n10561;
  assign n10563 = ~n10559 & n10562;
  assign n10564 = x524 & n10563;
  assign n10565 = n10557 & n10558;
  assign n10566 = ~n10564 & ~n10565;
  assign n10567 = n10559 & ~n10562;
  assign n10568 = ~x524 & n10567;
  assign n10569 = n10566 & ~n10568;
  assign n10570 = ~x523 & ~n10569;
  assign n10571 = n10560 & n10561;
  assign n10572 = n9400 & n10571;
  assign n10573 = n10563 ^ x524;
  assign n10574 = n10573 ^ n10563;
  assign n10575 = ~n10565 & ~n10567;
  assign n10576 = n10575 ^ n10563;
  assign n10577 = n10574 & n10576;
  assign n10578 = n10577 ^ n10563;
  assign n10579 = x523 & n10578;
  assign n10580 = ~n10572 & ~n10579;
  assign n10581 = ~n10570 & n10580;
  assign n10532 = x531 & x532;
  assign n10533 = x533 & x534;
  assign n10534 = ~n10532 & ~n10533;
  assign n10535 = ~x531 & ~x532;
  assign n10536 = ~x533 & ~x534;
  assign n10537 = ~n10535 & ~n10536;
  assign n10538 = ~n10534 & n10537;
  assign n10539 = x530 & n10538;
  assign n10540 = n10532 & n10533;
  assign n10541 = ~n10539 & ~n10540;
  assign n10542 = n10534 & ~n10537;
  assign n10543 = ~x530 & n10542;
  assign n10544 = n10541 & ~n10543;
  assign n10545 = ~x529 & ~n10544;
  assign n10546 = n10535 & n10536;
  assign n10547 = n9405 & n10546;
  assign n10548 = n10538 ^ x530;
  assign n10549 = n10548 ^ n10538;
  assign n10550 = ~n10540 & ~n10542;
  assign n10551 = n10550 ^ n10538;
  assign n10552 = n10549 & n10551;
  assign n10553 = n10552 ^ n10538;
  assign n10554 = x529 & n10553;
  assign n10555 = ~n10547 & ~n10554;
  assign n10556 = ~n10545 & n10555;
  assign n10582 = n10581 ^ n10556;
  assign n10643 = n10642 ^ n10582;
  assign n10998 = n10643 ^ n10642;
  assign n10999 = n10642 ^ n10583;
  assign n11000 = n10998 & ~n10999;
  assign n11001 = n11000 ^ n10642;
  assign n11002 = ~n10997 & n11001;
  assign n11003 = ~n10996 & n11002;
  assign n11337 = n10983 & n11003;
  assign n11336 = n10984 & n10985;
  assign n11338 = n11337 ^ n11336;
  assign n10991 = n10582 & n10583;
  assign n10992 = n10556 & n10581;
  assign n10993 = ~n10991 & ~n10992;
  assign n10989 = n10566 & ~n10579;
  assign n10988 = n10541 & ~n10554;
  assign n10990 = n10989 ^ n10988;
  assign n10994 = n10993 ^ n10990;
  assign n11339 = ~n10983 & ~n11003;
  assign n11340 = ~n10994 & ~n11339;
  assign n11341 = n11340 ^ n11336;
  assign n11342 = n11341 ^ n11340;
  assign n11343 = n11340 ^ n10994;
  assign n11344 = ~n11342 & n11343;
  assign n11345 = n11344 ^ n11340;
  assign n11346 = n11338 & ~n11345;
  assign n11347 = n11339 ^ n10994;
  assign n11349 = n11348 ^ n10994;
  assign n11350 = ~n11347 & n11349;
  assign n11351 = ~n11346 & ~n11350;
  assign n11333 = n10993 ^ n10989;
  assign n11334 = ~n10990 & n11333;
  assign n11335 = n11334 ^ n10993;
  assign n11352 = n11351 ^ n11335;
  assign n11586 = ~n11348 & ~n11352;
  assign n11587 = n11335 & ~n11340;
  assign n11588 = ~n11586 & ~n11587;
  assign n10511 = x551 & x552;
  assign n10512 = x549 & x550;
  assign n10513 = n10511 & n10512;
  assign n10516 = x547 & x548;
  assign n10518 = ~n10513 & n10516;
  assign n9380 = x552 ^ x551;
  assign n10505 = x551 ^ x550;
  assign n10506 = ~n9380 & n10505;
  assign n10507 = n10506 ^ x550;
  assign n10519 = n10518 ^ n10507;
  assign n10502 = ~x551 & ~x552;
  assign n10503 = ~x550 & n10502;
  assign n10504 = x549 & ~n10503;
  assign n10520 = n10518 ^ n10504;
  assign n10521 = n10520 ^ n10504;
  assign n9381 = x550 ^ x549;
  assign n9382 = n9381 ^ n9380;
  assign n9383 = x548 ^ x547;
  assign n10522 = n9382 & n9383;
  assign n10523 = n10522 ^ n10504;
  assign n10524 = ~n10521 & ~n10523;
  assign n10525 = n10524 ^ n10504;
  assign n10526 = n10519 & n10525;
  assign n10527 = n10526 ^ n10507;
  assign n11013 = ~n10513 & ~n10527;
  assign n9376 = x556 ^ x555;
  assign n10479 = x557 & x558;
  assign n10480 = n10479 ^ x556;
  assign n10481 = ~n9376 & ~n10480;
  assign n10483 = x555 & x556;
  assign n10484 = ~x557 & ~x558;
  assign n10485 = ~n10483 & n10484;
  assign n10493 = x553 & x554;
  assign n10494 = ~n10485 & n10493;
  assign n10495 = ~n10481 & n10494;
  assign n9377 = x554 ^ x553;
  assign n10488 = ~x555 & ~x556;
  assign n10496 = n10479 & ~n10488;
  assign n10497 = n10483 & ~n10484;
  assign n10498 = ~n10496 & ~n10497;
  assign n10499 = n9377 & ~n10498;
  assign n10500 = ~n10495 & ~n10499;
  assign n11011 = n10479 & n10483;
  assign n11012 = n10500 & ~n11011;
  assign n11014 = n11013 ^ n11012;
  assign n9378 = n9377 ^ n9376;
  assign n9375 = x558 ^ x557;
  assign n9379 = n9378 ^ n9375;
  assign n9384 = n9383 ^ n9382;
  assign n10462 = n9379 & n9384;
  assign n10508 = ~n10504 & ~n10507;
  assign n10509 = ~n9383 & n10508;
  assign n10510 = ~x549 & n10503;
  assign n10514 = ~n10510 & ~n10513;
  assign n10515 = ~n10509 & n10514;
  assign n10517 = ~n10515 & ~n10516;
  assign n10528 = ~n10517 & ~n10527;
  assign n10482 = ~x553 & n10481;
  assign n10486 = ~x554 & n10485;
  assign n10487 = ~n10482 & ~n10486;
  assign n10489 = x553 & ~n10488;
  assign n10490 = x554 & ~n10484;
  assign n10491 = ~n10489 & ~n10490;
  assign n10492 = ~n10487 & n10491;
  assign n10501 = ~n10492 & n10500;
  assign n10529 = n10528 ^ n10501;
  assign n11015 = ~n10462 & n10529;
  assign n11016 = ~n10501 & ~n10528;
  assign n11017 = ~n11015 & ~n11016;
  assign n11354 = n11017 ^ n11013;
  assign n11355 = ~n11014 & ~n11354;
  assign n11356 = n11355 ^ n11017;
  assign n10402 = x539 & x540;
  assign n10403 = x537 & x538;
  assign n10404 = ~n10402 & ~n10403;
  assign n10405 = ~x539 & ~x540;
  assign n10406 = ~x537 & ~x538;
  assign n10407 = ~n10405 & ~n10406;
  assign n10408 = ~n10404 & n10407;
  assign n10409 = x536 & n10408;
  assign n10410 = n10402 & n10403;
  assign n10411 = ~n10409 & ~n10410;
  assign n10418 = n10408 ^ x536;
  assign n10419 = n10418 ^ n10408;
  assign n10412 = n10404 & ~n10407;
  assign n10420 = ~n10410 & ~n10412;
  assign n10421 = n10420 ^ n10408;
  assign n10422 = n10419 & n10421;
  assign n10423 = n10422 ^ n10408;
  assign n10424 = x535 & n10423;
  assign n11005 = n10411 & ~n10424;
  assign n10427 = x543 & x544;
  assign n10428 = ~x545 & ~x546;
  assign n10429 = ~n10427 & n10428;
  assign n10430 = x545 & x546;
  assign n10431 = ~x543 & ~x544;
  assign n10432 = ~n10430 & n10431;
  assign n10433 = ~n10429 & ~n10432;
  assign n10434 = n10427 & n10430;
  assign n10435 = n10433 & ~n10434;
  assign n10436 = x542 & ~n10435;
  assign n9370 = x544 ^ x543;
  assign n10437 = n10430 ^ x544;
  assign n10438 = n9370 & ~n10437;
  assign n10439 = n10438 ^ x543;
  assign n10440 = n10439 ^ n10428;
  assign n10441 = n10428 ^ x541;
  assign n10442 = ~n10428 & ~n10441;
  assign n10443 = n10442 ^ n10428;
  assign n10444 = ~n10440 & ~n10443;
  assign n10445 = n10444 ^ n10442;
  assign n10446 = n10445 ^ n10428;
  assign n10447 = n10446 ^ x541;
  assign n10448 = ~x542 & ~n10447;
  assign n10449 = n10448 ^ x541;
  assign n10450 = ~n10436 & n10449;
  assign n10451 = x542 & ~n10428;
  assign n10452 = ~n10434 & ~n10451;
  assign n10453 = n10439 & ~n10452;
  assign n11006 = ~n10450 & ~n10453;
  assign n11358 = ~n11005 & ~n11006;
  assign n10454 = n10432 & ~n10451;
  assign n10455 = ~n10453 & ~n10454;
  assign n10456 = ~x541 & ~n10455;
  assign n10457 = ~n10450 & ~n10456;
  assign n9371 = x546 ^ x545;
  assign n9372 = n9371 ^ n9370;
  assign n9369 = x542 ^ x541;
  assign n9373 = n9372 ^ n9369;
  assign n10458 = ~x542 & n10429;
  assign n10459 = n9373 & n10458;
  assign n10460 = n10457 & ~n10459;
  assign n10413 = ~x536 & n10412;
  assign n10414 = n10411 & ~n10413;
  assign n10415 = ~x535 & ~n10414;
  assign n9366 = x536 ^ x535;
  assign n10416 = n10405 & n10406;
  assign n10417 = n9366 & n10416;
  assign n10425 = ~n10417 & ~n10424;
  assign n10426 = ~n10415 & n10425;
  assign n10461 = n10460 ^ n10426;
  assign n9365 = x538 ^ x537;
  assign n9367 = n9366 ^ n9365;
  assign n9364 = x540 ^ x539;
  assign n9368 = n9367 ^ n9364;
  assign n10463 = n9368 & n9373;
  assign n11008 = n10463 ^ n10460;
  assign n11009 = ~n10461 & n11008;
  assign n11010 = n11009 ^ n10463;
  assign n11018 = n11017 ^ n11014;
  assign n11357 = n11010 & n11018;
  assign n11359 = n11358 ^ n11357;
  assign n10464 = n10462 & n10463;
  assign n9374 = n9373 ^ n9368;
  assign n10465 = n9384 ^ n9374;
  assign n9385 = n9384 ^ n9379;
  assign n10466 = n10465 ^ n9385;
  assign n10467 = n9379 ^ n9373;
  assign n10468 = n10467 ^ n9384;
  assign n10469 = n10468 ^ n9384;
  assign n10470 = ~n9374 & n10469;
  assign n10471 = n10470 ^ n9374;
  assign n10472 = n10468 & ~n10471;
  assign n10473 = n10472 ^ n9384;
  assign n10474 = n10466 & n10473;
  assign n10475 = n10474 ^ n10470;
  assign n10476 = n10475 ^ n9384;
  assign n10477 = n10476 ^ n9385;
  assign n10478 = ~n10464 & n10477;
  assign n10530 = n10529 ^ n10478;
  assign n11020 = ~n10461 & n10530;
  assign n11021 = n10477 ^ n10462;
  assign n11022 = ~n10529 & ~n11021;
  assign n11023 = n11022 ^ n10462;
  assign n11024 = ~n11020 & ~n11023;
  assign n11025 = n10461 & n10463;
  assign n11026 = n11024 & ~n11025;
  assign n11360 = n11357 ^ n11026;
  assign n11361 = n11360 ^ n11026;
  assign n11362 = ~n11010 & ~n11018;
  assign n11363 = n11026 & ~n11362;
  assign n11364 = n11363 ^ n11026;
  assign n11365 = ~n11361 & ~n11364;
  assign n11366 = n11365 ^ n11026;
  assign n11367 = n11359 & n11366;
  assign n11368 = n11367 ^ n11358;
  assign n11369 = ~n11356 & ~n11368;
  assign n11019 = n11018 ^ n11010;
  assign n11027 = n11026 ^ n11019;
  assign n11370 = n11005 & n11006;
  assign n11371 = n11027 & n11370;
  assign n11372 = ~n11026 & ~n11358;
  assign n11373 = n11362 & n11372;
  assign n11374 = ~n11371 & ~n11373;
  assign n11375 = ~n11369 & n11374;
  assign n11589 = n11588 ^ n11375;
  assign n11007 = n11006 ^ n11005;
  assign n11028 = n11027 ^ n11007;
  assign n10986 = n10985 ^ n10984;
  assign n10987 = n10986 ^ n10983;
  assign n10995 = n10994 ^ n10987;
  assign n11004 = n11003 ^ n10995;
  assign n11029 = n11028 ^ n11004;
  assign n10531 = n10530 ^ n10461;
  assign n10644 = n10643 ^ n10531;
  assign n9386 = n9385 ^ n9374;
  assign n9409 = n9408 ^ n9397;
  assign n10974 = n9386 & n9409;
  assign n10978 = n10974 ^ n10531;
  assign n10979 = ~n10644 & ~n10978;
  assign n10980 = n10979 ^ n10643;
  assign n11330 = n11004 ^ n10980;
  assign n11331 = ~n11029 & ~n11330;
  assign n11332 = n11331 ^ n11028;
  assign n11353 = n11352 ^ n11332;
  assign n11376 = n11018 & n11026;
  assign n11377 = n11375 & n11376;
  assign n11378 = ~n11363 & n11371;
  assign n11379 = n11357 & n11358;
  assign n11380 = ~n11373 & ~n11379;
  assign n11381 = ~n11378 & n11380;
  assign n11382 = ~n11377 & n11381;
  assign n11383 = n11382 ^ n11356;
  assign n11583 = n11383 ^ n11352;
  assign n11584 = n11353 & ~n11583;
  assign n11585 = n11584 ^ n11383;
  assign n11590 = n11589 ^ n11585;
  assign n10197 = x501 & x502;
  assign n10198 = x503 & x504;
  assign n10199 = ~n10197 & ~n10198;
  assign n10200 = ~x501 & ~x502;
  assign n10201 = ~x503 & ~x504;
  assign n10202 = ~n10200 & ~n10201;
  assign n10203 = ~n10199 & n10202;
  assign n10204 = x500 & n10203;
  assign n10205 = n10197 & n10198;
  assign n10206 = ~n10204 & ~n10205;
  assign n10213 = n10203 ^ x500;
  assign n10214 = n10213 ^ n10203;
  assign n10207 = n10199 & ~n10202;
  assign n10215 = ~n10205 & ~n10207;
  assign n10216 = n10215 ^ n10203;
  assign n10217 = n10214 & n10216;
  assign n10218 = n10217 ^ n10203;
  assign n10219 = x499 & n10218;
  assign n10954 = n10206 & ~n10219;
  assign n10230 = x509 & x510;
  assign n10231 = x508 & n10230;
  assign n10232 = x507 & n10231;
  assign n10235 = x505 & x506;
  assign n10238 = ~n10232 & n10235;
  assign n9345 = x510 ^ x509;
  assign n10225 = x509 ^ x508;
  assign n10226 = ~n9345 & n10225;
  assign n10227 = n10226 ^ x508;
  assign n10239 = n10238 ^ n10227;
  assign n10222 = ~x509 & ~x510;
  assign n10223 = ~x508 & n10222;
  assign n10224 = x507 & ~n10223;
  assign n10240 = n10238 ^ n10224;
  assign n10241 = n10240 ^ n10224;
  assign n9347 = x506 ^ x505;
  assign n10242 = ~x507 & ~n10231;
  assign n10243 = n9347 & ~n10242;
  assign n10244 = n10243 ^ n10224;
  assign n10245 = ~n10241 & ~n10244;
  assign n10246 = n10245 ^ n10224;
  assign n10247 = n10239 & n10246;
  assign n10248 = n10247 ^ n10227;
  assign n10953 = ~n10232 & ~n10248;
  assign n10955 = n10954 ^ n10953;
  assign n10228 = ~n10224 & ~n10227;
  assign n10229 = ~x506 & n10228;
  assign n10233 = ~n10229 & ~n10232;
  assign n10234 = ~x505 & ~n10233;
  assign n10236 = ~x507 & ~n10235;
  assign n10237 = n10223 & n10236;
  assign n10249 = ~n10237 & ~n10248;
  assign n10250 = ~n10234 & n10249;
  assign n10208 = ~x500 & n10207;
  assign n10209 = n10206 & ~n10208;
  assign n10210 = ~x499 & ~n10209;
  assign n9342 = x500 ^ x499;
  assign n10211 = n10200 & n10201;
  assign n10212 = n9342 & n10211;
  assign n10220 = ~n10212 & ~n10219;
  assign n10221 = ~n10210 & n10220;
  assign n10251 = n10250 ^ n10221;
  assign n9341 = x502 ^ x501;
  assign n9343 = n9342 ^ n9341;
  assign n9340 = x504 ^ x503;
  assign n9344 = n9343 ^ n9340;
  assign n9346 = x508 ^ x507;
  assign n9348 = n9347 ^ n9346;
  assign n9349 = n9348 ^ n9345;
  assign n10141 = n9344 & n9349;
  assign n10950 = n10221 ^ n10141;
  assign n10951 = n10251 & ~n10950;
  assign n10952 = n10951 ^ n10250;
  assign n10956 = n10955 ^ n10952;
  assign n9353 = x494 ^ x493;
  assign n10167 = x495 & x496;
  assign n10168 = x497 & x498;
  assign n10169 = ~n10167 & ~n10168;
  assign n10170 = ~x495 & ~x496;
  assign n10171 = ~x497 & ~x498;
  assign n10172 = ~n10170 & ~n10171;
  assign n10173 = n10169 & ~n10172;
  assign n10174 = ~n9353 & n10173;
  assign n10175 = n10167 & n10168;
  assign n10176 = n10170 & n10171;
  assign n10177 = ~n10175 & ~n10176;
  assign n10178 = ~n10174 & n10177;
  assign n10179 = x493 & x494;
  assign n10180 = ~n10178 & ~n10179;
  assign n10181 = ~n10175 & n10179;
  assign n10182 = n10181 ^ n10172;
  assign n10183 = n10181 ^ n9353;
  assign n10184 = n10172 ^ n10169;
  assign n10185 = n10184 ^ n10181;
  assign n10186 = ~n10181 & ~n10185;
  assign n10187 = n10186 ^ n10181;
  assign n10188 = n10183 & ~n10187;
  assign n10189 = n10188 ^ n10186;
  assign n10190 = n10189 ^ n10181;
  assign n10191 = n10190 ^ n10184;
  assign n10192 = n10182 & ~n10191;
  assign n10193 = n10192 ^ n10181;
  assign n10194 = ~n10180 & ~n10193;
  assign n9359 = x488 ^ x487;
  assign n10143 = x489 & x490;
  assign n10144 = ~x491 & ~x492;
  assign n10145 = ~n10143 & n10144;
  assign n10146 = ~x489 & ~x490;
  assign n10147 = x491 & x492;
  assign n10148 = n10146 & ~n10147;
  assign n10149 = ~n10145 & ~n10148;
  assign n10150 = ~n9359 & ~n10149;
  assign n10151 = n10143 & n10147;
  assign n10152 = n10144 & n10146;
  assign n10153 = ~n10151 & ~n10152;
  assign n10154 = ~n10150 & n10153;
  assign n10155 = x487 & x488;
  assign n10156 = ~n10154 & ~n10155;
  assign n9357 = x490 ^ x489;
  assign n9356 = x492 ^ x491;
  assign n9358 = n9357 ^ n9356;
  assign n10157 = n9358 ^ x488;
  assign n10158 = n10157 ^ n9358;
  assign n10159 = n10151 ^ n9358;
  assign n10160 = n10159 ^ n9358;
  assign n10161 = n10158 & ~n10160;
  assign n10162 = n10161 ^ n9358;
  assign n10163 = ~n9359 & n10162;
  assign n10164 = n10163 ^ n9358;
  assign n10165 = n10149 & n10164;
  assign n10166 = ~n10156 & ~n10165;
  assign n10195 = n10194 ^ n10166;
  assign n9360 = n9359 ^ n9358;
  assign n9352 = x496 ^ x495;
  assign n9354 = n9353 ^ n9352;
  assign n9351 = x498 ^ x497;
  assign n9355 = n9354 ^ n9351;
  assign n9361 = n9360 ^ n9355;
  assign n9350 = n9349 ^ n9344;
  assign n10138 = n9355 ^ n9350;
  assign n10139 = n9361 & ~n10138;
  assign n10140 = n10139 ^ n9360;
  assign n10142 = n10141 ^ n10140;
  assign n10196 = n10195 ^ n10142;
  assign n10959 = n10196 & ~n10251;
  assign n10945 = n9355 & n9360;
  assign n10960 = n10945 ^ n10140;
  assign n10961 = n10195 & ~n10960;
  assign n10962 = n10961 ^ n10140;
  assign n10963 = ~n10959 & n10962;
  assign n10964 = n10141 & n10251;
  assign n10965 = n10963 & ~n10964;
  assign n10958 = ~n10175 & ~n10193;
  assign n10966 = n10965 ^ n10958;
  assign n10946 = n10195 & n10945;
  assign n10947 = n10166 & n10194;
  assign n10948 = ~n10946 & ~n10947;
  assign n10944 = ~n10151 & ~n10165;
  assign n10949 = n10948 ^ n10944;
  assign n10957 = n10956 ^ n10949;
  assign n10967 = n10966 ^ n10957;
  assign n11307 = n10956 & n10967;
  assign n11308 = ~n10944 & ~n10948;
  assign n11309 = ~n11307 & ~n11308;
  assign n11310 = n10958 & ~n10965;
  assign n11311 = n11309 & n11310;
  assign n11312 = n10948 & ~n10956;
  assign n11313 = n10944 & n11312;
  assign n11314 = n11313 ^ n11307;
  assign n11315 = n11313 ^ n11308;
  assign n11316 = ~n10958 & n10965;
  assign n11317 = n11316 ^ n11313;
  assign n11318 = ~n11313 & n11317;
  assign n11319 = n11318 ^ n11313;
  assign n11320 = ~n11315 & ~n11319;
  assign n11321 = n11320 ^ n11318;
  assign n11322 = n11321 ^ n11313;
  assign n11323 = n11322 ^ n11316;
  assign n11324 = n11314 & n11323;
  assign n11325 = n11324 ^ n11307;
  assign n11326 = ~n11311 & ~n11325;
  assign n11304 = n10954 ^ n10952;
  assign n11305 = ~n10955 & ~n11304;
  assign n11306 = n11305 ^ n10952;
  assign n11327 = n11326 ^ n11306;
  assign n10327 = x479 & x480;
  assign n10328 = x477 & x478;
  assign n10329 = ~n10327 & ~n10328;
  assign n10330 = ~x479 & ~x480;
  assign n10331 = ~x477 & ~x478;
  assign n10332 = ~n10330 & ~n10331;
  assign n10333 = ~n10329 & n10332;
  assign n10334 = x476 & n10333;
  assign n10335 = n10327 & n10328;
  assign n10336 = ~n10334 & ~n10335;
  assign n10343 = n10333 ^ x476;
  assign n10344 = n10343 ^ n10333;
  assign n10337 = n10329 & ~n10332;
  assign n10345 = ~n10335 & ~n10337;
  assign n10346 = n10345 ^ n10333;
  assign n10347 = n10344 & n10346;
  assign n10348 = n10347 ^ n10333;
  assign n10349 = x475 & n10348;
  assign n10931 = n10336 & ~n10349;
  assign n10353 = x485 & x486;
  assign n10352 = x483 & x484;
  assign n10354 = n10353 ^ n10352;
  assign n10355 = ~x485 & ~x486;
  assign n10356 = ~x483 & ~x484;
  assign n10357 = ~n10355 & ~n10356;
  assign n10358 = n10357 ^ n10352;
  assign n10359 = n10358 ^ n10352;
  assign n10360 = n10352 ^ x482;
  assign n10361 = n10360 ^ n10352;
  assign n10362 = n10359 & n10361;
  assign n10363 = n10362 ^ n10352;
  assign n10364 = n10354 & ~n10363;
  assign n10365 = n10364 ^ n10353;
  assign n9324 = x482 ^ x481;
  assign n10367 = ~n10352 & ~n10353;
  assign n10378 = n10357 & ~n10367;
  assign n10379 = n9324 & n10378;
  assign n10380 = ~n10357 & n10367;
  assign n10381 = x481 & x482;
  assign n10382 = n10352 & n10381;
  assign n10383 = x486 & n10382;
  assign n10384 = n10383 ^ n10381;
  assign n10385 = ~n10380 & n10384;
  assign n10386 = ~n10379 & ~n10385;
  assign n10930 = ~n10365 & n10386;
  assign n10932 = n10931 ^ n10930;
  assign n10366 = n10356 ^ n10355;
  assign n10368 = n10367 ^ n10356;
  assign n10369 = n10368 ^ n10356;
  assign n10370 = n10356 ^ x482;
  assign n10371 = n10370 ^ n10356;
  assign n10372 = n10369 & ~n10371;
  assign n10373 = n10372 ^ n10356;
  assign n10374 = n10366 & ~n10373;
  assign n10375 = n10374 ^ n10355;
  assign n10376 = ~n10365 & ~n10375;
  assign n10377 = ~x481 & ~n10376;
  assign n9323 = x484 ^ x483;
  assign n10387 = n10381 ^ x484;
  assign n10388 = n10387 ^ n10381;
  assign n10389 = ~x482 & ~x486;
  assign n10390 = n10389 ^ n10381;
  assign n10391 = ~n10388 & n10390;
  assign n10392 = n10391 ^ n10381;
  assign n10393 = ~n9323 & n10392;
  assign n10394 = ~x485 & n10393;
  assign n10395 = n10386 & ~n10394;
  assign n10396 = ~n10377 & n10395;
  assign n10338 = ~x476 & n10337;
  assign n10339 = n10336 & ~n10338;
  assign n10340 = ~x475 & ~n10339;
  assign n9319 = x476 ^ x475;
  assign n10341 = n10330 & n10331;
  assign n10342 = n9319 & n10341;
  assign n10350 = ~n10342 & ~n10349;
  assign n10351 = ~n10340 & n10350;
  assign n10397 = n10396 ^ n10351;
  assign n9318 = x478 ^ x477;
  assign n9320 = n9319 ^ n9318;
  assign n9317 = x480 ^ x479;
  assign n9321 = n9320 ^ n9317;
  assign n9325 = n9324 ^ n9323;
  assign n9322 = x486 ^ x485;
  assign n9326 = n9325 ^ n9322;
  assign n10323 = n9321 & n9326;
  assign n10927 = n10351 ^ n10323;
  assign n10928 = n10397 & ~n10927;
  assign n10929 = n10928 ^ n10396;
  assign n10933 = n10932 ^ n10929;
  assign n10293 = x467 & x468;
  assign n10294 = x465 & x466;
  assign n10295 = ~n10293 & ~n10294;
  assign n10296 = ~x467 & ~x468;
  assign n10297 = ~x465 & ~x466;
  assign n10298 = ~n10296 & ~n10297;
  assign n10299 = ~n10295 & n10298;
  assign n10300 = x464 & n10299;
  assign n10301 = n10293 & n10294;
  assign n10302 = ~n10300 & ~n10301;
  assign n10309 = n10299 ^ x464;
  assign n10310 = n10309 ^ n10299;
  assign n10303 = n10295 & ~n10298;
  assign n10311 = ~n10301 & ~n10303;
  assign n10312 = n10311 ^ n10299;
  assign n10313 = n10310 & n10312;
  assign n10314 = n10313 ^ n10299;
  assign n10315 = x463 & n10314;
  assign n10924 = n10302 & ~n10315;
  assign n10253 = x471 & x472;
  assign n10258 = x473 & x474;
  assign n10263 = n10253 & n10258;
  assign n10254 = ~x473 & ~x474;
  assign n10264 = x470 & ~n10254;
  assign n10265 = ~n10263 & ~n10264;
  assign n9334 = x472 ^ x471;
  assign n10266 = n10258 ^ x472;
  assign n10267 = n9334 & ~n10266;
  assign n10268 = n10267 ^ x471;
  assign n10269 = ~n10265 & n10268;
  assign n10280 = ~n10254 & n10268;
  assign n10259 = ~x471 & ~x472;
  assign n10260 = ~n10258 & n10259;
  assign n10277 = x469 & ~n10260;
  assign n10255 = ~n10253 & n10254;
  assign n10278 = ~n10255 & ~n10263;
  assign n10279 = n10277 & n10278;
  assign n10281 = n10280 ^ n10279;
  assign n10282 = n10279 ^ x469;
  assign n10283 = n10279 ^ x470;
  assign n10284 = ~n10279 & n10283;
  assign n10285 = n10284 ^ n10279;
  assign n10286 = n10282 & ~n10285;
  assign n10287 = n10286 ^ n10284;
  assign n10288 = n10287 ^ n10279;
  assign n10289 = n10288 ^ x470;
  assign n10290 = n10281 & n10289;
  assign n10291 = n10290 ^ n10279;
  assign n10923 = ~n10269 & ~n10291;
  assign n10925 = n10924 ^ n10923;
  assign n10304 = ~x464 & n10303;
  assign n10305 = n10302 & ~n10304;
  assign n10306 = ~x463 & ~n10305;
  assign n9330 = x464 ^ x463;
  assign n10307 = n10296 & n10297;
  assign n10308 = n9330 & n10307;
  assign n10316 = ~n10308 & ~n10315;
  assign n10317 = ~n10306 & n10316;
  assign n10256 = ~x470 & n10255;
  assign n10257 = n10256 ^ x469;
  assign n10261 = n10260 ^ n10256;
  assign n10262 = n10261 ^ n10260;
  assign n10270 = n10260 & ~n10264;
  assign n10271 = ~n10269 & ~n10270;
  assign n10272 = n10271 ^ n10260;
  assign n10273 = ~n10262 & n10272;
  assign n10274 = n10273 ^ n10260;
  assign n10275 = ~n10257 & n10274;
  assign n10276 = n10275 ^ x469;
  assign n10292 = n10276 & ~n10291;
  assign n10318 = n10317 ^ n10292;
  assign n9329 = x468 ^ x467;
  assign n9331 = n9330 ^ n9329;
  assign n9328 = x466 ^ x465;
  assign n9332 = n9331 ^ n9328;
  assign n9335 = x474 ^ x473;
  assign n9336 = n9335 ^ n9334;
  assign n9333 = x470 ^ x469;
  assign n9337 = n9336 ^ n9333;
  assign n10319 = n9332 & n9337;
  assign n10920 = n10319 ^ n10317;
  assign n10921 = ~n10318 & n10920;
  assign n10922 = n10921 ^ n10319;
  assign n10926 = n10925 ^ n10922;
  assign n10934 = n10933 ^ n10926;
  assign n10935 = n10323 & n10397;
  assign n9327 = n9326 ^ n9321;
  assign n9338 = n9337 ^ n9332;
  assign n10320 = n9338 ^ n9326;
  assign n10321 = ~n9327 & n10320;
  assign n10322 = n10321 ^ n9338;
  assign n10936 = ~n10322 & ~n10397;
  assign n10324 = n10323 ^ n10322;
  assign n10325 = ~n10319 & ~n10324;
  assign n10326 = n10325 ^ n10323;
  assign n10398 = n10397 ^ n10326;
  assign n10399 = n10398 ^ n10318;
  assign n10937 = n10399 ^ n10398;
  assign n10938 = n10398 ^ n10319;
  assign n10939 = n10937 & ~n10938;
  assign n10940 = n10939 ^ n10398;
  assign n10941 = ~n10936 & n10940;
  assign n10942 = ~n10935 & n10941;
  assign n11279 = n10934 & n10942;
  assign n11280 = n10922 & n10933;
  assign n11281 = ~n11279 & ~n11280;
  assign n11282 = n10923 & n10924;
  assign n11283 = n11281 & n11282;
  assign n11284 = ~n10923 & ~n10924;
  assign n11285 = ~n10922 & ~n11284;
  assign n11286 = ~n11282 & ~n11285;
  assign n11287 = n10942 & n11286;
  assign n11288 = n10933 & n11287;
  assign n11289 = n11284 ^ n10922;
  assign n11290 = n11284 ^ n10942;
  assign n11291 = n10933 ^ n10922;
  assign n11292 = n11291 ^ n11284;
  assign n11293 = ~n11284 & n11292;
  assign n11294 = n11293 ^ n11284;
  assign n11295 = ~n11290 & ~n11294;
  assign n11296 = n11295 ^ n11293;
  assign n11297 = n11296 ^ n11284;
  assign n11298 = n11297 ^ n11291;
  assign n11299 = ~n11289 & n11298;
  assign n11300 = ~n11288 & ~n11299;
  assign n11301 = ~n11283 & n11300;
  assign n11276 = n10931 ^ n10929;
  assign n11277 = ~n10932 & ~n11276;
  assign n11278 = n11277 ^ n10929;
  assign n11302 = n11301 ^ n11278;
  assign n10943 = n10942 ^ n10934;
  assign n10968 = n10967 ^ n10943;
  assign n10252 = n10251 ^ n10196;
  assign n10400 = n10399 ^ n10252;
  assign n9339 = n9338 ^ n9327;
  assign n9362 = n9361 ^ n9350;
  assign n10916 = n9339 & n9362;
  assign n10917 = n10916 ^ n10252;
  assign n10918 = ~n10400 & ~n10917;
  assign n10919 = n10918 ^ n10399;
  assign n11273 = n10943 ^ n10919;
  assign n11274 = ~n10968 & n11273;
  assign n11275 = n11274 ^ n10967;
  assign n11303 = n11302 ^ n11275;
  assign n11328 = n11327 ^ n11303;
  assign n11030 = n11029 ^ n10980;
  assign n10970 = n10400 & n10644;
  assign n9363 = n9362 ^ n9339;
  assign n9410 = n9409 ^ n9386;
  assign n10971 = n9363 & n9410;
  assign n10972 = ~n10970 & n10971;
  assign n10973 = n10916 ^ n10400;
  assign n10975 = n10974 ^ n10644;
  assign n10976 = ~n10973 & ~n10975;
  assign n10977 = ~n10972 & ~n10976;
  assign n11031 = n11030 ^ n10977;
  assign n10969 = n10968 ^ n10919;
  assign n11270 = n10977 ^ n10969;
  assign n11271 = ~n11031 & n11270;
  assign n11272 = n11271 ^ n11030;
  assign n11329 = n11328 ^ n11272;
  assign n11384 = n11383 ^ n11353;
  assign n11580 = n11384 ^ n11272;
  assign n11581 = n11329 & ~n11580;
  assign n11582 = n11581 ^ n11384;
  assign n11591 = n11590 ^ n11582;
  assign n11598 = ~n10944 & ~n11327;
  assign n11599 = n11306 & ~n11312;
  assign n11600 = ~n11598 & ~n11599;
  assign n11601 = ~n11310 & ~n11600;
  assign n11602 = ~n11309 & ~n11327;
  assign n11603 = n11306 & n11316;
  assign n11604 = ~n11602 & ~n11603;
  assign n11605 = ~n11601 & n11604;
  assign n11595 = ~n11284 & n11302;
  assign n11596 = ~n11278 & n11281;
  assign n11597 = ~n11595 & ~n11596;
  assign n11606 = n11605 ^ n11597;
  assign n11592 = n11327 ^ n11302;
  assign n11593 = n11303 & n11592;
  assign n11594 = n11593 ^ n11327;
  assign n11607 = n11606 ^ n11594;
  assign n11752 = n11607 ^ n11590;
  assign n11753 = n11591 & ~n11752;
  assign n11754 = n11753 ^ n11607;
  assign n11755 = n11588 ^ n11585;
  assign n11756 = n11585 ^ n11375;
  assign n11757 = ~n11755 & n11756;
  assign n11758 = n11757 ^ n11375;
  assign n11759 = n11597 ^ n11594;
  assign n11760 = ~n11606 & ~n11759;
  assign n11761 = n11760 ^ n11605;
  assign n11828 = ~n11758 & n11761;
  assign n11829 = n11754 & n11828;
  assign n11608 = n11607 ^ n11591;
  assign n11268 = n11267 ^ n11218;
  assign n11032 = n11031 ^ n10969;
  assign n9411 = n9410 ^ n9363;
  assign n9509 = ~n9411 & ~n9508;
  assign n9510 = ~n9434 & ~n9457;
  assign n9511 = ~n9505 & n9510;
  assign n9512 = ~n9509 & ~n9511;
  assign n10133 = n9409 ^ n9339;
  assign n10135 = n10133 ^ n9386;
  assign n10136 = ~n9362 & n10135;
  assign n10134 = ~n9410 & ~n10133;
  assign n10137 = n10136 ^ n10134;
  assign n10401 = n10400 ^ n10137;
  assign n10645 = n10644 ^ n10401;
  assign n10900 = n9457 & n9505;
  assign n10901 = n10645 & ~n10900;
  assign n10902 = n9512 & ~n10901;
  assign n10903 = ~n10131 & ~n10902;
  assign n10904 = n9508 & n10131;
  assign n10905 = n10904 ^ n10645;
  assign n9514 = n9411 & n9505;
  assign n10906 = ~n9458 & n9514;
  assign n10907 = n10906 ^ n10904;
  assign n10908 = n10907 ^ n10906;
  assign n10649 = n9505 ^ n9458;
  assign n10909 = n9411 & n10649;
  assign n10910 = n10909 ^ n10906;
  assign n10911 = ~n10908 & ~n10910;
  assign n10912 = n10911 ^ n10906;
  assign n10913 = n10905 & ~n10912;
  assign n10914 = n10913 ^ n10645;
  assign n10915 = ~n10903 & ~n10914;
  assign n11033 = n11032 ^ n10915;
  assign n11102 = n11101 ^ n11038;
  assign n11164 = n11163 ^ n11102;
  assign n11169 = n11164 ^ n10915;
  assign n11170 = ~n11033 & n11169;
  assign n11171 = n11170 ^ n11032;
  assign n11269 = n11268 ^ n11171;
  assign n11385 = n11384 ^ n11329;
  assign n11577 = n11385 ^ n11171;
  assign n11578 = n11269 & ~n11577;
  assign n11579 = n11578 ^ n11385;
  assign n11609 = n11608 ^ n11579;
  assign n11749 = n11639 ^ n11608;
  assign n11750 = ~n11609 & ~n11749;
  assign n11751 = n11750 ^ n11639;
  assign n11762 = n11761 ^ n11758;
  assign n11822 = n11761 ^ n11754;
  assign n11823 = n11762 & n11822;
  assign n11824 = n11823 ^ n11754;
  assign n11834 = n11751 & n11824;
  assign n11835 = ~n11829 & ~n11834;
  assign n11836 = n11835 ^ n11777;
  assign n11837 = ~n11781 & n11836;
  assign n11815 = n11614 & n11618;
  assign n11816 = n11781 & ~n11815;
  assign n11817 = ~n11766 & ~n11775;
  assign n11818 = ~n11816 & ~n11817;
  assign n11819 = n11758 & ~n11761;
  assign n11820 = ~n11754 & n11819;
  assign n11821 = ~n11818 & n11820;
  assign n11825 = ~n11751 & ~n11824;
  assign n11826 = ~n11821 & ~n11825;
  assign n11844 = n11818 & ~n11829;
  assign n11845 = n11826 & ~n11844;
  assign n11846 = ~n11837 & ~n11845;
  assign n11859 = n11858 ^ n11846;
  assign n11797 = ~n11714 & ~n11745;
  assign n11710 = n11709 ^ n11706;
  assign n11798 = n11709 ^ n11703;
  assign n11799 = n11710 & n11798;
  assign n11800 = n11799 ^ n11703;
  assign n11801 = n11797 & n11800;
  assign n11804 = n11802 & n11803;
  assign n11805 = ~n11801 & ~n11804;
  assign n11807 = ~n11706 & n11806;
  assign n11808 = n11807 ^ n11800;
  assign n11809 = n11714 & ~n11808;
  assign n11810 = n11745 & n11809;
  assign n11811 = n11810 ^ n11807;
  assign n11812 = n11805 & ~n11811;
  assign n11813 = n11812 ^ n11796;
  assign n11711 = n11710 ^ n11703;
  assign n11747 = n11746 ^ n11711;
  assign n11640 = n11639 ^ n11609;
  assign n11386 = n11385 ^ n11269;
  assign n10898 = n10897 ^ n10893;
  assign n9515 = n9513 & n9514;
  assign n9516 = n9512 & ~n9515;
  assign n10132 = n10131 ^ n9516;
  assign n10646 = n10645 ^ n10132;
  assign n9316 = n9315 ^ n8002;
  assign n10647 = n10646 ^ n9316;
  assign n10648 = ~n7906 & ~n8001;
  assign n10650 = n10649 ^ n9411;
  assign n10651 = ~n10648 & n10650;
  assign n10652 = n10651 ^ n10646;
  assign n10653 = n10652 ^ n10646;
  assign n10654 = n10646 ^ n8002;
  assign n10655 = n10654 ^ n10646;
  assign n10656 = n10653 & ~n10655;
  assign n10657 = n10656 ^ n10646;
  assign n10658 = n10647 & ~n10657;
  assign n10659 = n10658 ^ n10646;
  assign n10899 = n10898 ^ n10659;
  assign n11165 = n11164 ^ n11033;
  assign n11166 = n11165 ^ n10659;
  assign n11167 = n10899 & n11166;
  assign n11168 = n11167 ^ n10898;
  assign n11387 = n11386 ^ n11168;
  assign n11573 = n11572 ^ n11479;
  assign n11574 = n11573 ^ n11168;
  assign n11575 = n11387 & ~n11574;
  assign n11576 = n11575 ^ n11386;
  assign n11641 = n11640 ^ n11576;
  assign n11697 = n11696 ^ n11644;
  assign n11698 = n11697 ^ n11640;
  assign n11699 = ~n11641 & ~n11698;
  assign n11700 = n11699 ^ n11697;
  assign n11748 = n11747 ^ n11700;
  assign n11763 = n11762 ^ n11754;
  assign n11764 = n11763 ^ n11751;
  assign n11782 = n11781 ^ n11764;
  assign n11783 = n11782 ^ n11700;
  assign n11784 = n11748 & n11783;
  assign n11785 = n11784 ^ n11747;
  assign n11814 = n11813 ^ n11785;
  assign n11827 = n11781 & n11826;
  assign n11830 = ~n11818 & ~n11829;
  assign n11831 = n11751 & ~n11820;
  assign n11832 = ~n11830 & n11831;
  assign n11833 = n11827 & ~n11832;
  assign n11838 = n11818 & n11829;
  assign n11839 = ~n11837 & ~n11838;
  assign n11840 = ~n11833 & n11839;
  assign n11841 = n11840 ^ n11785;
  assign n11842 = n11814 & n11841;
  assign n11843 = n11842 ^ n11813;
  assign n11860 = n11859 ^ n11843;
  assign n11862 = n11861 ^ n11860;
  assign n11905 = n7737 ^ n7698;
  assign n11864 = n7676 ^ n7545;
  assign n11863 = n11782 ^ n11748;
  assign n11865 = n11864 ^ n11863;
  assign n11896 = n7500 ^ n7331;
  assign n11866 = n7212 ^ n6881;
  assign n11867 = n11573 ^ n11387;
  assign n11868 = n11866 & ~n11867;
  assign n11870 = n6604 ^ n6092;
  assign n11869 = n11165 ^ n10899;
  assign n11871 = n11870 ^ n11869;
  assign n11876 = n3179 ^ n2988;
  assign n11877 = n3182 ^ n3179;
  assign n11878 = n11876 & ~n11877;
  assign n11879 = n11878 ^ n2988;
  assign n11880 = n11879 ^ n2797;
  assign n11881 = n11880 ^ n5758;
  assign n11872 = n10651 ^ n9314;
  assign n11873 = ~n8002 & ~n11872;
  assign n11874 = n11873 ^ n9313;
  assign n11875 = n11874 ^ n10646;
  assign n11882 = n11881 ^ n11875;
  assign n11883 = n11876 ^ n3182;
  assign n11884 = n8001 ^ n7906;
  assign n11885 = n11884 ^ n10650;
  assign n11886 = n11883 & n11885;
  assign n11887 = n11886 ^ n11875;
  assign n11888 = ~n11882 & n11887;
  assign n11889 = n11888 ^ n11881;
  assign n11890 = n11889 ^ n11869;
  assign n11891 = ~n11871 & ~n11890;
  assign n11892 = n11891 ^ n11870;
  assign n11893 = ~n11868 & n11892;
  assign n11894 = ~n11866 & n11867;
  assign n11895 = ~n11893 & ~n11894;
  assign n11897 = n11896 ^ n11895;
  assign n11898 = n11697 ^ n11641;
  assign n11899 = n11898 ^ n11895;
  assign n11900 = n11897 & ~n11899;
  assign n11901 = n11900 ^ n11896;
  assign n11902 = n11901 ^ n11863;
  assign n11903 = ~n11865 & n11902;
  assign n11904 = n11903 ^ n11864;
  assign n11906 = n11905 ^ n11904;
  assign n11907 = n11840 ^ n11814;
  assign n11908 = n11907 ^ n11905;
  assign n11909 = n11906 & n11908;
  assign n11910 = n11909 ^ n11904;
  assign n11911 = n11910 ^ n11860;
  assign n11912 = ~n11862 & ~n11911;
  assign n11913 = n11912 ^ n11861;
  assign n11914 = n11913 ^ n7794;
  assign n11915 = n7811 & n11914;
  assign n11916 = n11915 ^ n11913;
  assign n11920 = n7794 & ~n7810;
  assign n11921 = n11913 & n11920;
  assign n11917 = n11858 ^ n11843;
  assign n11918 = ~n11859 & n11917;
  assign n11919 = n11918 ^ n11843;
  assign n11922 = n11921 ^ n11919;
  assign n11923 = ~n11904 & ~n11905;
  assign n11924 = n11907 & n11923;
  assign n11925 = n11893 & ~n11894;
  assign n11926 = n11867 ^ n11866;
  assign n11927 = ~n11869 & n11870;
  assign n11928 = ~n11889 & n11927;
  assign n11929 = n11885 ^ n11883;
  assign n11930 = n11885 ^ n11882;
  assign n11931 = ~n11929 & n11930;
  assign n11932 = ~x1000 & n11931;
  assign n11933 = ~n11928 & ~n11932;
  assign n11934 = n11892 & ~n11933;
  assign n11935 = n11926 & ~n11934;
  assign n11936 = n11869 & ~n11870;
  assign n11937 = n11889 & ~n11932;
  assign n11938 = n11936 & n11937;
  assign n11939 = ~n11935 & ~n11938;
  assign n11940 = ~n11925 & n11939;
  assign n11941 = ~n11895 & ~n11896;
  assign n11942 = ~n11898 & n11941;
  assign n11943 = ~n11901 & ~n11942;
  assign n11944 = n11943 ^ n11865;
  assign n11945 = n11944 ^ n11943;
  assign n11946 = n11895 & n11896;
  assign n11947 = n11898 & n11946;
  assign n11948 = n11947 ^ n11943;
  assign n11949 = n11945 & n11948;
  assign n11950 = n11949 ^ n11943;
  assign n11951 = ~n11940 & n11950;
  assign n11952 = ~n11924 & n11951;
  assign n11953 = n11910 ^ n11862;
  assign n11954 = n11953 ^ n11910;
  assign n11955 = n11904 & n11905;
  assign n11956 = ~n11907 & n11955;
  assign n11957 = n11956 ^ n11910;
  assign n11958 = n11954 & ~n11957;
  assign n11959 = n11958 ^ n11910;
  assign n11960 = n11952 & ~n11959;
  assign n11961 = n11960 ^ n11919;
  assign n11962 = ~n11922 & n11961;
  assign n11963 = n11962 ^ n11919;
  assign n11964 = n11916 & ~n11963;
  assign y0 = ~n11964;
endmodule
