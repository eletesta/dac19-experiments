// Benchmark "top" written by ABC on Mon Nov 19 13:33:26 2018

module top ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10;
  wire n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
    n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
    n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
    n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
    n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
    n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
    n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
    n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
    n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
    n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
    n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
    n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
    n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
    n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
    n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
    n215, n216, n217, n218, n219, n220, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
    n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
    n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
    n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
    n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
    n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
    n300, n301, n302, n303, n304, n305, n306, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
    n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
    n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
    n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n361,
    n362, n363, n364, n365, n366, n368, n369, n370, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
    n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
    n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
    n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
    n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
    n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
    n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
    n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n508, n509,
    n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n545, n546,
    n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n570, n571,
    n572, n573;
  assign n23 = ~pi0 & pi7;
  assign n24 = ~pi2 & ~pi8;
  assign n25 = pi2 & pi8;
  assign n26 = pi8 & ~pi9;
  assign n27 = n25 & ~pi9;
  assign n28 = ~n27 & ~n24;
  assign n29 = ~n28 & n23;
  assign n30 = pi0 & pi9;
  assign n31 = ~pi2 & pi8;
  assign n32 = pi8 & pi9;
  assign n33 = pi0 & ~pi2;
  assign n34 = n30 & n31;
  assign n35 = ~n29 & ~n34;
  assign n36 = ~n35 & ~pi3;
  assign n37 = ~pi3 & pi9;
  assign n38 = pi2 & ~pi3;
  assign n39 = n32 & n38;
  assign n40 = pi3 & ~pi9;
  assign n41 = ~pi8 & ~pi9;
  assign n42 = ~pi2 & pi3;
  assign n43 = n41 & n42;
  assign n44 = ~n39 & ~n43;
  assign n45 = ~n44 & ~pi0;
  assign n46 = ~n40 & pi2;
  assign n47 = ~n42 & pi0;
  assign n48 = n47 & ~n41;
  assign n49 = n48 & ~n46;
  assign n50 = pi2 & pi3;
  assign n51 = ~pi2 & ~pi3;
  assign n52 = ~n45 & ~n49;
  assign n53 = ~n52 & ~pi7;
  assign n54 = ~n36 & ~n53;
  assign n55 = ~n54 & ~pi1;
  assign n56 = ~pi7 & ~pi8;
  assign n57 = ~pi8 & pi9;
  assign n58 = ~pi7 & ~pi9;
  assign n59 = n51 & ~n58;
  assign n60 = ~n57 ^ pi0;
  assign n61 = n59 & ~n60;
  assign n62 = ~n61 & ~n56;
  assign n63 = ~pi5 & ~pi6;
  assign n64 = ~n55 ^ ~n62;
  assign n65 = ~n64 & n63;
  assign n66 = ~pi5 & pi8;
  assign n67 = pi0 & pi1;
  assign n68 = n67 & pi8;
  assign n69 = ~pi1 & ~pi2;
  assign n70 = n69 & ~pi5;
  assign n71 = pi5 & ~pi8;
  assign n72 = ~n51 & ~n71;
  assign n73 = ~n70 & n72;
  assign n74 = ~n73 & ~n68;
  assign n75 = ~n74 & ~n66;
  assign n76 = ~n42 & ~pi5;
  assign n77 = ~pi0 & ~pi1;
  assign n78 = ~n71 & n77;
  assign n79 = ~n76 & n78;
  assign n80 = n32 & ~n38;
  assign n81 = pi5 & pi9;
  assign n82 = ~n30 & ~n81;
  assign n83 = ~n80 & n82;
  assign n84 = ~n79 & ~n83;
  assign n85 = ~n75 & n84;
  assign n86 = ~n25 & ~pi3;
  assign n87 = ~pi1 & pi2;
  assign n88 = ~n87 & ~pi8;
  assign n89 = ~n86 & ~n88;
  assign n90 = ~pi1 & pi8;
  assign n91 = ~n90 & ~pi0;
  assign n92 = ~n89 & n91;
  assign n93 = ~n87 & pi8;
  assign n94 = ~pi1 & ~pi8;
  assign n95 = ~n94 & ~pi3;
  assign n96 = ~n93 & pi0;
  assign n97 = n96 & ~n95;
  assign n98 = ~pi5 & ~pi9;
  assign n99 = ~n92 & n98;
  assign n100 = n99 & ~n97;
  assign n101 = ~pi0 & ~pi2;
  assign n102 = n77 & ~pi2;
  assign n103 = n51 & n77;
  assign n104 = n41 & pi5;
  assign n105 = ~n103 & n104;
  assign n106 = pi6 & ~pi7;
  assign n107 = ~n105 & n106;
  assign n108 = ~n85 & n107;
  assign n109 = n108 & ~n100;
  assign n110 = pi0 & ~pi1;
  assign n111 = ~pi1 & pi9;
  assign n112 = ~n111 ^ ~pi2;
  assign n113 = n112 & n110;
  assign n114 = ~n113 & n86;
  assign n115 = n33 & ~pi9;
  assign n116 = n57 & pi2;
  assign n117 = ~n115 & ~n116;
  assign n118 = ~n117 & pi1;
  assign n119 = ~n31 & pi3;
  assign n120 = ~n118 & n119;
  assign n121 = ~n120 & ~n114;
  assign n122 = ~pi0 & ~pi9;
  assign n123 = ~pi0 ^ pi9;
  assign n124 = n123 & pi1;
  assign n125 = ~n124 & pi8;
  assign n126 = pi5 & ~pi6;
  assign n127 = n126 & ~pi7;
  assign n128 = ~n125 & n127;
  assign n129 = ~n121 & n128;
  assign n130 = ~n109 & ~n129;
  assign n131 = ~n65 & n130;
  assign n132 = ~n103 & pi4;
  assign n133 = ~pi3 & ~pi4;
  assign n134 = ~n41 & ~pi4;
  assign n135 = n103 & n134;
  assign n136 = ~pi5 & pi6;
  assign n137 = ~pi5 ^ ~pi6;
  assign n138 = n41 & pi4;
  assign n139 = n138 & ~n137;
  assign n140 = ~n132 & ~n139;
  assign n141 = n140 & ~n135;
  assign po00 = ~n131 & n141;
  assign n143 = n24 & n77;
  assign n144 = n25 & n110;
  assign n145 = ~n143 & n58;
  assign n146 = n145 & ~n144;
  assign n147 = ~pi3 & ~pi9;
  assign n148 = ~pi0 & pi8;
  assign n149 = pi1 & ~pi2;
  assign n150 = n148 & n149;
  assign n151 = ~pi7 & pi8;
  assign n152 = ~n24 & ~n151;
  assign n153 = ~n152 & n110;
  assign n154 = ~n153 & ~n150;
  assign n155 = ~n154 & n147;
  assign n156 = ~n69 & ~pi3;
  assign n157 = ~n33 & ~n77;
  assign n158 = n32 & pi7;
  assign n159 = ~n32 ^ ~pi7;
  assign n160 = n156 & n159;
  assign n161 = n160 & ~n157;
  assign n162 = ~n155 & ~n161;
  assign n163 = ~n162 ^ n146;
  assign n164 = n163 & n63;
  assign n165 = ~pi3 ^ ~pi9;
  assign n166 = ~n165 & pi1;
  assign n167 = ~n40 & pi1;
  assign n168 = ~n66 & ~pi9;
  assign n169 = n166 & ~n168;
  assign n170 = ~pi8 ^ ~pi9;
  assign n171 = ~pi1 & ~pi5;
  assign n172 = n165 & pi8;
  assign n173 = ~n41 & pi0;
  assign n174 = ~n173 & ~pi3;
  assign n175 = ~n174 & ~n172;
  assign n176 = ~n175 & n171;
  assign n177 = n51 & n67;
  assign n178 = ~n98 & ~pi2;
  assign n179 = ~n177 & ~n178;
  assign n180 = ~n148 & pi1;
  assign n181 = n180 & n81;
  assign n182 = ~n179 & ~n181;
  assign n183 = n57 & n110;
  assign n184 = ~n77 & ~pi3;
  assign n185 = pi0 & ~pi8;
  assign n186 = pi1 & pi9;
  assign n187 = n57 & n67;
  assign n188 = n184 & ~n187;
  assign n189 = ~n81 & pi2;
  assign n190 = ~n169 & n189;
  assign n191 = ~n176 & n190;
  assign n192 = ~n81 & pi3;
  assign n193 = ~n183 & n192;
  assign n194 = ~n188 & ~n193;
  assign n195 = n182 & ~n194;
  assign n196 = ~n195 & n106;
  assign n197 = ~n191 & n196;
  assign n198 = n144 & ~pi3;
  assign n199 = n50 & n57;
  assign n200 = ~n199 & ~n147;
  assign n201 = ~n200 & pi1;
  assign n202 = ~n201 & ~n198;
  assign n203 = ~n32 & ~n111;
  assign n204 = ~n51 & pi9;
  assign n205 = n203 & ~n204;
  assign n206 = n205 & ~pi0;
  assign n207 = ~n31 & pi1;
  assign n208 = ~n38 & ~pi9;
  assign n209 = ~n207 & n208;
  assign n210 = ~n206 & ~n209;
  assign n211 = n202 & n210;
  assign n212 = ~n211 & n127;
  assign n213 = ~n197 & ~n212;
  assign n214 = ~n164 & n213;
  assign n215 = ~pi0 & ~pi6;
  assign n216 = ~n215 & ~pi9;
  assign n217 = n69 & ~pi3;
  assign n218 = ~n216 & n217;
  assign n219 = ~n218 & pi4;
  assign n220 = ~n219 & ~n135;
  assign po01 = ~n214 & n220;
  assign n222 = ~pi6 & pi9;
  assign n223 = ~n136 & ~n222;
  assign n224 = ~n223 & n90;
  assign n225 = ~n27 & n66;
  assign n226 = ~n225 & ~n148;
  assign n227 = n226 & ~n224;
  assign n228 = pi2 & ~pi5;
  assign n229 = ~pi2 & ~pi6;
  assign n230 = ~n228 & ~n229;
  assign n231 = n230 & ~pi1;
  assign n232 = pi1 & ~pi9;
  assign n233 = n228 & n232;
  assign n234 = pi5 & pi6;
  assign n235 = ~n234 & ~pi0;
  assign n236 = ~n178 & n235;
  assign n237 = n236 & ~n233;
  assign n238 = n237 & ~n231;
  assign n239 = ~n227 & ~n238;
  assign n240 = pi1 & pi6;
  assign n241 = n240 & ~pi0;
  assign n242 = ~pi0 & pi2;
  assign n243 = n241 & n228;
  assign n244 = n30 & ~n240;
  assign n245 = ~n243 & ~n244;
  assign n246 = n232 & pi5;
  assign n247 = ~n230 & ~n246;
  assign n248 = ~n247 & pi0;
  assign n249 = ~n230 & n122;
  assign n250 = ~n249 & ~pi8;
  assign n251 = ~n248 & n250;
  assign n252 = n251 & n245;
  assign n253 = ~n239 & ~n252;
  assign n254 = pi3 & ~pi4;
  assign n255 = ~n253 & n254;
  assign n256 = n136 & ~pi8;
  assign n257 = n102 & ~n256;
  assign n258 = ~n257 ^ pi4;
  assign n259 = n258 & ~pi3;
  assign n260 = ~n255 & ~n259;
  assign n261 = ~pi6 & pi8;
  assign n262 = ~n31 & ~n229;
  assign n263 = n262 & ~n261;
  assign n264 = ~n263 & n186;
  assign n265 = ~n264 & ~pi0;
  assign n266 = ~n24 & pi0;
  assign n267 = ~n266 & n37;
  assign n268 = pi1 & ~pi6;
  assign n269 = ~n26 & n268;
  assign n270 = pi2 & ~pi6;
  assign n271 = ~n270 & ~pi3;
  assign n272 = ~n269 & n271;
  assign n273 = ~n267 & ~n272;
  assign n274 = ~n265 & ~n273;
  assign n275 = ~n274 & ~pi7;
  assign n276 = n173 & n149;
  assign n277 = ~n261 & ~pi1;
  assign n278 = n115 & n277;
  assign n279 = n32 & ~pi0;
  assign n280 = n32 & n242;
  assign n281 = ~n278 & ~n280;
  assign n282 = n281 & ~n276;
  assign n283 = ~n215 & ~pi8;
  assign n284 = ~n283 & ~n229;
  assign n285 = ~n270 & pi0;
  assign n286 = ~n285 & n232;
  assign n287 = ~n284 & n286;
  assign n288 = ~n25 & ~pi9;
  assign n289 = ~n32 & ~pi6;
  assign n290 = ~n289 & n77;
  assign n291 = n290 & ~n288;
  assign n292 = ~n287 & ~n291;
  assign n293 = n282 & n292;
  assign n294 = ~pi5 & ~pi7;
  assign n295 = n232 & pi0;
  assign n296 = ~n57 & n63;
  assign n297 = ~n295 & n296;
  assign n298 = ~n297 & ~n294;
  assign n299 = ~n23 & ~pi3;
  assign n300 = ~n299 & ~n147;
  assign n301 = n58 & ~pi0;
  assign n302 = n301 & n268;
  assign n303 = ~n300 & ~n302;
  assign n304 = ~n298 & n303;
  assign n305 = ~n293 & n304;
  assign n306 = ~n275 ^ ~n305;
  assign po02 = ~n260 & n306;
  assign n308 = pi0 & pi5;
  assign n309 = ~n170 & ~pi2;
  assign n310 = ~n41 & pi2;
  assign n311 = ~n309 & pi1;
  assign n312 = n311 & ~n310;
  assign n313 = ~pi1 & ~pi6;
  assign n314 = n69 & ~pi6;
  assign n315 = n314 & n41;
  assign n316 = ~n315 & ~n240;
  assign n317 = ~n312 & n316;
  assign n318 = ~n317 & n308;
  assign n319 = ~n148 & ~pi9;
  assign n320 = ~n111 & ~n148;
  assign n321 = ~n232 & pi6;
  assign n322 = ~n320 & n321;
  assign n323 = ~n322 & ~pi5;
  assign n324 = n32 & n77;
  assign n325 = ~n324 & ~pi6;
  assign n326 = ~n325 & ~n270;
  assign n327 = n323 & n326;
  assign n328 = n25 & n186;
  assign n329 = ~n328 & ~pi6;
  assign n330 = ~pi0 & pi5;
  assign n331 = ~n240 & n330;
  assign n332 = n136 & pi2;
  assign n333 = ~n331 & ~n332;
  assign n334 = ~n329 & ~n333;
  assign n335 = n233 & ~n148;
  assign n336 = ~n335 & ~pi3;
  assign n337 = ~n334 & n336;
  assign n338 = ~n327 & n337;
  assign n339 = ~n318 & n338;
  assign n340 = ~n261 & n330;
  assign n341 = ~n26 & ~pi5;
  assign n342 = ~n222 & pi0;
  assign n343 = n341 & n342;
  assign n344 = ~n343 & ~n340;
  assign n345 = ~n344 & pi1;
  assign n346 = ~n308 & pi1;
  assign n347 = n32 & ~pi6;
  assign n348 = ~n346 & n347;
  assign n349 = n110 & ~n126;
  assign n350 = ~n341 & n349;
  assign n351 = ~n348 & ~n350;
  assign n352 = ~n345 & n351;
  assign n353 = ~n112 & ~n234;
  assign n354 = ~n353 & pi3;
  assign n355 = ~n352 & n354;
  assign n356 = n217 & ~n137;
  assign n357 = ~n356 ^ ~pi4;
  assign n358 = ~n357 & ~pi7;
  assign n359 = ~n339 & n358;
  assign po03 = n359 & ~n355;
  assign n361 = n234 & ~pi7;
  assign n362 = ~n217 ^ ~pi4;
  assign n363 = ~n362 & n102;
  assign n364 = pi2 & ~pi4;
  assign n365 = ~n77 & n364;
  assign n366 = ~n363 & ~n365;
  assign po04 = ~n366 & n361;
  assign n368 = ~n102 & n254;
  assign n369 = n103 & pi4;
  assign n370 = ~n368 & ~n369;
  assign po05 = ~n370 & n361;
  assign n372 = n294 & ~pi2;
  assign n373 = n372 & ~n41;
  assign n374 = ~n373 & pi6;
  assign n375 = ~n328 & ~pi7;
  assign n376 = ~n375 & pi5;
  assign n377 = n372 & n222;
  assign n378 = ~n376 & ~n377;
  assign n379 = ~n374 & pi0;
  assign n380 = n378 & n379;
  assign n381 = ~n41 & ~pi7;
  assign n382 = ~n381 & pi2;
  assign n383 = n58 & n66;
  assign n384 = pi7 & ~pi8;
  assign n385 = ~n58 & ~pi2;
  assign n386 = ~n384 & pi1;
  assign n387 = ~n383 & n386;
  assign n388 = ~n382 & n387;
  assign n389 = ~n104 & ~n385;
  assign n390 = ~n158 & ~pi1;
  assign n391 = n389 & n390;
  assign n392 = ~n388 & ~n391;
  assign n393 = n380 & ~n392;
  assign n394 = ~n268 & pi5;
  assign n395 = ~n394 & ~n186;
  assign n396 = ~n395 & ~pi7;
  assign n397 = n98 & ~n240;
  assign n398 = ~n397 & n151;
  assign n399 = ~n32 & ~pi5;
  assign n400 = ~n151 & n313;
  assign n401 = ~n32 & n63;
  assign n402 = n399 & n400;
  assign n403 = ~n398 & pi2;
  assign n404 = ~n396 & ~n402;
  assign n405 = n404 & n403;
  assign n406 = n63 & ~pi1;
  assign n407 = n406 & ~n384;
  assign n408 = ~n56 & ~n63;
  assign n409 = ~n408 & ~pi9;
  assign n410 = ~n407 & n409;
  assign n411 = n56 & n240;
  assign n412 = ~n361 & ~pi2;
  assign n413 = n412 & ~n411;
  assign n414 = ~n410 & n413;
  assign n415 = ~n405 & ~n414;
  assign n416 = ~n393 ^ n415;
  assign n417 = ~n416 & n133;
  assign n418 = ~n67 & n71;
  assign n419 = n418 & ~n149;
  assign n420 = n419 & ~n115;
  assign n421 = n111 & n242;
  assign n422 = pi5 & pi8;
  assign n423 = ~n232 & n422;
  assign n424 = ~n421 & n423;
  assign n425 = ~n424 & ~pi4;
  assign n426 = ~n420 & n425;
  assign n427 = ~n426 & ~n234;
  assign n428 = ~pi2 & pi6;
  assign n429 = ~n148 & n428;
  assign n430 = ~n122 & ~n428;
  assign n431 = ~n429 & ~n430;
  assign n432 = ~n25 & ~n222;
  assign n433 = ~n432 & pi0;
  assign n434 = ~n57 & ~pi1;
  assign n435 = ~n431 & n434;
  assign n436 = n435 & ~n433;
  assign n437 = ~n263 & n279;
  assign n438 = ~n148 & ~pi2;
  assign n439 = n216 & n438;
  assign n440 = ~n439 & pi1;
  assign n441 = ~n437 & n440;
  assign n442 = ~n436 & ~n441;
  assign n443 = n442 & ~pi5;
  assign n444 = ~n443 & ~n427;
  assign n445 = ~n444 & ~n369;
  assign n446 = ~n133 & ~pi7;
  assign n447 = ~n445 & n446;
  assign po06 = ~n447 & ~n417;
  assign n449 = n124 & pi8;
  assign n450 = ~n449 & ~pi3;
  assign n451 = ~n95 & ~n90;
  assign n452 = n451 & ~n203;
  assign n453 = ~n279 & ~n77;
  assign n454 = ~n450 & n453;
  assign n455 = n454 & ~n452;
  assign n456 = ~n455 & ~pi2;
  assign n457 = n25 & n165;
  assign n458 = ~n37 & n185;
  assign n459 = n458 & ~n42;
  assign n460 = ~n459 & ~n457;
  assign n461 = ~n460 & pi1;
  assign n462 = ~n101 & ~pi3;
  assign n463 = n170 & n313;
  assign n464 = n462 & n463;
  assign n465 = ~n464 & n126;
  assign n466 = ~n461 & n465;
  assign n467 = ~n456 & n466;
  assign n468 = ~pi0 & pi3;
  assign n469 = ~n170 & n468;
  assign n470 = ~n310 & ~n469;
  assign n471 = ~n470 & ~pi1;
  assign n472 = n184 & n41;
  assign n473 = ~n41 & ~pi1;
  assign n474 = n203 & ~n90;
  assign n475 = ~n472 & n474;
  assign n476 = n173 & ~n111;
  assign n477 = ~n475 & ~n476;
  assign n478 = ~n477 & ~pi2;
  assign n479 = ~n471 & ~n39;
  assign n480 = ~n478 & n479;
  assign n481 = ~n480 & ~pi4;
  assign n482 = ~n37 & ~n242;
  assign n483 = n167 & ~n482;
  assign n484 = ~n111 & pi3;
  assign n485 = ~n484 & n33;
  assign n486 = ~n483 & ~n485;
  assign n487 = ~n486 & pi8;
  assign n488 = n38 & n186;
  assign n489 = ~n86 & ~n122;
  assign n490 = ~n24 & pi3;
  assign n491 = ~n490 & ~pi1;
  assign n492 = ~n489 & n491;
  assign n493 = ~n492 & ~n488;
  assign n494 = ~n487 & n493;
  assign n495 = ~n494 & ~pi4;
  assign n496 = ~n495 & ~pi6;
  assign n497 = ~n481 ^ n496;
  assign n498 = ~n497 & ~pi5;
  assign n499 = ~n498 & ~n467;
  assign n500 = ~n464 & pi7;
  assign n501 = n31 & n58;
  assign n502 = ~n501 & ~n384;
  assign n503 = n313 & pi0;
  assign n504 = ~n502 & n503;
  assign n505 = ~n500 & ~n504;
  assign n506 = n505 & ~n132;
  assign po07 = n499 | ~n506;
  assign n508 = n369 & n294;
  assign n509 = ~n246 & ~n30;
  assign n510 = ~n26 & n110;
  assign n511 = n320 & ~n510;
  assign n512 = n509 & n511;
  assign n513 = ~n512 & ~pi2;
  assign n514 = ~n288 & ~pi1;
  assign n515 = n514 & ~n399;
  assign n516 = ~n289 & ~n63;
  assign n517 = n336 & ~n515;
  assign n518 = ~n513 & n517;
  assign n519 = n518 & ~n516;
  assign n520 = n474 & ~n77;
  assign n521 = n42 & n126;
  assign n522 = ~n324 & n521;
  assign n523 = ~n520 & n522;
  assign n524 = ~pi2 ^ ~pi6;
  assign n525 = n524 & pi9;
  assign n526 = ~n180 & n525;
  assign n527 = ~n102 & ~n313;
  assign n528 = ~n283 & ~pi9;
  assign n529 = ~n527 & n528;
  assign n530 = ~n90 & n229;
  assign n531 = pi3 & ~pi5;
  assign n532 = ~n530 & n531;
  assign n533 = ~n526 & n532;
  assign n534 = ~n529 & n533;
  assign n535 = ~n523 & ~n534;
  assign n536 = ~n519 & n535;
  assign n537 = ~n232 & ~pi2;
  assign n538 = n310 & n77;
  assign n539 = ~n538 & ~n537;
  assign n540 = ~n539 & n401;
  assign n541 = ~n540 & pi7;
  assign n542 = ~n541 & ~pi4;
  assign n543 = ~n536 & n542;
  assign po08 = ~n543 & ~n508;
  assign n545 = ~n323 & ~n325;
  assign n546 = n453 & ~n473;
  assign n547 = n546 & n63;
  assign n548 = ~n545 & ~n547;
  assign n549 = ~n63 & ~pi2;
  assign n550 = ~n137 & pi2;
  assign n551 = ~n549 & ~n550;
  assign n552 = ~n548 & ~n551;
  assign n553 = pi3 & ~pi7;
  assign n554 = ~n552 & n553;
  assign n555 = n474 & n270;
  assign n556 = ~n63 & ~n69;
  assign n557 = ~n555 & n556;
  assign n558 = n110 & ~pi2;
  assign n559 = ~n319 & n149;
  assign n560 = ~n558 & ~pi7;
  assign n561 = ~n559 & n560;
  assign n562 = ~n561 & ~n538;
  assign n563 = n25 & n111;
  assign n564 = ~n563 & ~pi3;
  assign n565 = ~n356 & n564;
  assign n566 = ~n562 & n565;
  assign n567 = n566 & ~n557;
  assign n568 = ~n554 & ~n567;
  assign po09 = ~n568 & ~n362;
  assign n570 = n546 & n50;
  assign n571 = ~n570 & ~pi4;
  assign n572 = n63 & ~pi7;
  assign n573 = ~n132 & n572;
  assign po10 = ~n571 & n573;
endmodule


