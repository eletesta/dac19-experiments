module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128;
  wire n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103;
  assign n257 = x128 ^ x0;
  assign n259 = x0 & x128;
  assign n258 = x129 ^ x1;
  assign n260 = n259 ^ n258;
  assign n264 = x130 ^ x2;
  assign n261 = n259 ^ x129;
  assign n262 = n258 & ~n261;
  assign n263 = n262 ^ x1;
  assign n265 = n264 ^ n263;
  assign n269 = x131 ^ x3;
  assign n266 = n263 ^ x130;
  assign n267 = n264 & ~n266;
  assign n268 = n267 ^ x2;
  assign n270 = n269 ^ n268;
  assign n274 = x132 ^ x4;
  assign n271 = n268 ^ x131;
  assign n272 = n269 & ~n271;
  assign n273 = n272 ^ x3;
  assign n275 = n274 ^ n273;
  assign n277 = n269 & n274;
  assign n278 = n268 & n277;
  assign n279 = x3 & x131;
  assign n280 = n279 ^ x132;
  assign n281 = n274 & ~n280;
  assign n282 = n281 ^ x4;
  assign n283 = ~n278 & ~n282;
  assign n276 = x133 ^ x5;
  assign n284 = n283 ^ n276;
  assign n288 = x134 ^ x6;
  assign n285 = n283 ^ x133;
  assign n286 = n276 & n285;
  assign n287 = n286 ^ x5;
  assign n289 = n288 ^ n287;
  assign n291 = n276 & n288;
  assign n292 = ~n283 & n291;
  assign n293 = x5 & x133;
  assign n294 = n293 ^ x134;
  assign n295 = n288 & ~n294;
  assign n296 = n295 ^ x6;
  assign n297 = ~n292 & ~n296;
  assign n290 = x135 ^ x7;
  assign n298 = n297 ^ n290;
  assign n302 = x136 ^ x8;
  assign n299 = n297 ^ x135;
  assign n300 = n290 & n299;
  assign n301 = n300 ^ x7;
  assign n303 = n302 ^ n301;
  assign n305 = n290 & n302;
  assign n306 = ~n297 & n305;
  assign n307 = x7 & x135;
  assign n308 = n307 ^ x136;
  assign n309 = n302 & ~n308;
  assign n310 = n309 ^ x8;
  assign n311 = ~n306 & ~n310;
  assign n304 = x137 ^ x9;
  assign n312 = n311 ^ n304;
  assign n314 = x9 & x137;
  assign n315 = n304 & ~n311;
  assign n316 = ~n314 & ~n315;
  assign n313 = x138 ^ x10;
  assign n317 = n316 ^ n313;
  assign n326 = x139 ^ x11;
  assign n318 = n315 ^ x138;
  assign n319 = n318 ^ x138;
  assign n320 = n314 ^ x138;
  assign n321 = n320 ^ x138;
  assign n322 = ~n319 & ~n321;
  assign n323 = n322 ^ x138;
  assign n324 = n313 & n323;
  assign n325 = n324 ^ x10;
  assign n327 = n326 ^ n325;
  assign n331 = x140 ^ x12;
  assign n328 = n325 ^ x139;
  assign n329 = n326 & ~n328;
  assign n330 = n329 ^ x11;
  assign n332 = n331 ^ n330;
  assign n334 = n326 & n331;
  assign n335 = n325 & n334;
  assign n336 = x11 & x139;
  assign n337 = n336 ^ x140;
  assign n338 = n331 & ~n337;
  assign n339 = n338 ^ x12;
  assign n340 = ~n335 & ~n339;
  assign n333 = x141 ^ x13;
  assign n341 = n340 ^ n333;
  assign n345 = x142 ^ x14;
  assign n342 = n340 ^ x141;
  assign n343 = n333 & n342;
  assign n344 = n343 ^ x13;
  assign n346 = n345 ^ n344;
  assign n348 = n333 & n345;
  assign n349 = ~n340 & n348;
  assign n350 = x13 & x141;
  assign n351 = n350 ^ x142;
  assign n352 = n345 & ~n351;
  assign n353 = n352 ^ x14;
  assign n354 = ~n349 & ~n353;
  assign n347 = x143 ^ x15;
  assign n355 = n354 ^ n347;
  assign n359 = x144 ^ x16;
  assign n356 = n354 ^ x143;
  assign n357 = n347 & n356;
  assign n358 = n357 ^ x15;
  assign n360 = n359 ^ n358;
  assign n362 = n347 & n359;
  assign n363 = ~n354 & n362;
  assign n364 = x15 & x143;
  assign n365 = n364 ^ x144;
  assign n366 = n359 & ~n365;
  assign n367 = n366 ^ x16;
  assign n368 = ~n363 & ~n367;
  assign n361 = x145 ^ x17;
  assign n369 = n368 ^ n361;
  assign n373 = x146 ^ x18;
  assign n370 = n368 ^ x145;
  assign n371 = n361 & n370;
  assign n372 = n371 ^ x17;
  assign n374 = n373 ^ n372;
  assign n376 = n361 & n373;
  assign n377 = ~n368 & n376;
  assign n378 = x17 & x145;
  assign n379 = n378 ^ x146;
  assign n380 = n373 & ~n379;
  assign n381 = n380 ^ x18;
  assign n382 = ~n377 & ~n381;
  assign n375 = x147 ^ x19;
  assign n383 = n382 ^ n375;
  assign n385 = x19 & x147;
  assign n386 = n375 & ~n382;
  assign n387 = ~n385 & ~n386;
  assign n384 = x148 ^ x20;
  assign n388 = n387 ^ n384;
  assign n397 = x149 ^ x21;
  assign n389 = n386 ^ x148;
  assign n390 = n389 ^ x148;
  assign n391 = n385 ^ x148;
  assign n392 = n391 ^ x148;
  assign n393 = ~n390 & ~n392;
  assign n394 = n393 ^ x148;
  assign n395 = n384 & n394;
  assign n396 = n395 ^ x20;
  assign n398 = n397 ^ n396;
  assign n402 = x150 ^ x22;
  assign n399 = n396 ^ x149;
  assign n400 = n397 & ~n399;
  assign n401 = n400 ^ x21;
  assign n403 = n402 ^ n401;
  assign n405 = n397 & n402;
  assign n406 = n396 & n405;
  assign n407 = x21 & x149;
  assign n408 = n407 ^ x150;
  assign n409 = n402 & ~n408;
  assign n410 = n409 ^ x22;
  assign n411 = ~n406 & ~n410;
  assign n404 = x151 ^ x23;
  assign n412 = n411 ^ n404;
  assign n416 = x152 ^ x24;
  assign n413 = n411 ^ x151;
  assign n414 = n404 & n413;
  assign n415 = n414 ^ x23;
  assign n417 = n416 ^ n415;
  assign n419 = n404 & n416;
  assign n420 = ~n411 & n419;
  assign n421 = x23 & x151;
  assign n422 = n421 ^ x152;
  assign n423 = n416 & ~n422;
  assign n424 = n423 ^ x24;
  assign n425 = ~n420 & ~n424;
  assign n418 = x153 ^ x25;
  assign n426 = n425 ^ n418;
  assign n430 = x154 ^ x26;
  assign n427 = n425 ^ x153;
  assign n428 = n418 & n427;
  assign n429 = n428 ^ x25;
  assign n431 = n430 ^ n429;
  assign n433 = n418 & n430;
  assign n434 = ~n425 & n433;
  assign n435 = x25 & x153;
  assign n436 = n435 ^ x154;
  assign n437 = n430 & ~n436;
  assign n438 = n437 ^ x26;
  assign n439 = ~n434 & ~n438;
  assign n432 = x155 ^ x27;
  assign n440 = n439 ^ n432;
  assign n444 = x156 ^ x28;
  assign n441 = n439 ^ x155;
  assign n442 = n432 & n441;
  assign n443 = n442 ^ x27;
  assign n445 = n444 ^ n443;
  assign n447 = n432 & n444;
  assign n448 = ~n439 & n447;
  assign n449 = x27 & x155;
  assign n450 = n449 ^ x156;
  assign n451 = n444 & ~n450;
  assign n452 = n451 ^ x28;
  assign n453 = ~n448 & ~n452;
  assign n446 = x157 ^ x29;
  assign n454 = n453 ^ n446;
  assign n456 = x29 & x157;
  assign n457 = n446 & ~n453;
  assign n458 = ~n456 & ~n457;
  assign n455 = x158 ^ x30;
  assign n459 = n458 ^ n455;
  assign n468 = x159 ^ x31;
  assign n460 = n457 ^ x158;
  assign n461 = n460 ^ x158;
  assign n462 = n456 ^ x158;
  assign n463 = n462 ^ x158;
  assign n464 = ~n461 & ~n463;
  assign n465 = n464 ^ x158;
  assign n466 = n455 & n465;
  assign n467 = n466 ^ x30;
  assign n469 = n468 ^ n467;
  assign n473 = x160 ^ x32;
  assign n470 = n467 ^ x159;
  assign n471 = n468 & ~n470;
  assign n472 = n471 ^ x31;
  assign n474 = n473 ^ n472;
  assign n476 = n468 & n473;
  assign n477 = n467 & n476;
  assign n478 = x31 & x159;
  assign n479 = n478 ^ x160;
  assign n480 = n473 & ~n479;
  assign n481 = n480 ^ x32;
  assign n482 = ~n477 & ~n481;
  assign n475 = x161 ^ x33;
  assign n483 = n482 ^ n475;
  assign n487 = x162 ^ x34;
  assign n484 = n482 ^ x161;
  assign n485 = n475 & n484;
  assign n486 = n485 ^ x33;
  assign n488 = n487 ^ n486;
  assign n490 = n475 & n487;
  assign n491 = ~n482 & n490;
  assign n492 = x33 & x161;
  assign n493 = n492 ^ x162;
  assign n494 = n487 & ~n493;
  assign n495 = n494 ^ x34;
  assign n496 = ~n491 & ~n495;
  assign n489 = x163 ^ x35;
  assign n497 = n496 ^ n489;
  assign n501 = x164 ^ x36;
  assign n498 = n496 ^ x163;
  assign n499 = n489 & n498;
  assign n500 = n499 ^ x35;
  assign n502 = n501 ^ n500;
  assign n504 = n489 & n501;
  assign n505 = ~n496 & n504;
  assign n506 = x35 & x163;
  assign n507 = n506 ^ x164;
  assign n508 = n501 & ~n507;
  assign n509 = n508 ^ x36;
  assign n510 = ~n505 & ~n509;
  assign n503 = x165 ^ x37;
  assign n511 = n510 ^ n503;
  assign n515 = x166 ^ x38;
  assign n512 = n510 ^ x165;
  assign n513 = n503 & n512;
  assign n514 = n513 ^ x37;
  assign n516 = n515 ^ n514;
  assign n518 = n503 & n515;
  assign n519 = ~n510 & n518;
  assign n520 = x37 & x165;
  assign n521 = n520 ^ x166;
  assign n522 = n515 & ~n521;
  assign n523 = n522 ^ x38;
  assign n524 = ~n519 & ~n523;
  assign n517 = x167 ^ x39;
  assign n525 = n524 ^ n517;
  assign n527 = x39 & x167;
  assign n528 = n517 & ~n524;
  assign n529 = ~n527 & ~n528;
  assign n526 = x168 ^ x40;
  assign n530 = n529 ^ n526;
  assign n539 = x169 ^ x41;
  assign n531 = n528 ^ x168;
  assign n532 = n531 ^ x168;
  assign n533 = n527 ^ x168;
  assign n534 = n533 ^ x168;
  assign n535 = ~n532 & ~n534;
  assign n536 = n535 ^ x168;
  assign n537 = n526 & n536;
  assign n538 = n537 ^ x40;
  assign n540 = n539 ^ n538;
  assign n544 = x170 ^ x42;
  assign n541 = n538 ^ x169;
  assign n542 = n539 & ~n541;
  assign n543 = n542 ^ x41;
  assign n545 = n544 ^ n543;
  assign n547 = n539 & n544;
  assign n548 = n538 & n547;
  assign n549 = x41 & x169;
  assign n550 = n549 ^ x170;
  assign n551 = n544 & ~n550;
  assign n552 = n551 ^ x42;
  assign n553 = ~n548 & ~n552;
  assign n546 = x171 ^ x43;
  assign n554 = n553 ^ n546;
  assign n558 = x172 ^ x44;
  assign n555 = n553 ^ x171;
  assign n556 = n546 & n555;
  assign n557 = n556 ^ x43;
  assign n559 = n558 ^ n557;
  assign n561 = n546 & n558;
  assign n562 = ~n553 & n561;
  assign n563 = x43 & x171;
  assign n564 = n563 ^ x172;
  assign n565 = n558 & ~n564;
  assign n566 = n565 ^ x44;
  assign n567 = ~n562 & ~n566;
  assign n560 = x173 ^ x45;
  assign n568 = n567 ^ n560;
  assign n572 = x174 ^ x46;
  assign n569 = n567 ^ x173;
  assign n570 = n560 & n569;
  assign n571 = n570 ^ x45;
  assign n573 = n572 ^ n571;
  assign n575 = n560 & n572;
  assign n576 = ~n567 & n575;
  assign n577 = x45 & x173;
  assign n578 = n577 ^ x174;
  assign n579 = n572 & ~n578;
  assign n580 = n579 ^ x46;
  assign n581 = ~n576 & ~n580;
  assign n574 = x175 ^ x47;
  assign n582 = n581 ^ n574;
  assign n586 = x176 ^ x48;
  assign n583 = n581 ^ x175;
  assign n584 = n574 & n583;
  assign n585 = n584 ^ x47;
  assign n587 = n586 ^ n585;
  assign n589 = n574 & n586;
  assign n590 = ~n581 & n589;
  assign n591 = x47 & x175;
  assign n592 = n591 ^ x176;
  assign n593 = n586 & ~n592;
  assign n594 = n593 ^ x48;
  assign n595 = ~n590 & ~n594;
  assign n588 = x177 ^ x49;
  assign n596 = n595 ^ n588;
  assign n598 = x49 & x177;
  assign n599 = n588 & ~n595;
  assign n600 = ~n598 & ~n599;
  assign n597 = x178 ^ x50;
  assign n601 = n600 ^ n597;
  assign n610 = x179 ^ x51;
  assign n602 = n599 ^ x178;
  assign n603 = n602 ^ x178;
  assign n604 = n598 ^ x178;
  assign n605 = n604 ^ x178;
  assign n606 = ~n603 & ~n605;
  assign n607 = n606 ^ x178;
  assign n608 = n597 & n607;
  assign n609 = n608 ^ x50;
  assign n611 = n610 ^ n609;
  assign n615 = x180 ^ x52;
  assign n612 = n609 ^ x179;
  assign n613 = n610 & ~n612;
  assign n614 = n613 ^ x51;
  assign n616 = n615 ^ n614;
  assign n618 = n610 & n615;
  assign n619 = n609 & n618;
  assign n620 = x51 & x179;
  assign n621 = n620 ^ x180;
  assign n622 = n615 & ~n621;
  assign n623 = n622 ^ x52;
  assign n624 = ~n619 & ~n623;
  assign n617 = x181 ^ x53;
  assign n625 = n624 ^ n617;
  assign n629 = x182 ^ x54;
  assign n626 = n624 ^ x181;
  assign n627 = n617 & n626;
  assign n628 = n627 ^ x53;
  assign n630 = n629 ^ n628;
  assign n632 = n617 & n629;
  assign n633 = ~n624 & n632;
  assign n634 = x53 & x181;
  assign n635 = n634 ^ x182;
  assign n636 = n629 & ~n635;
  assign n637 = n636 ^ x54;
  assign n638 = ~n633 & ~n637;
  assign n631 = x183 ^ x55;
  assign n639 = n638 ^ n631;
  assign n643 = x184 ^ x56;
  assign n640 = n638 ^ x183;
  assign n641 = n631 & n640;
  assign n642 = n641 ^ x55;
  assign n644 = n643 ^ n642;
  assign n646 = n631 & n643;
  assign n647 = ~n638 & n646;
  assign n648 = x55 & x183;
  assign n649 = n648 ^ x184;
  assign n650 = n643 & ~n649;
  assign n651 = n650 ^ x56;
  assign n652 = ~n647 & ~n651;
  assign n645 = x185 ^ x57;
  assign n653 = n652 ^ n645;
  assign n657 = x186 ^ x58;
  assign n654 = n652 ^ x185;
  assign n655 = n645 & n654;
  assign n656 = n655 ^ x57;
  assign n658 = n657 ^ n656;
  assign n660 = n645 & n657;
  assign n661 = ~n652 & n660;
  assign n662 = x57 & x185;
  assign n663 = n662 ^ x186;
  assign n664 = n657 & ~n663;
  assign n665 = n664 ^ x58;
  assign n666 = ~n661 & ~n665;
  assign n659 = x187 ^ x59;
  assign n667 = n666 ^ n659;
  assign n669 = x59 & x187;
  assign n670 = n659 & ~n666;
  assign n671 = ~n669 & ~n670;
  assign n668 = x188 ^ x60;
  assign n672 = n671 ^ n668;
  assign n681 = x189 ^ x61;
  assign n673 = n670 ^ x188;
  assign n674 = n673 ^ x188;
  assign n675 = n669 ^ x188;
  assign n676 = n675 ^ x188;
  assign n677 = ~n674 & ~n676;
  assign n678 = n677 ^ x188;
  assign n679 = n668 & n678;
  assign n680 = n679 ^ x60;
  assign n682 = n681 ^ n680;
  assign n686 = x190 ^ x62;
  assign n683 = n680 ^ x189;
  assign n684 = n681 & ~n683;
  assign n685 = n684 ^ x61;
  assign n687 = n686 ^ n685;
  assign n689 = n681 & n686;
  assign n690 = n680 & n689;
  assign n691 = x61 & x189;
  assign n692 = n691 ^ x190;
  assign n693 = n686 & ~n692;
  assign n694 = n693 ^ x62;
  assign n695 = ~n690 & ~n694;
  assign n688 = x191 ^ x63;
  assign n696 = n695 ^ n688;
  assign n700 = x192 ^ x64;
  assign n697 = n695 ^ x191;
  assign n698 = n688 & n697;
  assign n699 = n698 ^ x63;
  assign n701 = n700 ^ n699;
  assign n703 = n688 & n700;
  assign n704 = ~n695 & n703;
  assign n705 = x63 & x191;
  assign n706 = n705 ^ x192;
  assign n707 = n700 & ~n706;
  assign n708 = n707 ^ x64;
  assign n709 = ~n704 & ~n708;
  assign n702 = x193 ^ x65;
  assign n710 = n709 ^ n702;
  assign n714 = x194 ^ x66;
  assign n711 = n709 ^ x193;
  assign n712 = n702 & n711;
  assign n713 = n712 ^ x65;
  assign n715 = n714 ^ n713;
  assign n717 = n702 & n714;
  assign n718 = ~n709 & n717;
  assign n719 = x65 & x193;
  assign n720 = n719 ^ x194;
  assign n721 = n714 & ~n720;
  assign n722 = n721 ^ x66;
  assign n723 = ~n718 & ~n722;
  assign n716 = x195 ^ x67;
  assign n724 = n723 ^ n716;
  assign n728 = x196 ^ x68;
  assign n725 = n723 ^ x195;
  assign n726 = n716 & n725;
  assign n727 = n726 ^ x67;
  assign n729 = n728 ^ n727;
  assign n731 = n716 & n728;
  assign n732 = ~n723 & n731;
  assign n733 = x67 & x195;
  assign n734 = n733 ^ x196;
  assign n735 = n728 & ~n734;
  assign n736 = n735 ^ x68;
  assign n737 = ~n732 & ~n736;
  assign n730 = x197 ^ x69;
  assign n738 = n737 ^ n730;
  assign n740 = x69 & x197;
  assign n741 = n730 & ~n737;
  assign n742 = ~n740 & ~n741;
  assign n739 = x198 ^ x70;
  assign n743 = n742 ^ n739;
  assign n752 = x199 ^ x71;
  assign n744 = n741 ^ x198;
  assign n745 = n744 ^ x198;
  assign n746 = n740 ^ x198;
  assign n747 = n746 ^ x198;
  assign n748 = ~n745 & ~n747;
  assign n749 = n748 ^ x198;
  assign n750 = n739 & n749;
  assign n751 = n750 ^ x70;
  assign n753 = n752 ^ n751;
  assign n757 = x200 ^ x72;
  assign n754 = n751 ^ x199;
  assign n755 = n752 & ~n754;
  assign n756 = n755 ^ x71;
  assign n758 = n757 ^ n756;
  assign n760 = n752 & n757;
  assign n761 = n751 & n760;
  assign n762 = x71 & x199;
  assign n763 = n762 ^ x200;
  assign n764 = n757 & ~n763;
  assign n765 = n764 ^ x72;
  assign n766 = ~n761 & ~n765;
  assign n759 = x201 ^ x73;
  assign n767 = n766 ^ n759;
  assign n771 = x202 ^ x74;
  assign n768 = n766 ^ x201;
  assign n769 = n759 & n768;
  assign n770 = n769 ^ x73;
  assign n772 = n771 ^ n770;
  assign n774 = n759 & n771;
  assign n775 = ~n766 & n774;
  assign n776 = x73 & x201;
  assign n777 = n776 ^ x202;
  assign n778 = n771 & ~n777;
  assign n779 = n778 ^ x74;
  assign n780 = ~n775 & ~n779;
  assign n773 = x203 ^ x75;
  assign n781 = n780 ^ n773;
  assign n785 = x204 ^ x76;
  assign n782 = n780 ^ x203;
  assign n783 = n773 & n782;
  assign n784 = n783 ^ x75;
  assign n786 = n785 ^ n784;
  assign n788 = n773 & n785;
  assign n789 = ~n780 & n788;
  assign n790 = x75 & x203;
  assign n791 = n790 ^ x204;
  assign n792 = n785 & ~n791;
  assign n793 = n792 ^ x76;
  assign n794 = ~n789 & ~n793;
  assign n787 = x205 ^ x77;
  assign n795 = n794 ^ n787;
  assign n799 = x206 ^ x78;
  assign n796 = n794 ^ x205;
  assign n797 = n787 & n796;
  assign n798 = n797 ^ x77;
  assign n800 = n799 ^ n798;
  assign n802 = n787 & n799;
  assign n803 = ~n794 & n802;
  assign n804 = x77 & x205;
  assign n805 = n804 ^ x206;
  assign n806 = n799 & ~n805;
  assign n807 = n806 ^ x78;
  assign n808 = ~n803 & ~n807;
  assign n801 = x207 ^ x79;
  assign n809 = n808 ^ n801;
  assign n811 = x79 & x207;
  assign n812 = n801 & ~n808;
  assign n813 = ~n811 & ~n812;
  assign n810 = x208 ^ x80;
  assign n814 = n813 ^ n810;
  assign n823 = x209 ^ x81;
  assign n815 = n812 ^ x208;
  assign n816 = n815 ^ x208;
  assign n817 = n811 ^ x208;
  assign n818 = n817 ^ x208;
  assign n819 = ~n816 & ~n818;
  assign n820 = n819 ^ x208;
  assign n821 = n810 & n820;
  assign n822 = n821 ^ x80;
  assign n824 = n823 ^ n822;
  assign n828 = x210 ^ x82;
  assign n825 = n822 ^ x209;
  assign n826 = n823 & ~n825;
  assign n827 = n826 ^ x81;
  assign n829 = n828 ^ n827;
  assign n831 = n823 & n828;
  assign n832 = n822 & n831;
  assign n833 = x81 & x209;
  assign n834 = n833 ^ x210;
  assign n835 = n828 & ~n834;
  assign n836 = n835 ^ x82;
  assign n837 = ~n832 & ~n836;
  assign n830 = x211 ^ x83;
  assign n838 = n837 ^ n830;
  assign n842 = x212 ^ x84;
  assign n839 = n837 ^ x211;
  assign n840 = n830 & n839;
  assign n841 = n840 ^ x83;
  assign n843 = n842 ^ n841;
  assign n845 = n830 & n842;
  assign n846 = ~n837 & n845;
  assign n847 = x83 & x211;
  assign n848 = n847 ^ x212;
  assign n849 = n842 & ~n848;
  assign n850 = n849 ^ x84;
  assign n851 = ~n846 & ~n850;
  assign n844 = x213 ^ x85;
  assign n852 = n851 ^ n844;
  assign n856 = x214 ^ x86;
  assign n853 = n851 ^ x213;
  assign n854 = n844 & n853;
  assign n855 = n854 ^ x85;
  assign n857 = n856 ^ n855;
  assign n859 = n844 & n856;
  assign n860 = ~n851 & n859;
  assign n861 = x85 & x213;
  assign n862 = n861 ^ x214;
  assign n863 = n856 & ~n862;
  assign n864 = n863 ^ x86;
  assign n865 = ~n860 & ~n864;
  assign n858 = x215 ^ x87;
  assign n866 = n865 ^ n858;
  assign n870 = x216 ^ x88;
  assign n867 = n865 ^ x215;
  assign n868 = n858 & n867;
  assign n869 = n868 ^ x87;
  assign n871 = n870 ^ n869;
  assign n873 = n858 & n870;
  assign n874 = ~n865 & n873;
  assign n875 = x87 & x215;
  assign n876 = n875 ^ x216;
  assign n877 = n870 & ~n876;
  assign n878 = n877 ^ x88;
  assign n879 = ~n874 & ~n878;
  assign n872 = x217 ^ x89;
  assign n880 = n879 ^ n872;
  assign n882 = x89 & x217;
  assign n883 = n872 & ~n879;
  assign n884 = ~n882 & ~n883;
  assign n881 = x218 ^ x90;
  assign n885 = n884 ^ n881;
  assign n894 = x219 ^ x91;
  assign n886 = n883 ^ x218;
  assign n887 = n886 ^ x218;
  assign n888 = n882 ^ x218;
  assign n889 = n888 ^ x218;
  assign n890 = ~n887 & ~n889;
  assign n891 = n890 ^ x218;
  assign n892 = n881 & n891;
  assign n893 = n892 ^ x90;
  assign n895 = n894 ^ n893;
  assign n897 = x91 & x219;
  assign n898 = n893 & n894;
  assign n899 = ~n897 & ~n898;
  assign n896 = x220 ^ x92;
  assign n900 = n899 ^ n896;
  assign n909 = x221 ^ x93;
  assign n901 = n898 ^ x220;
  assign n902 = n901 ^ x220;
  assign n903 = n897 ^ x220;
  assign n904 = n903 ^ x220;
  assign n905 = ~n902 & ~n904;
  assign n906 = n905 ^ x220;
  assign n907 = n896 & n906;
  assign n908 = n907 ^ x92;
  assign n910 = n909 ^ n908;
  assign n914 = x222 ^ x94;
  assign n911 = n908 ^ x221;
  assign n912 = n909 & ~n911;
  assign n913 = n912 ^ x93;
  assign n915 = n914 ^ n913;
  assign n919 = x223 ^ x95;
  assign n916 = n913 ^ x222;
  assign n917 = n914 & ~n916;
  assign n918 = n917 ^ x94;
  assign n920 = n919 ^ n918;
  assign n924 = x224 ^ x96;
  assign n921 = n918 ^ x223;
  assign n922 = n919 & ~n921;
  assign n923 = n922 ^ x95;
  assign n925 = n924 ^ n923;
  assign n929 = x225 ^ x97;
  assign n926 = n923 ^ x224;
  assign n927 = n924 & ~n926;
  assign n928 = n927 ^ x96;
  assign n930 = n929 ^ n928;
  assign n934 = x226 ^ x98;
  assign n931 = n928 ^ x225;
  assign n932 = n929 & ~n931;
  assign n933 = n932 ^ x97;
  assign n935 = n934 ^ n933;
  assign n937 = n929 & n934;
  assign n938 = n928 & n937;
  assign n939 = x97 & x225;
  assign n940 = n939 ^ x226;
  assign n941 = n934 & ~n940;
  assign n942 = n941 ^ x98;
  assign n943 = ~n938 & ~n942;
  assign n936 = x227 ^ x99;
  assign n944 = n943 ^ n936;
  assign n948 = x228 ^ x100;
  assign n945 = n943 ^ x227;
  assign n946 = n936 & n945;
  assign n947 = n946 ^ x99;
  assign n949 = n948 ^ n947;
  assign n951 = n936 & n948;
  assign n952 = ~n943 & n951;
  assign n953 = x99 & x227;
  assign n954 = n953 ^ x228;
  assign n955 = n948 & ~n954;
  assign n956 = n955 ^ x100;
  assign n957 = ~n952 & ~n956;
  assign n950 = x229 ^ x101;
  assign n958 = n957 ^ n950;
  assign n962 = x230 ^ x102;
  assign n959 = n957 ^ x229;
  assign n960 = n950 & n959;
  assign n961 = n960 ^ x101;
  assign n963 = n962 ^ n961;
  assign n965 = n950 & n962;
  assign n966 = ~n957 & n965;
  assign n967 = x101 & x229;
  assign n968 = n967 ^ x230;
  assign n969 = n962 & ~n968;
  assign n970 = n969 ^ x102;
  assign n971 = ~n966 & ~n970;
  assign n964 = x231 ^ x103;
  assign n972 = n971 ^ n964;
  assign n976 = x232 ^ x104;
  assign n973 = n971 ^ x231;
  assign n974 = n964 & n973;
  assign n975 = n974 ^ x103;
  assign n977 = n976 ^ n975;
  assign n981 = x233 ^ x105;
  assign n978 = n975 ^ x232;
  assign n979 = n976 & ~n978;
  assign n980 = n979 ^ x104;
  assign n982 = n981 ^ n980;
  assign n986 = x234 ^ x106;
  assign n983 = n980 ^ x233;
  assign n984 = n981 & ~n983;
  assign n985 = n984 ^ x105;
  assign n987 = n986 ^ n985;
  assign n989 = n981 & n986;
  assign n990 = n980 & n989;
  assign n991 = x105 & x233;
  assign n992 = n991 ^ x234;
  assign n993 = n986 & ~n992;
  assign n994 = n993 ^ x106;
  assign n995 = ~n990 & ~n994;
  assign n988 = x235 ^ x107;
  assign n996 = n995 ^ n988;
  assign n1000 = x236 ^ x108;
  assign n997 = n995 ^ x235;
  assign n998 = n988 & n997;
  assign n999 = n998 ^ x107;
  assign n1001 = n1000 ^ n999;
  assign n1005 = x237 ^ x109;
  assign n1002 = n999 ^ x236;
  assign n1003 = n1000 & ~n1002;
  assign n1004 = n1003 ^ x108;
  assign n1006 = n1005 ^ n1004;
  assign n1010 = x238 ^ x110;
  assign n1007 = n1004 ^ x237;
  assign n1008 = n1005 & ~n1007;
  assign n1009 = n1008 ^ x109;
  assign n1011 = n1010 ^ n1009;
  assign n1013 = n1005 & n1010;
  assign n1014 = n1004 & n1013;
  assign n1015 = x109 & x237;
  assign n1016 = n1015 ^ x238;
  assign n1017 = n1010 & ~n1016;
  assign n1018 = n1017 ^ x110;
  assign n1019 = ~n1014 & ~n1018;
  assign n1012 = x239 ^ x111;
  assign n1020 = n1019 ^ n1012;
  assign n1024 = x240 ^ x112;
  assign n1021 = n1019 ^ x239;
  assign n1022 = n1012 & n1021;
  assign n1023 = n1022 ^ x111;
  assign n1025 = n1024 ^ n1023;
  assign n1029 = x241 ^ x113;
  assign n1026 = n1023 ^ x240;
  assign n1027 = n1024 & ~n1026;
  assign n1028 = n1027 ^ x112;
  assign n1030 = n1029 ^ n1028;
  assign n1034 = x242 ^ x114;
  assign n1031 = n1028 ^ x241;
  assign n1032 = n1029 & ~n1031;
  assign n1033 = n1032 ^ x113;
  assign n1035 = n1034 ^ n1033;
  assign n1039 = x243 ^ x115;
  assign n1036 = n1033 ^ x242;
  assign n1037 = n1034 & ~n1036;
  assign n1038 = n1037 ^ x114;
  assign n1040 = n1039 ^ n1038;
  assign n1044 = x244 ^ x116;
  assign n1041 = n1038 ^ x243;
  assign n1042 = n1039 & ~n1041;
  assign n1043 = n1042 ^ x115;
  assign n1045 = n1044 ^ n1043;
  assign n1049 = x245 ^ x117;
  assign n1046 = n1043 ^ x244;
  assign n1047 = n1044 & ~n1046;
  assign n1048 = n1047 ^ x116;
  assign n1050 = n1049 ^ n1048;
  assign n1054 = x246 ^ x118;
  assign n1051 = n1048 ^ x245;
  assign n1052 = n1049 & ~n1051;
  assign n1053 = n1052 ^ x117;
  assign n1055 = n1054 ^ n1053;
  assign n1059 = x247 ^ x119;
  assign n1056 = n1053 ^ x246;
  assign n1057 = n1054 & ~n1056;
  assign n1058 = n1057 ^ x118;
  assign n1060 = n1059 ^ n1058;
  assign n1064 = x248 ^ x120;
  assign n1061 = n1058 ^ x247;
  assign n1062 = n1059 & ~n1061;
  assign n1063 = n1062 ^ x119;
  assign n1065 = n1064 ^ n1063;
  assign n1069 = x249 ^ x121;
  assign n1066 = n1063 ^ x248;
  assign n1067 = n1064 & ~n1066;
  assign n1068 = n1067 ^ x120;
  assign n1070 = n1069 ^ n1068;
  assign n1074 = x250 ^ x122;
  assign n1071 = n1068 ^ x249;
  assign n1072 = n1069 & ~n1071;
  assign n1073 = n1072 ^ x121;
  assign n1075 = n1074 ^ n1073;
  assign n1079 = x251 ^ x123;
  assign n1076 = n1073 ^ x250;
  assign n1077 = n1074 & ~n1076;
  assign n1078 = n1077 ^ x122;
  assign n1080 = n1079 ^ n1078;
  assign n1084 = x252 ^ x124;
  assign n1081 = n1078 ^ x251;
  assign n1082 = n1079 & ~n1081;
  assign n1083 = n1082 ^ x123;
  assign n1085 = n1084 ^ n1083;
  assign n1089 = x253 ^ x125;
  assign n1086 = n1083 ^ x252;
  assign n1087 = n1084 & ~n1086;
  assign n1088 = n1087 ^ x124;
  assign n1090 = n1089 ^ n1088;
  assign n1094 = x254 ^ x126;
  assign n1091 = n1088 ^ x253;
  assign n1092 = n1089 & ~n1091;
  assign n1093 = n1092 ^ x125;
  assign n1095 = n1094 ^ n1093;
  assign n1099 = x255 ^ x127;
  assign n1096 = n1093 ^ x254;
  assign n1097 = n1094 & ~n1096;
  assign n1098 = n1097 ^ x126;
  assign n1100 = n1099 ^ n1098;
  assign n1101 = n1098 ^ x255;
  assign n1102 = n1099 & ~n1101;
  assign n1103 = n1102 ^ x127;
  assign y0 = n257;
  assign y1 = n260;
  assign y2 = n265;
  assign y3 = n270;
  assign y4 = n275;
  assign y5 = ~n284;
  assign y6 = n289;
  assign y7 = ~n298;
  assign y8 = n303;
  assign y9 = ~n312;
  assign y10 = ~n317;
  assign y11 = n327;
  assign y12 = n332;
  assign y13 = ~n341;
  assign y14 = n346;
  assign y15 = ~n355;
  assign y16 = n360;
  assign y17 = ~n369;
  assign y18 = n374;
  assign y19 = ~n383;
  assign y20 = ~n388;
  assign y21 = n398;
  assign y22 = n403;
  assign y23 = ~n412;
  assign y24 = n417;
  assign y25 = ~n426;
  assign y26 = n431;
  assign y27 = ~n440;
  assign y28 = n445;
  assign y29 = ~n454;
  assign y30 = ~n459;
  assign y31 = n469;
  assign y32 = n474;
  assign y33 = ~n483;
  assign y34 = n488;
  assign y35 = ~n497;
  assign y36 = n502;
  assign y37 = ~n511;
  assign y38 = n516;
  assign y39 = ~n525;
  assign y40 = ~n530;
  assign y41 = n540;
  assign y42 = n545;
  assign y43 = ~n554;
  assign y44 = n559;
  assign y45 = ~n568;
  assign y46 = n573;
  assign y47 = ~n582;
  assign y48 = n587;
  assign y49 = ~n596;
  assign y50 = ~n601;
  assign y51 = n611;
  assign y52 = n616;
  assign y53 = ~n625;
  assign y54 = n630;
  assign y55 = ~n639;
  assign y56 = n644;
  assign y57 = ~n653;
  assign y58 = n658;
  assign y59 = ~n667;
  assign y60 = ~n672;
  assign y61 = n682;
  assign y62 = n687;
  assign y63 = ~n696;
  assign y64 = n701;
  assign y65 = ~n710;
  assign y66 = n715;
  assign y67 = ~n724;
  assign y68 = n729;
  assign y69 = ~n738;
  assign y70 = ~n743;
  assign y71 = n753;
  assign y72 = n758;
  assign y73 = ~n767;
  assign y74 = n772;
  assign y75 = ~n781;
  assign y76 = n786;
  assign y77 = ~n795;
  assign y78 = n800;
  assign y79 = ~n809;
  assign y80 = ~n814;
  assign y81 = n824;
  assign y82 = n829;
  assign y83 = ~n838;
  assign y84 = n843;
  assign y85 = ~n852;
  assign y86 = n857;
  assign y87 = ~n866;
  assign y88 = n871;
  assign y89 = ~n880;
  assign y90 = ~n885;
  assign y91 = n895;
  assign y92 = ~n900;
  assign y93 = n910;
  assign y94 = n915;
  assign y95 = n920;
  assign y96 = n925;
  assign y97 = n930;
  assign y98 = n935;
  assign y99 = ~n944;
  assign y100 = n949;
  assign y101 = ~n958;
  assign y102 = n963;
  assign y103 = ~n972;
  assign y104 = n977;
  assign y105 = n982;
  assign y106 = n987;
  assign y107 = ~n996;
  assign y108 = n1001;
  assign y109 = n1006;
  assign y110 = n1011;
  assign y111 = ~n1020;
  assign y112 = n1025;
  assign y113 = n1030;
  assign y114 = n1035;
  assign y115 = n1040;
  assign y116 = n1045;
  assign y117 = n1050;
  assign y118 = n1055;
  assign y119 = n1060;
  assign y120 = n1065;
  assign y121 = n1070;
  assign y122 = n1075;
  assign y123 = n1080;
  assign y124 = n1085;
  assign y125 = n1090;
  assign y126 = n1095;
  assign y127 = n1100;
  assign y128 = n1103;
endmodule
