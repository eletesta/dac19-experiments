module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64;
  wire n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488;
  assign n129 = x64 ^ x0;
  assign n131 = x0 & x64;
  assign n130 = x65 ^ x1;
  assign n132 = n131 ^ n130;
  assign n133 = x1 & x65;
  assign n134 = ~x1 & ~x65;
  assign n135 = n131 & ~n134;
  assign n136 = ~n133 & ~n135;
  assign n137 = n136 ^ x2;
  assign n138 = n137 ^ x66;
  assign n139 = x66 ^ x2;
  assign n140 = n136 ^ x66;
  assign n141 = n139 & n140;
  assign n142 = n141 ^ x2;
  assign n143 = n142 ^ x67;
  assign n144 = n143 ^ x3;
  assign n145 = x67 ^ x3;
  assign n146 = ~n143 & n145;
  assign n147 = n146 ^ x3;
  assign n148 = n147 ^ x4;
  assign n149 = n148 ^ x68;
  assign n150 = x68 ^ x4;
  assign n151 = n147 ^ x68;
  assign n152 = n150 & ~n151;
  assign n153 = n152 ^ x4;
  assign n154 = n153 ^ x5;
  assign n155 = n154 ^ x69;
  assign n156 = x69 ^ x5;
  assign n157 = n153 ^ x69;
  assign n158 = n156 & ~n157;
  assign n159 = n158 ^ x5;
  assign n160 = n159 ^ x6;
  assign n161 = n160 ^ x70;
  assign n162 = x70 ^ x6;
  assign n163 = n159 ^ x70;
  assign n164 = n162 & ~n163;
  assign n165 = n164 ^ x6;
  assign n166 = n165 ^ x7;
  assign n167 = n166 ^ x71;
  assign n168 = x71 ^ x7;
  assign n169 = n165 ^ x71;
  assign n170 = n168 & ~n169;
  assign n171 = n170 ^ x7;
  assign n172 = n171 ^ x8;
  assign n173 = n172 ^ x72;
  assign n174 = x72 ^ x8;
  assign n175 = n171 ^ x72;
  assign n176 = n174 & ~n175;
  assign n177 = n176 ^ x8;
  assign n178 = n177 ^ x9;
  assign n179 = n178 ^ x73;
  assign n180 = x73 ^ x9;
  assign n181 = n177 ^ x73;
  assign n182 = n180 & ~n181;
  assign n183 = n182 ^ x9;
  assign n184 = n183 ^ x10;
  assign n185 = n184 ^ x74;
  assign n186 = x74 ^ x10;
  assign n187 = n183 ^ x74;
  assign n188 = n186 & ~n187;
  assign n189 = n188 ^ x10;
  assign n190 = n189 ^ x11;
  assign n191 = n190 ^ x75;
  assign n192 = x75 ^ x11;
  assign n193 = n189 ^ x75;
  assign n194 = n192 & ~n193;
  assign n195 = n194 ^ x11;
  assign n196 = n195 ^ x12;
  assign n197 = n196 ^ x76;
  assign n198 = x76 ^ x12;
  assign n199 = n195 ^ x76;
  assign n200 = n198 & ~n199;
  assign n201 = n200 ^ x12;
  assign n202 = n201 ^ x13;
  assign n203 = n202 ^ x77;
  assign n204 = x77 ^ x13;
  assign n205 = n201 ^ x77;
  assign n206 = n204 & ~n205;
  assign n207 = n206 ^ x13;
  assign n208 = n207 ^ x14;
  assign n209 = n208 ^ x78;
  assign n210 = x78 ^ x14;
  assign n211 = n207 ^ x78;
  assign n212 = n210 & ~n211;
  assign n213 = n212 ^ x14;
  assign n214 = n213 ^ x15;
  assign n215 = n214 ^ x79;
  assign n216 = x79 ^ x15;
  assign n217 = n213 ^ x79;
  assign n218 = n216 & ~n217;
  assign n219 = n218 ^ x15;
  assign n220 = n219 ^ x80;
  assign n221 = n220 ^ x16;
  assign n222 = x80 ^ x16;
  assign n223 = ~n220 & n222;
  assign n224 = n223 ^ x16;
  assign n225 = n224 ^ x17;
  assign n226 = n225 ^ x81;
  assign n227 = x81 ^ x17;
  assign n228 = n224 ^ x81;
  assign n229 = n227 & ~n228;
  assign n230 = n229 ^ x17;
  assign n231 = n230 ^ x82;
  assign n232 = n231 ^ x18;
  assign n233 = x82 ^ x18;
  assign n234 = ~n231 & n233;
  assign n235 = n234 ^ x18;
  assign n236 = n235 ^ x19;
  assign n237 = n236 ^ x83;
  assign n238 = x83 ^ x19;
  assign n239 = n235 ^ x83;
  assign n240 = n238 & ~n239;
  assign n241 = n240 ^ x19;
  assign n242 = n241 ^ x20;
  assign n243 = n242 ^ x84;
  assign n244 = x84 ^ x20;
  assign n245 = n241 ^ x84;
  assign n246 = n244 & ~n245;
  assign n247 = n246 ^ x20;
  assign n248 = n247 ^ x21;
  assign n249 = n248 ^ x85;
  assign n250 = x85 ^ x21;
  assign n251 = n247 ^ x85;
  assign n252 = n250 & ~n251;
  assign n253 = n252 ^ x21;
  assign n254 = n253 ^ x22;
  assign n255 = n254 ^ x86;
  assign n256 = x86 ^ x22;
  assign n257 = n253 ^ x86;
  assign n258 = n256 & ~n257;
  assign n259 = n258 ^ x22;
  assign n260 = n259 ^ x87;
  assign n261 = n260 ^ x23;
  assign n262 = x87 ^ x23;
  assign n263 = ~n260 & n262;
  assign n264 = n263 ^ x23;
  assign n265 = n264 ^ x88;
  assign n266 = n265 ^ x24;
  assign n267 = x88 ^ x24;
  assign n268 = ~n265 & n267;
  assign n269 = n268 ^ x24;
  assign n270 = n269 ^ x25;
  assign n271 = n270 ^ x89;
  assign n272 = x89 ^ x25;
  assign n273 = n269 ^ x89;
  assign n274 = n272 & ~n273;
  assign n275 = n274 ^ x25;
  assign n276 = n275 ^ x26;
  assign n277 = n276 ^ x90;
  assign n278 = x90 ^ x26;
  assign n279 = n275 ^ x90;
  assign n280 = n278 & ~n279;
  assign n281 = n280 ^ x26;
  assign n282 = n281 ^ x27;
  assign n283 = n282 ^ x91;
  assign n284 = x91 ^ x27;
  assign n285 = n281 ^ x91;
  assign n286 = n284 & ~n285;
  assign n287 = n286 ^ x27;
  assign n288 = n287 ^ x28;
  assign n289 = n288 ^ x92;
  assign n290 = x92 ^ x28;
  assign n291 = n287 ^ x92;
  assign n292 = n290 & ~n291;
  assign n293 = n292 ^ x28;
  assign n294 = n293 ^ x93;
  assign n295 = n294 ^ x29;
  assign n296 = x93 ^ x29;
  assign n297 = ~n294 & n296;
  assign n298 = n297 ^ x29;
  assign n299 = n298 ^ x30;
  assign n300 = n299 ^ x94;
  assign n301 = x94 ^ x30;
  assign n302 = n298 ^ x94;
  assign n303 = n301 & ~n302;
  assign n304 = n303 ^ x30;
  assign n305 = n304 ^ x31;
  assign n306 = n305 ^ x95;
  assign n308 = x95 ^ x31;
  assign n309 = n304 ^ x95;
  assign n310 = n308 & ~n309;
  assign n311 = n310 ^ x31;
  assign n307 = x96 ^ x32;
  assign n312 = n311 ^ n307;
  assign n313 = x32 & x96;
  assign n314 = ~x32 & ~x96;
  assign n315 = n311 & ~n314;
  assign n316 = ~n313 & ~n315;
  assign n317 = n316 ^ x97;
  assign n318 = n317 ^ x33;
  assign n320 = x97 ^ x33;
  assign n321 = n317 & n320;
  assign n322 = n321 ^ x33;
  assign n319 = x98 ^ x34;
  assign n323 = n322 ^ n319;
  assign n325 = x34 & x98;
  assign n326 = ~x34 & ~x98;
  assign n327 = n322 & ~n326;
  assign n328 = ~n325 & ~n327;
  assign n324 = x99 ^ x35;
  assign n329 = n328 ^ n324;
  assign n330 = x35 & x99;
  assign n331 = ~x35 & ~x99;
  assign n332 = ~n328 & ~n331;
  assign n333 = ~n330 & ~n332;
  assign n334 = n333 ^ x100;
  assign n335 = n334 ^ x36;
  assign n337 = x100 ^ x36;
  assign n338 = n334 & n337;
  assign n339 = n338 ^ x36;
  assign n336 = x101 ^ x37;
  assign n340 = n339 ^ n336;
  assign n341 = x37 & x101;
  assign n342 = ~x37 & ~x101;
  assign n343 = n339 & ~n342;
  assign n344 = ~n341 & ~n343;
  assign n345 = n344 ^ x38;
  assign n346 = n345 ^ x102;
  assign n347 = x102 ^ x38;
  assign n348 = n344 ^ x102;
  assign n349 = n347 & n348;
  assign n350 = n349 ^ x38;
  assign n351 = n350 ^ x39;
  assign n352 = n351 ^ x103;
  assign n353 = x103 ^ x39;
  assign n354 = n350 ^ x103;
  assign n355 = n353 & ~n354;
  assign n356 = n355 ^ x39;
  assign n357 = n356 ^ x104;
  assign n358 = n357 ^ x40;
  assign n359 = x104 ^ x40;
  assign n360 = ~n357 & n359;
  assign n361 = n360 ^ x40;
  assign n362 = n361 ^ x41;
  assign n363 = n362 ^ x105;
  assign n364 = x105 ^ x41;
  assign n365 = n361 ^ x105;
  assign n366 = n364 & ~n365;
  assign n367 = n366 ^ x41;
  assign n368 = n367 ^ x106;
  assign n369 = n368 ^ x42;
  assign n370 = x106 ^ x42;
  assign n371 = ~n368 & n370;
  assign n372 = n371 ^ x42;
  assign n373 = n372 ^ x43;
  assign n374 = n373 ^ x107;
  assign n375 = x107 ^ x43;
  assign n376 = n372 ^ x107;
  assign n377 = n375 & ~n376;
  assign n378 = n377 ^ x43;
  assign n379 = n378 ^ x108;
  assign n380 = n379 ^ x44;
  assign n381 = x108 ^ x44;
  assign n382 = ~n379 & n381;
  assign n383 = n382 ^ x44;
  assign n384 = n383 ^ x109;
  assign n385 = n384 ^ x45;
  assign n386 = x109 ^ x45;
  assign n387 = ~n384 & n386;
  assign n388 = n387 ^ x45;
  assign n389 = n388 ^ x46;
  assign n390 = n389 ^ x110;
  assign n391 = x110 ^ x46;
  assign n392 = n388 ^ x110;
  assign n393 = n391 & ~n392;
  assign n394 = n393 ^ x46;
  assign n395 = n394 ^ x47;
  assign n396 = n395 ^ x111;
  assign n401 = x112 ^ x48;
  assign n397 = x111 ^ x47;
  assign n398 = n394 ^ x111;
  assign n399 = n397 & ~n398;
  assign n400 = n399 ^ x47;
  assign n402 = n401 ^ n400;
  assign n406 = x113 ^ x49;
  assign n403 = n400 ^ x112;
  assign n404 = n401 & ~n403;
  assign n405 = n404 ^ x48;
  assign n407 = n406 ^ n405;
  assign n411 = x114 ^ x50;
  assign n408 = n405 ^ x113;
  assign n409 = n406 & ~n408;
  assign n410 = n409 ^ x49;
  assign n412 = n411 ^ n410;
  assign n414 = n410 ^ x114;
  assign n415 = n411 & ~n414;
  assign n416 = n415 ^ x50;
  assign n413 = x115 ^ x51;
  assign n417 = n416 ^ n413;
  assign n422 = x116 ^ x52;
  assign n418 = ~x51 & ~x115;
  assign n419 = x51 & x115;
  assign n420 = ~n416 & ~n419;
  assign n421 = ~n418 & ~n420;
  assign n423 = n422 ^ n421;
  assign n427 = x117 ^ x53;
  assign n424 = n421 ^ x116;
  assign n425 = n422 & ~n424;
  assign n426 = n425 ^ x52;
  assign n428 = n427 ^ n426;
  assign n432 = x118 ^ x54;
  assign n429 = n426 ^ x117;
  assign n430 = n427 & ~n429;
  assign n431 = n430 ^ x53;
  assign n433 = n432 ^ n431;
  assign n435 = n431 ^ x118;
  assign n436 = n432 & ~n435;
  assign n437 = n436 ^ x54;
  assign n434 = x119 ^ x55;
  assign n438 = n437 ^ n434;
  assign n443 = x120 ^ x56;
  assign n439 = ~x55 & ~x119;
  assign n440 = x55 & x119;
  assign n441 = ~n437 & ~n440;
  assign n442 = ~n439 & ~n441;
  assign n444 = n443 ^ n442;
  assign n445 = n442 ^ x120;
  assign n446 = n443 & ~n445;
  assign n447 = n446 ^ x56;
  assign n448 = n447 ^ x57;
  assign n449 = n448 ^ x121;
  assign n454 = x122 ^ x58;
  assign n450 = x121 ^ x57;
  assign n451 = n447 ^ x121;
  assign n452 = n450 & ~n451;
  assign n453 = n452 ^ x57;
  assign n455 = n454 ^ n453;
  assign n457 = n453 ^ x122;
  assign n458 = n454 & ~n457;
  assign n459 = n458 ^ x58;
  assign n456 = x123 ^ x59;
  assign n460 = n459 ^ n456;
  assign n462 = x59 & x123;
  assign n463 = ~x59 & ~x123;
  assign n464 = n459 & ~n463;
  assign n465 = ~n462 & ~n464;
  assign n461 = x124 ^ x60;
  assign n466 = n465 ^ n461;
  assign n468 = x60 & x124;
  assign n469 = ~x60 & ~x124;
  assign n470 = ~n465 & ~n469;
  assign n471 = ~n468 & ~n470;
  assign n467 = x125 ^ x61;
  assign n472 = n471 ^ n467;
  assign n474 = x61 & x125;
  assign n475 = ~x61 & ~x125;
  assign n476 = ~n471 & ~n475;
  assign n477 = ~n474 & ~n476;
  assign n473 = x126 ^ x62;
  assign n478 = n477 ^ n473;
  assign n480 = x62 & x126;
  assign n481 = ~x62 & ~x126;
  assign n482 = ~n477 & ~n481;
  assign n483 = ~n480 & ~n482;
  assign n479 = x127 ^ x63;
  assign n484 = n483 ^ n479;
  assign n485 = x63 & x127;
  assign n486 = ~x63 & ~x127;
  assign n487 = ~n483 & ~n486;
  assign n488 = ~n485 & ~n487;
  assign y0 = n129;
  assign y1 = n132;
  assign y2 = ~n138;
  assign y3 = n144;
  assign y4 = n149;
  assign y5 = n155;
  assign y6 = n161;
  assign y7 = n167;
  assign y8 = n173;
  assign y9 = n179;
  assign y10 = n185;
  assign y11 = n191;
  assign y12 = n197;
  assign y13 = n203;
  assign y14 = n209;
  assign y15 = n215;
  assign y16 = n221;
  assign y17 = n226;
  assign y18 = n232;
  assign y19 = n237;
  assign y20 = n243;
  assign y21 = n249;
  assign y22 = n255;
  assign y23 = n261;
  assign y24 = n266;
  assign y25 = n271;
  assign y26 = n277;
  assign y27 = n283;
  assign y28 = n289;
  assign y29 = n295;
  assign y30 = n300;
  assign y31 = n306;
  assign y32 = n312;
  assign y33 = ~n318;
  assign y34 = n323;
  assign y35 = ~n329;
  assign y36 = ~n335;
  assign y37 = n340;
  assign y38 = ~n346;
  assign y39 = n352;
  assign y40 = n358;
  assign y41 = n363;
  assign y42 = n369;
  assign y43 = n374;
  assign y44 = n380;
  assign y45 = n385;
  assign y46 = n390;
  assign y47 = n396;
  assign y48 = n402;
  assign y49 = n407;
  assign y50 = n412;
  assign y51 = n417;
  assign y52 = n423;
  assign y53 = n428;
  assign y54 = n433;
  assign y55 = n438;
  assign y56 = n444;
  assign y57 = n449;
  assign y58 = n455;
  assign y59 = n460;
  assign y60 = ~n466;
  assign y61 = ~n472;
  assign y62 = ~n478;
  assign y63 = ~n484;
  assign y64 = ~n488;
endmodule
