module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700, x701, x702, x703, x704, x705, x706, x707, x708, x709, x710, x711, x712, x713, x714, x715, x716, x717, x718, x719, x720, x721, x722, x723, x724, x725, x726, x727, x728, x729, x730, x731, x732, x733, x734, x735, x736, x737, x738, x739, x740, x741, x742, x743, x744, x745, x746, x747, x748, x749, x750, x751, x752, x753, x754, x755, x756, x757, x758, x759, x760, x761, x762, x763, x764, x765, x766, x767, x768, x769, x770, x771, x772, x773, x774, x775, x776, x777, x778, x779, x780, x781, x782, x783, x784, x785, x786, x787, x788, x789, x790, x791, x792, x793, x794, x795, x796, x797, x798, x799, x800, x801, x802, x803, x804, x805, x806, x807, x808, x809, x810, x811, x812, x813, x814, x815, x816, x817, x818, x819, x820, x821, x822, x823, x824, x825, x826, x827, x828, x829, x830, x831, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700, x701, x702, x703, x704, x705, x706, x707, x708, x709, x710, x711, x712, x713, x714, x715, x716, x717, x718, x719, x720, x721, x722, x723, x724, x725, x726, x727, x728, x729, x730, x731, x732, x733, x734, x735, x736, x737, x738, x739, x740, x741, x742, x743, x744, x745, x746, x747, x748, x749, x750, x751, x752, x753, x754, x755, x756, x757, x758, x759, x760, x761, x762, x763, x764, x765, x766, x767, x768, x769, x770, x771, x772, x773, x774, x775, x776, x777, x778, x779, x780, x781, x782, x783, x784, x785, x786, x787, x788, x789, x790, x791, x792, x793, x794, x795, x796, x797, x798, x799, x800, x801, x802, x803, x804, x805, x806, x807, x808, x809, x810, x811, x812, x813, x814, x815, x816, x817, x818, x819, x820, x821, x822, x823, x824, x825, x826, x827, x828, x829, x830, x831;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63;
  wire n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403;
  assign n833 = x70 ^ x32;
  assign n834 = x75 ^ x58;
  assign n835 = n833 & n834;
  assign n836 = x74 ^ x0;
  assign n837 = x72 ^ x16;
  assign n838 = n836 & n837;
  assign n839 = x71 ^ x24;
  assign n840 = x73 ^ x8;
  assign n841 = ~n839 & n840;
  assign n842 = n838 & n841;
  assign n843 = n835 & n842;
  assign n844 = ~n833 & n834;
  assign n845 = n836 & ~n837;
  assign n846 = n839 & ~n840;
  assign n847 = n845 & n846;
  assign n848 = n839 & n840;
  assign n849 = ~n836 & ~n837;
  assign n850 = n848 & n849;
  assign n851 = ~n847 & ~n850;
  assign n852 = n844 & ~n851;
  assign n853 = ~n839 & ~n840;
  assign n854 = n838 & n853;
  assign n855 = n841 & n849;
  assign n856 = ~n854 & ~n855;
  assign n857 = n844 & ~n856;
  assign n858 = n842 ^ n833;
  assign n859 = n858 ^ n842;
  assign n860 = n845 & n848;
  assign n861 = ~n836 & n837;
  assign n862 = n848 & n861;
  assign n863 = ~n860 & ~n862;
  assign n864 = n863 ^ n842;
  assign n865 = n859 & ~n864;
  assign n866 = n865 ^ n842;
  assign n867 = ~n834 & n866;
  assign n868 = ~n857 & ~n867;
  assign n869 = ~n833 & ~n834;
  assign n870 = n841 & n861;
  assign n871 = n869 & n870;
  assign n872 = n833 & ~n834;
  assign n873 = n849 & n853;
  assign n874 = ~n842 & ~n873;
  assign n875 = n872 & ~n874;
  assign n876 = ~n871 & ~n875;
  assign n877 = n845 & n853;
  assign n878 = n869 & n877;
  assign n879 = n853 & n861;
  assign n880 = n841 & n845;
  assign n881 = ~n879 & ~n880;
  assign n882 = n835 & ~n881;
  assign n883 = ~n878 & ~n882;
  assign n884 = n846 & n861;
  assign n885 = n838 & n846;
  assign n886 = ~n884 & ~n885;
  assign n887 = n851 & ~n870;
  assign n888 = n886 & n887;
  assign n889 = n835 & ~n888;
  assign n890 = n840 ^ n836;
  assign n891 = n839 ^ n837;
  assign n892 = ~n890 & ~n891;
  assign n893 = n844 & n892;
  assign n894 = ~n889 & ~n893;
  assign n895 = n846 & n849;
  assign n896 = n856 & ~n895;
  assign n897 = ~n885 & n896;
  assign n898 = n872 & ~n897;
  assign n899 = n851 & ~n862;
  assign n900 = ~n885 & n899;
  assign n901 = n900 ^ n879;
  assign n902 = n879 ^ n869;
  assign n903 = ~n879 & ~n902;
  assign n904 = n903 ^ n879;
  assign n905 = ~n901 & ~n904;
  assign n906 = n905 ^ n903;
  assign n907 = n906 ^ n879;
  assign n908 = n907 ^ n869;
  assign n909 = ~n898 & ~n908;
  assign n910 = n909 ^ n898;
  assign n911 = n894 & ~n910;
  assign n912 = n883 & n911;
  assign n913 = n876 & n912;
  assign n914 = n868 & n913;
  assign n915 = ~n852 & n914;
  assign n916 = ~n843 & n915;
  assign n917 = n916 ^ x27;
  assign n918 = n917 ^ x129;
  assign n919 = x93 ^ x28;
  assign n920 = x88 ^ x2;
  assign n921 = n919 & n920;
  assign n922 = x90 ^ x52;
  assign n923 = x91 ^ x44;
  assign n924 = n922 & n923;
  assign n925 = x89 ^ x60;
  assign n926 = x92 ^ x36;
  assign n927 = ~n925 & n926;
  assign n928 = n924 & n927;
  assign n929 = n921 & n928;
  assign n930 = n919 & ~n920;
  assign n931 = n925 & ~n926;
  assign n932 = n924 & n931;
  assign n933 = n922 & ~n923;
  assign n934 = n925 & n926;
  assign n935 = n933 & n934;
  assign n936 = ~n932 & ~n935;
  assign n937 = n930 & ~n936;
  assign n938 = ~n929 & ~n937;
  assign n939 = ~n922 & ~n923;
  assign n940 = ~n925 & ~n926;
  assign n941 = n939 & n940;
  assign n942 = n921 & n941;
  assign n943 = n924 & n940;
  assign n944 = n927 & n939;
  assign n945 = ~n943 & ~n944;
  assign n946 = n930 & ~n945;
  assign n947 = ~n942 & ~n946;
  assign n948 = ~n922 & n923;
  assign n949 = n927 & n948;
  assign n950 = n931 & n948;
  assign n951 = n934 & n948;
  assign n952 = ~n950 & ~n951;
  assign n953 = ~n949 & n952;
  assign n954 = n930 & ~n953;
  assign n955 = ~n919 & ~n920;
  assign n956 = n931 & n939;
  assign n957 = ~n943 & ~n956;
  assign n958 = n931 & n933;
  assign n959 = n924 & n934;
  assign n960 = ~n958 & ~n959;
  assign n961 = n957 & n960;
  assign n962 = n955 & ~n961;
  assign n963 = ~n954 & ~n962;
  assign n964 = n934 & n939;
  assign n965 = ~n919 & n920;
  assign n966 = ~n951 & ~n958;
  assign n967 = ~n965 & n966;
  assign n968 = ~n964 & n967;
  assign n969 = ~n928 & ~n964;
  assign n970 = n933 & n940;
  assign n971 = ~n949 & ~n970;
  assign n972 = n927 & n933;
  assign n973 = ~n950 & ~n972;
  assign n974 = ~n959 & n973;
  assign n975 = n971 & n974;
  assign n976 = n921 & ~n966;
  assign n977 = n975 & ~n976;
  assign n978 = n969 & n977;
  assign n979 = ~n956 & n978;
  assign n980 = ~n968 & ~n979;
  assign n981 = n920 & n980;
  assign n982 = n963 & ~n981;
  assign n983 = ~n944 & ~n972;
  assign n984 = n983 ^ n921;
  assign n985 = n983 ^ n955;
  assign n986 = n985 ^ n955;
  assign n987 = n940 & n948;
  assign n988 = n987 ^ n955;
  assign n989 = n986 & ~n988;
  assign n990 = n989 ^ n955;
  assign n991 = ~n984 & n990;
  assign n992 = n991 ^ n921;
  assign n993 = n982 & ~n992;
  assign n994 = n947 & n993;
  assign n995 = n938 & n994;
  assign n996 = n941 ^ n919;
  assign n997 = n996 ^ n941;
  assign n998 = ~n932 & ~n951;
  assign n999 = n998 ^ n941;
  assign n1000 = ~n997 & ~n999;
  assign n1001 = n1000 ^ n941;
  assign n1002 = ~n920 & n1001;
  assign n1003 = n995 & ~n1002;
  assign n1004 = n1003 ^ x1;
  assign n1005 = n1004 ^ x124;
  assign n1006 = ~n918 & n1005;
  assign n1007 = x82 ^ x34;
  assign n1008 = x87 ^ x60;
  assign n1009 = ~n1007 & ~n1008;
  assign n1010 = x85 ^ x10;
  assign n1012 = x84 ^ x18;
  assign n1011 = x86 ^ x2;
  assign n1013 = n1012 ^ n1011;
  assign n1014 = n1013 ^ n1011;
  assign n1015 = x83 ^ x26;
  assign n1016 = n1015 ^ n1012;
  assign n1017 = n1016 ^ n1011;
  assign n1018 = n1017 ^ n1011;
  assign n1019 = n1018 ^ n1011;
  assign n1020 = n1014 & ~n1019;
  assign n1021 = n1020 ^ n1011;
  assign n1022 = n1010 & n1021;
  assign n1023 = n1022 ^ n1017;
  assign n1024 = n1009 & ~n1023;
  assign n1025 = n1010 & n1012;
  assign n1026 = n1015 & n1025;
  assign n1027 = ~n1011 & n1026;
  assign n1028 = ~n1010 & n1012;
  assign n1029 = ~n1011 & ~n1015;
  assign n1030 = n1028 & n1029;
  assign n1031 = ~n1027 & ~n1030;
  assign n1032 = n1008 & ~n1031;
  assign n1033 = n1007 & n1008;
  assign n1034 = ~n1010 & ~n1012;
  assign n1035 = ~n1015 & n1034;
  assign n1036 = n1011 & n1015;
  assign n1037 = n1012 & n1036;
  assign n1038 = n1010 & ~n1012;
  assign n1039 = n1011 & n1038;
  assign n1040 = ~n1037 & ~n1039;
  assign n1041 = ~n1035 & n1040;
  assign n1042 = n1033 & ~n1041;
  assign n1043 = ~n1032 & ~n1042;
  assign n1044 = ~n1024 & n1043;
  assign n1045 = ~n1007 & n1008;
  assign n1046 = n1011 & n1028;
  assign n1047 = ~n1011 & n1038;
  assign n1048 = n1011 & n1025;
  assign n1049 = ~n1015 & n1048;
  assign n1050 = n1034 & n1036;
  assign n1051 = ~n1049 & ~n1050;
  assign n1052 = ~n1047 & n1051;
  assign n1053 = ~n1046 & n1052;
  assign n1054 = n1045 & ~n1053;
  assign n1055 = n1007 & ~n1008;
  assign n1056 = ~n1011 & n1028;
  assign n1057 = n1038 ^ n1015;
  assign n1058 = n1057 ^ n1038;
  assign n1059 = n1011 & n1034;
  assign n1060 = ~n1025 & ~n1059;
  assign n1061 = n1060 ^ n1038;
  assign n1062 = n1058 & ~n1061;
  assign n1063 = n1062 ^ n1038;
  assign n1064 = ~n1056 & ~n1063;
  assign n1065 = ~n1048 & n1064;
  assign n1066 = n1055 & n1065;
  assign n1067 = ~n1054 & ~n1066;
  assign n1068 = n1044 & n1067;
  assign n1069 = n1068 ^ x51;
  assign n1070 = n1069 ^ x126;
  assign n1071 = x67 ^ x40;
  assign n1072 = x66 ^ x48;
  assign n1073 = n1071 & n1072;
  assign n1074 = x65 ^ x56;
  assign n1075 = x68 ^ x32;
  assign n1076 = n1074 & ~n1075;
  assign n1077 = n1073 & n1076;
  assign n1078 = x69 ^ x24;
  assign n1079 = x64 ^ x6;
  assign n1080 = n1078 & n1079;
  assign n1081 = n1071 & ~n1072;
  assign n1082 = n1076 & n1081;
  assign n1083 = n1080 & n1082;
  assign n1084 = n1078 & ~n1079;
  assign n1085 = ~n1074 & n1075;
  assign n1086 = n1073 & n1085;
  assign n1087 = n1084 & n1086;
  assign n1088 = ~n1083 & ~n1087;
  assign n1089 = n1074 & n1075;
  assign n1090 = ~n1071 & n1072;
  assign n1091 = n1089 & n1090;
  assign n1092 = n1080 & n1091;
  assign n1093 = ~n1071 & ~n1072;
  assign n1094 = n1076 & n1093;
  assign n1095 = n1080 & n1094;
  assign n1096 = ~n1074 & ~n1075;
  assign n1097 = n1093 & n1096;
  assign n1098 = n1089 & n1093;
  assign n1099 = n1081 & n1085;
  assign n1100 = n1081 & n1096;
  assign n1101 = n1085 & n1090;
  assign n1102 = ~n1100 & ~n1101;
  assign n1103 = ~n1099 & n1102;
  assign n1104 = ~n1098 & n1103;
  assign n1105 = ~n1091 & n1104;
  assign n1106 = ~n1097 & n1105;
  assign n1107 = n1084 & ~n1106;
  assign n1108 = ~n1078 & ~n1079;
  assign n1109 = n1076 & n1090;
  assign n1110 = n1073 & n1089;
  assign n1111 = ~n1082 & ~n1110;
  assign n1112 = ~n1109 & n1111;
  assign n1113 = n1108 & ~n1112;
  assign n1114 = n1094 & n1108;
  assign n1115 = n1099 & n1108;
  assign n1116 = n1090 & n1096;
  assign n1117 = n1073 & n1096;
  assign n1118 = ~n1086 & ~n1099;
  assign n1119 = ~n1117 & n1118;
  assign n1120 = ~n1116 & n1119;
  assign n1121 = n1080 & ~n1120;
  assign n1122 = n1085 & n1093;
  assign n1123 = ~n1116 & ~n1122;
  assign n1124 = n1108 & ~n1123;
  assign n1125 = ~n1078 & n1079;
  assign n1126 = n1074 ^ n1071;
  assign n1127 = n1126 ^ n1072;
  assign n1128 = n1126 ^ n1071;
  assign n1129 = ~n1127 & ~n1128;
  assign n1130 = n1129 ^ n1126;
  assign n1131 = ~n1075 & ~n1130;
  assign n1132 = n1131 ^ n1126;
  assign n1133 = ~n1109 & n1132;
  assign n1134 = n1125 & ~n1133;
  assign n1135 = ~n1124 & ~n1134;
  assign n1136 = ~n1121 & n1135;
  assign n1137 = ~n1115 & n1136;
  assign n1138 = ~n1114 & n1137;
  assign n1139 = ~n1113 & n1138;
  assign n1140 = ~n1107 & n1139;
  assign n1141 = ~n1095 & n1140;
  assign n1142 = ~n1092 & n1141;
  assign n1143 = n1088 & n1142;
  assign n1144 = ~n1077 & n1143;
  assign n1145 = n1144 ^ x59;
  assign n1146 = n1145 ^ x125;
  assign n1147 = n1070 & n1146;
  assign n1148 = x100 ^ x4;
  assign n1149 = x105 ^ x30;
  assign n1150 = n1148 & n1149;
  assign n1151 = x101 ^ x62;
  assign n1152 = x103 ^ x46;
  assign n1153 = ~n1151 & ~n1152;
  assign n1154 = x102 ^ x54;
  assign n1155 = x104 ^ x38;
  assign n1156 = ~n1154 & n1155;
  assign n1157 = n1153 & n1156;
  assign n1158 = n1150 & n1157;
  assign n1159 = ~n1148 & n1149;
  assign n1160 = ~n1151 & n1152;
  assign n1161 = ~n1154 & ~n1155;
  assign n1162 = n1160 & n1161;
  assign n1163 = n1159 & n1162;
  assign n1164 = ~n1158 & ~n1163;
  assign n1165 = n1151 & ~n1152;
  assign n1166 = n1156 & n1165;
  assign n1167 = n1154 & ~n1155;
  assign n1168 = n1165 & n1167;
  assign n1169 = ~n1166 & ~n1168;
  assign n1170 = n1159 & ~n1169;
  assign n1171 = n1151 & n1152;
  assign n1172 = ~n1155 & n1171;
  assign n1173 = n1150 & n1172;
  assign n1174 = n1160 & n1167;
  assign n1175 = ~n1157 & ~n1174;
  assign n1176 = n1159 & ~n1175;
  assign n1177 = ~n1173 & ~n1176;
  assign n1178 = ~n1170 & n1177;
  assign n1179 = n1154 & n1155;
  assign n1180 = n1153 & n1179;
  assign n1181 = n1159 & n1180;
  assign n1182 = n1161 & n1165;
  assign n1183 = ~n1148 & ~n1149;
  assign n1184 = ~n1150 & ~n1183;
  assign n1185 = n1182 & ~n1184;
  assign n1186 = ~n1181 & ~n1185;
  assign n1187 = n1165 & n1179;
  assign n1188 = n1150 & n1187;
  assign n1189 = n1159 & n1171;
  assign n1190 = n1167 & n1189;
  assign n1191 = n1160 & n1179;
  assign n1192 = n1159 & n1191;
  assign n1193 = ~n1190 & ~n1192;
  assign n1194 = n1148 & ~n1149;
  assign n1195 = n1154 ^ n1152;
  assign n1196 = n1155 ^ n1152;
  assign n1197 = n1196 ^ n1155;
  assign n1198 = n1154 ^ n1151;
  assign n1199 = n1198 ^ n1155;
  assign n1200 = n1199 ^ n1155;
  assign n1201 = n1200 ^ n1155;
  assign n1202 = ~n1197 & n1201;
  assign n1203 = n1202 ^ n1155;
  assign n1204 = ~n1195 & n1203;
  assign n1205 = n1204 ^ n1199;
  assign n1206 = n1194 & ~n1205;
  assign n1207 = n1156 & n1160;
  assign n1208 = n1153 & n1167;
  assign n1209 = ~n1207 & ~n1208;
  assign n1210 = ~n1174 & n1209;
  assign n1211 = n1150 & ~n1210;
  assign n1212 = ~n1162 & ~n1180;
  assign n1213 = ~n1156 & ~n1167;
  assign n1214 = n1171 & n1213;
  assign n1215 = n1175 & ~n1214;
  assign n1216 = ~n1187 & n1215;
  assign n1217 = n1212 & n1216;
  assign n1218 = n1183 & ~n1217;
  assign n1219 = ~n1211 & ~n1218;
  assign n1220 = ~n1206 & n1219;
  assign n1221 = n1193 & n1220;
  assign n1222 = ~n1188 & n1221;
  assign n1223 = n1186 & n1222;
  assign n1224 = n1178 & n1223;
  assign n1225 = n1164 & n1224;
  assign n1226 = n1225 ^ x35;
  assign n1227 = n1226 ^ x128;
  assign n1228 = x99 ^ x62;
  assign n1229 = x94 ^ x36;
  assign n1230 = n1228 & ~n1229;
  assign n1231 = x96 ^ x20;
  assign n1232 = x95 ^ x28;
  assign n1233 = ~n1231 & ~n1232;
  assign n1234 = x98 ^ x4;
  assign n1235 = x97 ^ x12;
  assign n1236 = n1234 & ~n1235;
  assign n1237 = n1233 & n1236;
  assign n1238 = ~n1234 & ~n1235;
  assign n1239 = n1231 & ~n1232;
  assign n1240 = n1238 & n1239;
  assign n1241 = ~n1237 & ~n1240;
  assign n1242 = n1231 & n1232;
  assign n1243 = ~n1234 & n1235;
  assign n1244 = n1242 & n1243;
  assign n1245 = n1232 & n1236;
  assign n1246 = n1231 & n1245;
  assign n1247 = ~n1244 & ~n1246;
  assign n1248 = n1241 & n1247;
  assign n1249 = n1230 & ~n1248;
  assign n1250 = ~n1228 & ~n1229;
  assign n1251 = n1236 & n1239;
  assign n1252 = n1250 & n1251;
  assign n1253 = n1233 & n1238;
  assign n1254 = n1230 & n1253;
  assign n1255 = ~n1252 & ~n1254;
  assign n1256 = n1234 & n1235;
  assign n1257 = n1233 & n1256;
  assign n1258 = ~n1229 & n1257;
  assign n1259 = n1239 & n1243;
  assign n1260 = n1228 & n1229;
  assign n1261 = ~n1250 & ~n1260;
  assign n1262 = n1259 & ~n1261;
  assign n1263 = ~n1258 & ~n1262;
  assign n1264 = n1237 & n1260;
  assign n1265 = ~n1231 & n1232;
  assign n1266 = n1238 & n1265;
  assign n1267 = n1256 & n1265;
  assign n1268 = ~n1266 & ~n1267;
  assign n1269 = n1230 & ~n1268;
  assign n1270 = n1238 & n1242;
  assign n1271 = ~n1231 & n1245;
  assign n1272 = ~n1270 & ~n1271;
  assign n1273 = n1268 & n1272;
  assign n1274 = n1260 & ~n1273;
  assign n1275 = n1242 & n1256;
  assign n1276 = ~n1228 & n1229;
  assign n1277 = ~n1275 & ~n1276;
  assign n1278 = n1243 & n1265;
  assign n1279 = ~n1246 & ~n1270;
  assign n1280 = ~n1278 & n1279;
  assign n1281 = n1277 & n1280;
  assign n1282 = ~n1228 & ~n1281;
  assign n1283 = ~n1274 & ~n1282;
  assign n1284 = n1233 & n1243;
  assign n1285 = n1239 & n1256;
  assign n1286 = ~n1284 & ~n1285;
  assign n1287 = ~n1250 & n1268;
  assign n1288 = n1260 & ~n1272;
  assign n1289 = n1287 & ~n1288;
  assign n1290 = n1241 & n1289;
  assign n1291 = n1286 & n1290;
  assign n1292 = ~n1275 & n1291;
  assign n1293 = ~n1244 & n1292;
  assign n1294 = ~n1283 & ~n1293;
  assign n1295 = ~n1269 & ~n1294;
  assign n1296 = ~n1264 & n1295;
  assign n1297 = n1263 & n1296;
  assign n1298 = n1284 ^ n1260;
  assign n1299 = n1260 ^ n1250;
  assign n1300 = n1299 ^ n1250;
  assign n1301 = n1285 ^ n1250;
  assign n1302 = n1300 & ~n1301;
  assign n1303 = n1302 ^ n1250;
  assign n1304 = n1298 & ~n1303;
  assign n1305 = n1304 ^ n1284;
  assign n1306 = n1297 & ~n1305;
  assign n1307 = n1255 & n1306;
  assign n1308 = ~n1249 & n1307;
  assign n1309 = n1308 ^ x43;
  assign n1310 = n1309 ^ x127;
  assign n1311 = n1227 & n1310;
  assign n1312 = n1147 & n1311;
  assign n1313 = n1006 & n1312;
  assign n1314 = n1070 & ~n1146;
  assign n1315 = ~n1227 & n1310;
  assign n1316 = n1314 & n1315;
  assign n1317 = n918 & n1005;
  assign n1318 = ~n918 & ~n1005;
  assign n1319 = ~n1317 & ~n1318;
  assign n1320 = n1316 & ~n1319;
  assign n1321 = n918 & ~n1005;
  assign n1322 = ~n1070 & n1146;
  assign n1323 = n1311 & n1322;
  assign n1324 = n1321 & n1323;
  assign n1325 = n1005 ^ n918;
  assign n1326 = n1311 & n1314;
  assign n1327 = n1326 ^ n1005;
  assign n1328 = n1327 ^ n1326;
  assign n1329 = n1227 & ~n1310;
  assign n1330 = n1322 & n1329;
  assign n1331 = n1330 ^ n1326;
  assign n1332 = ~n1328 & n1331;
  assign n1333 = n1332 ^ n1326;
  assign n1334 = ~n1325 & n1333;
  assign n1335 = ~n1324 & ~n1334;
  assign n1336 = ~n1320 & n1335;
  assign n1337 = n1318 & n1326;
  assign n1338 = n1147 & n1329;
  assign n1339 = ~n1323 & ~n1338;
  assign n1340 = n1006 & ~n1339;
  assign n1341 = ~n1337 & ~n1340;
  assign n1342 = ~n1227 & ~n1310;
  assign n1343 = n1147 & n1342;
  assign n1344 = ~n1318 & n1343;
  assign n1345 = ~n1070 & ~n1146;
  assign n1346 = n1311 & n1345;
  assign n1347 = n1322 & n1342;
  assign n1348 = ~n1070 & n1315;
  assign n1349 = n1146 & n1348;
  assign n1350 = ~n1338 & ~n1349;
  assign n1351 = ~n1347 & n1350;
  assign n1352 = ~n1346 & n1351;
  assign n1353 = ~n1319 & ~n1352;
  assign n1354 = ~n1344 & ~n1353;
  assign n1355 = n1342 & n1345;
  assign n1356 = n1317 & n1355;
  assign n1357 = ~n1312 & ~n1330;
  assign n1358 = n1321 & ~n1357;
  assign n1359 = ~n1356 & ~n1358;
  assign n1360 = n1314 & n1342;
  assign n1361 = n1318 & n1360;
  assign n1362 = n1329 & n1345;
  assign n1363 = ~n1146 & n1348;
  assign n1364 = n1314 & n1329;
  assign n1365 = ~n1363 & ~n1364;
  assign n1366 = ~n1362 & n1365;
  assign n1367 = ~n1355 & n1366;
  assign n1368 = ~n1321 & n1367;
  assign n1369 = n1147 & n1315;
  assign n1370 = ~n1360 & ~n1362;
  assign n1371 = ~n1006 & n1370;
  assign n1372 = ~n1363 & n1371;
  assign n1373 = ~n1369 & n1372;
  assign n1374 = ~n1368 & ~n1373;
  assign n1375 = n1319 & n1374;
  assign n1376 = ~n1361 & ~n1375;
  assign n1377 = n1359 & n1376;
  assign n1378 = n1354 & n1377;
  assign n1379 = n1341 & n1378;
  assign n1380 = n1336 & n1379;
  assign n1381 = ~n1313 & n1380;
  assign n1382 = n1381 ^ x2;
  assign n1383 = n1382 ^ x184;
  assign n1384 = n1009 & ~n1053;
  assign n1385 = n1033 & ~n1065;
  assign n1386 = ~n1384 & ~n1385;
  assign n1387 = n1008 ^ n1007;
  assign n1388 = n1041 ^ n1008;
  assign n1389 = n1388 ^ n1041;
  assign n1390 = n1041 ^ n1023;
  assign n1391 = n1389 & ~n1390;
  assign n1392 = n1391 ^ n1041;
  assign n1393 = n1387 & ~n1392;
  assign n1394 = n1386 & ~n1393;
  assign n1395 = n1031 & n1394;
  assign n1396 = n1395 ^ x57;
  assign n1397 = n1396 ^ x159;
  assign n1398 = n850 & n869;
  assign n1399 = n884 ^ n833;
  assign n1400 = n1399 ^ n884;
  assign n1401 = n884 ^ n870;
  assign n1402 = ~n1400 & n1401;
  assign n1403 = n1402 ^ n884;
  assign n1404 = n834 & n1403;
  assign n1405 = ~n1398 & ~n1404;
  assign n1406 = n838 & n848;
  assign n1407 = n834 ^ n833;
  assign n1408 = n1406 & ~n1407;
  assign n1409 = ~n855 & ~n895;
  assign n1410 = ~n877 & n1409;
  assign n1411 = n835 & ~n1410;
  assign n1412 = ~n1408 & ~n1411;
  assign n1413 = n869 & ~n897;
  assign n1414 = ~n854 & ~n873;
  assign n1415 = n863 & n1414;
  assign n1416 = ~n885 & n1415;
  assign n1417 = n844 & ~n1416;
  assign n1418 = ~n847 & n886;
  assign n1419 = ~n862 & n1418;
  assign n1420 = n881 & n1419;
  assign n1421 = n872 & ~n1420;
  assign n1422 = ~n1417 & ~n1421;
  assign n1423 = ~n1413 & n1422;
  assign n1424 = n1412 & n1423;
  assign n1425 = n883 & n1424;
  assign n1426 = n876 & n1425;
  assign n1427 = n1405 & n1426;
  assign n1428 = ~n852 & n1427;
  assign n1429 = ~n843 & n1428;
  assign n1430 = n1429 ^ x39;
  assign n1431 = n1430 ^ x154;
  assign n1432 = ~n1397 & n1431;
  assign n1433 = x78 ^ x50;
  assign n1434 = x80 ^ x34;
  assign n1435 = ~n1433 & ~n1434;
  assign n1436 = x79 ^ x42;
  assign n1437 = x77 ^ x58;
  assign n1438 = n1436 & ~n1437;
  assign n1439 = n1435 & n1438;
  assign n1440 = ~n1436 & n1437;
  assign n1441 = n1435 & n1440;
  assign n1442 = x81 ^ x26;
  assign n1443 = x76 ^ x0;
  assign n1444 = n1442 & ~n1443;
  assign n1445 = ~n1442 & n1443;
  assign n1446 = ~n1444 & ~n1445;
  assign n1447 = n1441 & n1446;
  assign n1448 = n1433 & n1434;
  assign n1450 = ~n1436 & ~n1437;
  assign n1451 = n1448 & n1450;
  assign n1449 = n1440 & n1448;
  assign n1452 = n1451 ^ n1449;
  assign n1453 = n1452 ^ n1451;
  assign n1454 = n1451 ^ n1445;
  assign n1455 = n1454 ^ n1451;
  assign n1456 = n1453 & ~n1455;
  assign n1457 = n1456 ^ n1451;
  assign n1458 = ~n1444 & n1457;
  assign n1459 = n1458 ^ n1451;
  assign n1460 = ~n1447 & ~n1459;
  assign n1461 = n1442 & n1443;
  assign n1462 = ~n1433 & n1434;
  assign n1463 = n1438 & n1462;
  assign n1464 = n1435 & n1450;
  assign n1465 = ~n1463 & ~n1464;
  assign n1466 = n1461 & ~n1465;
  assign n1467 = n1436 & n1437;
  assign n1468 = n1448 & n1467;
  assign n1469 = n1435 & n1467;
  assign n1470 = ~n1468 & ~n1469;
  assign n1471 = n1444 & ~n1470;
  assign n1472 = ~n1466 & ~n1471;
  assign n1473 = ~n1446 & ~n1465;
  assign n1474 = n1433 & ~n1434;
  assign n1475 = n1450 & n1474;
  assign n1476 = n1445 & n1475;
  assign n1477 = n1440 & n1462;
  assign n1478 = n1440 & n1474;
  assign n1479 = ~n1477 & ~n1478;
  assign n1480 = n1444 & ~n1479;
  assign n1481 = ~n1476 & ~n1480;
  assign n1482 = ~n1442 & ~n1443;
  assign n1483 = n1450 & n1462;
  assign n1484 = n1438 & n1448;
  assign n1485 = ~n1477 & ~n1484;
  assign n1486 = ~n1483 & n1485;
  assign n1487 = n1470 & n1486;
  assign n1488 = n1482 & ~n1487;
  assign n1489 = n1438 & n1474;
  assign n1490 = ~n1451 & ~n1489;
  assign n1491 = ~n1439 & n1490;
  assign n1492 = ~n1468 & n1491;
  assign n1493 = n1461 & ~n1492;
  assign n1494 = n1462 & n1467;
  assign n1495 = n1479 & ~n1494;
  assign n1496 = ~n1484 & n1495;
  assign n1497 = n1445 & ~n1496;
  assign n1498 = ~n1493 & ~n1497;
  assign n1499 = ~n1488 & n1498;
  assign n1500 = n1481 & n1499;
  assign n1501 = ~n1473 & n1500;
  assign n1502 = n1472 & n1501;
  assign n1503 = n1460 & n1502;
  assign n1504 = ~n1439 & n1503;
  assign n1505 = n1504 ^ x23;
  assign n1506 = n1505 ^ x156;
  assign n1507 = ~n1097 & ~n1101;
  assign n1508 = n1080 & ~n1507;
  assign n1509 = ~n1102 & n1108;
  assign n1510 = ~n1508 & ~n1509;
  assign n1511 = n1081 & n1089;
  assign n1512 = ~n1077 & ~n1511;
  assign n1513 = ~n1091 & ~n1109;
  assign n1514 = n1512 & n1513;
  assign n1515 = n1514 ^ n1086;
  assign n1516 = n1515 ^ n1086;
  assign n1517 = n1086 ^ n1078;
  assign n1518 = n1517 ^ n1086;
  assign n1519 = ~n1516 & n1518;
  assign n1520 = n1519 ^ n1086;
  assign n1521 = ~n1079 & n1520;
  assign n1522 = n1521 ^ n1086;
  assign n1523 = n1510 & ~n1522;
  assign n1524 = ~n1080 & ~n1108;
  assign n1525 = n1117 & ~n1524;
  assign n1526 = ~n1094 & n1123;
  assign n1527 = n1125 & ~n1526;
  assign n1528 = n1108 & ~n1513;
  assign n1529 = ~n1095 & ~n1528;
  assign n1530 = ~n1100 & ~n1122;
  assign n1531 = ~n1117 & n1530;
  assign n1532 = n1084 & ~n1531;
  assign n1533 = ~n1109 & n1512;
  assign n1534 = ~n1082 & n1533;
  assign n1535 = n1125 & ~n1534;
  assign n1536 = ~n1532 & ~n1535;
  assign n1537 = n1110 ^ n1080;
  assign n1538 = n1110 ^ n1108;
  assign n1539 = n1538 ^ n1108;
  assign n1540 = n1108 ^ n1098;
  assign n1541 = ~n1539 & ~n1540;
  assign n1542 = n1541 ^ n1108;
  assign n1543 = n1537 & n1542;
  assign n1544 = n1543 ^ n1080;
  assign n1545 = n1536 & ~n1544;
  assign n1546 = n1529 & n1545;
  assign n1547 = ~n1114 & n1546;
  assign n1548 = n1088 & n1547;
  assign n1549 = ~n1527 & n1548;
  assign n1550 = ~n1525 & n1549;
  assign n1551 = n1523 & n1550;
  assign n1552 = ~n1115 & n1551;
  assign n1553 = n1552 ^ x15;
  assign n1554 = n1553 ^ x157;
  assign n1555 = ~n1506 & n1554;
  assign n1556 = n1159 & n1207;
  assign n1557 = n1179 & n1189;
  assign n1558 = ~n1188 & ~n1557;
  assign n1559 = ~n1166 & ~n1191;
  assign n1560 = n1150 & ~n1559;
  assign n1561 = n1150 & n1208;
  assign n1562 = n1161 & n1189;
  assign n1563 = ~n1561 & ~n1562;
  assign n1564 = n1159 & n1208;
  assign n1565 = n1183 & ~n1205;
  assign n1566 = ~n1564 & ~n1565;
  assign n1567 = n1153 & n1161;
  assign n1568 = ~n1180 & ~n1567;
  assign n1569 = n1148 & ~n1568;
  assign n1570 = ~n1168 & n1216;
  assign n1571 = n1194 & ~n1570;
  assign n1572 = ~n1569 & ~n1571;
  assign n1573 = n1566 & n1572;
  assign n1574 = n1563 & n1573;
  assign n1575 = ~n1560 & n1574;
  assign n1576 = n1558 & n1575;
  assign n1577 = n1178 & n1576;
  assign n1578 = ~n1556 & n1577;
  assign n1579 = n1578 ^ x7;
  assign n1580 = n1579 ^ x158;
  assign n1581 = n1230 & n1259;
  assign n1582 = ~n1241 & ~n1261;
  assign n1583 = ~n1581 & ~n1582;
  assign n1584 = ~n1257 & ~n1275;
  assign n1585 = n1272 & n1584;
  assign n1586 = n1247 & n1585;
  assign n1587 = n1230 & ~n1586;
  assign n1588 = ~n1278 & ~n1285;
  assign n1589 = ~n1266 & n1588;
  assign n1590 = n1277 & n1589;
  assign n1591 = ~n1260 & n1590;
  assign n1592 = n1247 & ~n1278;
  assign n1593 = ~n1266 & n1592;
  assign n1594 = n1593 ^ n1228;
  assign n1595 = n1594 ^ n1593;
  assign n1596 = n1234 ^ n1231;
  assign n1597 = n1596 ^ n1232;
  assign n1598 = n1597 ^ n1235;
  assign n1599 = ~n1232 & n1598;
  assign n1600 = ~n1234 & n1599;
  assign n1601 = n1600 ^ n1597;
  assign n1602 = n1601 ^ n1593;
  assign n1603 = ~n1595 & ~n1602;
  assign n1604 = n1603 ^ n1593;
  assign n1605 = n1229 & ~n1604;
  assign n1606 = n1605 ^ n1228;
  assign n1607 = ~n1591 & ~n1606;
  assign n1608 = ~n1587 & ~n1607;
  assign n1609 = n1583 & n1608;
  assign n1610 = ~n1305 & n1609;
  assign n1611 = n1255 & n1610;
  assign n1612 = n1611 ^ x31;
  assign n1613 = n1612 ^ x155;
  assign n1614 = n1580 & n1613;
  assign n1615 = n1555 & n1614;
  assign n1616 = n1432 & n1615;
  assign n1617 = n1397 & ~n1431;
  assign n1618 = n1506 & n1554;
  assign n1619 = n1614 & n1618;
  assign n1620 = ~n1506 & ~n1554;
  assign n1621 = ~n1580 & n1613;
  assign n1622 = n1620 & n1621;
  assign n1623 = ~n1619 & ~n1622;
  assign n1624 = n1617 & ~n1623;
  assign n1625 = n1397 & n1431;
  assign n1626 = n1580 & ~n1613;
  assign n1627 = n1618 & n1626;
  assign n1628 = ~n1580 & ~n1613;
  assign n1629 = n1555 & n1628;
  assign n1630 = ~n1627 & ~n1629;
  assign n1631 = n1625 & ~n1630;
  assign n1632 = ~n1624 & ~n1631;
  assign n1633 = ~n1613 & n1620;
  assign n1634 = ~n1580 & n1633;
  assign n1635 = n1432 & n1634;
  assign n1636 = n1614 & n1620;
  assign n1637 = n1625 & n1636;
  assign n1638 = n1555 & n1621;
  assign n1639 = n1432 & n1638;
  assign n1640 = ~n1637 & ~n1639;
  assign n1641 = ~n1635 & n1640;
  assign n1642 = ~n1397 & ~n1431;
  assign n1643 = n1638 & n1642;
  assign n1644 = n1618 & n1628;
  assign n1645 = n1617 & n1644;
  assign n1646 = ~n1643 & ~n1645;
  assign n1647 = n1506 & ~n1554;
  assign n1648 = n1614 & n1647;
  assign n1649 = ~n1622 & ~n1648;
  assign n1650 = n1432 & ~n1649;
  assign n1651 = n1618 & n1621;
  assign n1652 = ~n1648 & ~n1651;
  assign n1653 = n1617 & ~n1652;
  assign n1654 = ~n1650 & ~n1653;
  assign n1655 = ~n1619 & ~n1636;
  assign n1656 = n1642 & ~n1655;
  assign n1657 = n1628 & n1647;
  assign n1658 = n1626 & n1647;
  assign n1659 = ~n1627 & ~n1658;
  assign n1660 = ~n1657 & n1659;
  assign n1661 = n1432 & ~n1660;
  assign n1662 = ~n1656 & ~n1661;
  assign n1663 = n1431 ^ n1397;
  assign n1664 = n1621 & n1647;
  assign n1665 = ~n1663 & n1664;
  assign n1666 = ~n1615 & ~n1657;
  assign n1667 = n1625 & ~n1666;
  assign n1668 = n1580 & n1633;
  assign n1669 = ~n1658 & ~n1668;
  assign n1670 = ~n1638 & n1669;
  assign n1671 = n1617 & ~n1670;
  assign n1672 = ~n1628 & ~n1642;
  assign n1673 = n1555 & n1626;
  assign n1674 = ~n1644 & ~n1673;
  assign n1675 = ~n1633 & n1674;
  assign n1676 = ~n1672 & ~n1675;
  assign n1677 = ~n1663 & n1676;
  assign n1678 = ~n1671 & ~n1677;
  assign n1679 = ~n1667 & n1678;
  assign n1680 = ~n1665 & n1679;
  assign n1681 = n1662 & n1680;
  assign n1682 = n1654 & n1681;
  assign n1683 = n1646 & n1682;
  assign n1684 = n1641 & n1683;
  assign n1685 = n1632 & n1684;
  assign n1686 = ~n1616 & n1685;
  assign n1687 = n1686 ^ x28;
  assign n1688 = n1687 ^ x189;
  assign n1689 = ~n1383 & n1688;
  assign n1690 = n1250 & n1259;
  assign n1691 = ~n1229 & n1266;
  assign n1692 = ~n1690 & ~n1691;
  assign n1693 = ~n1237 & ~n1251;
  assign n1694 = ~n1261 & ~n1693;
  assign n1695 = ~n1257 & n1286;
  assign n1696 = ~n1240 & ~n1244;
  assign n1697 = n1272 & n1696;
  assign n1698 = n1695 & n1697;
  assign n1699 = n1230 & ~n1698;
  assign n1700 = ~n1694 & ~n1699;
  assign n1701 = ~n1253 & ~n1284;
  assign n1702 = n1260 & ~n1701;
  assign n1703 = ~n1267 & n1280;
  assign n1704 = n1228 & n1703;
  assign n1705 = ~n1260 & n1592;
  assign n1706 = ~n1267 & n1705;
  assign n1707 = ~n1261 & ~n1706;
  assign n1708 = n1585 & n1589;
  assign n1709 = ~n1240 & n1708;
  assign n1710 = n1276 & ~n1709;
  assign n1711 = ~n1707 & ~n1710;
  assign n1712 = ~n1704 & ~n1711;
  assign n1713 = ~n1702 & ~n1712;
  assign n1714 = n1700 & n1713;
  assign n1715 = n1692 & n1714;
  assign n1716 = n1715 ^ x33;
  assign n1717 = n1716 ^ x118;
  assign n1718 = n1145 ^ x123;
  assign n1719 = ~n1717 & n1718;
  assign n1720 = n1444 & n1475;
  assign n1721 = n1446 & n1494;
  assign n1722 = ~n1720 & ~n1721;
  assign n1723 = n1445 & ~n1490;
  assign n1724 = ~n1473 & ~n1723;
  assign n1725 = n1443 ^ n1441;
  assign n1726 = n1725 ^ n1441;
  assign n1727 = n1449 ^ n1441;
  assign n1728 = n1727 ^ n1441;
  assign n1729 = n1726 & n1728;
  assign n1730 = n1729 ^ n1441;
  assign n1731 = n1442 & n1730;
  assign n1732 = n1731 ^ n1441;
  assign n1733 = n1724 & ~n1732;
  assign n1734 = n1482 & ~n1491;
  assign n1735 = n1484 ^ n1461;
  assign n1736 = n1484 ^ n1482;
  assign n1737 = n1736 ^ n1482;
  assign n1738 = ~n1451 & ~n1464;
  assign n1739 = ~n1439 & n1738;
  assign n1740 = n1739 ^ n1482;
  assign n1741 = ~n1737 & n1740;
  assign n1742 = n1741 ^ n1482;
  assign n1743 = n1735 & n1742;
  assign n1744 = n1743 ^ n1461;
  assign n1745 = ~n1734 & ~n1744;
  assign n1746 = n1479 ^ n1444;
  assign n1747 = n1746 ^ n1479;
  assign n1748 = n1467 & n1474;
  assign n1749 = ~n1449 & ~n1748;
  assign n1750 = n1470 & n1749;
  assign n1751 = n1750 ^ n1479;
  assign n1752 = n1747 & n1751;
  assign n1753 = n1752 ^ n1479;
  assign n1754 = n1745 & n1753;
  assign n1755 = n1733 & n1754;
  assign n1756 = n1443 ^ n1442;
  assign n1757 = n1468 ^ n1443;
  assign n1758 = n1757 ^ n1468;
  assign n1759 = n1483 ^ n1468;
  assign n1760 = ~n1758 & n1759;
  assign n1761 = n1760 ^ n1468;
  assign n1762 = n1756 & n1761;
  assign n1763 = n1755 & ~n1762;
  assign n1764 = n1722 & n1763;
  assign n1765 = n1764 ^ x17;
  assign n1766 = n1765 ^ x120;
  assign n1767 = x111 ^ x56;
  assign n1768 = x106 ^ x38;
  assign n1769 = n1767 & n1768;
  assign n1770 = x109 ^ x14;
  assign n1771 = x108 ^ x22;
  assign n1772 = ~n1770 & n1771;
  assign n1773 = x110 ^ x6;
  assign n1774 = x107 ^ x30;
  assign n1775 = ~n1773 & n1774;
  assign n1776 = n1772 & n1775;
  assign n1777 = n1769 & n1776;
  assign n1778 = ~n1767 & n1768;
  assign n1779 = ~n1770 & ~n1771;
  assign n1780 = n1775 & n1779;
  assign n1781 = n1773 & n1774;
  assign n1782 = n1772 & n1781;
  assign n1783 = ~n1780 & ~n1782;
  assign n1784 = n1778 & ~n1783;
  assign n1785 = ~n1767 & ~n1768;
  assign n1786 = n1770 & n1771;
  assign n1787 = n1781 & n1786;
  assign n1788 = n1770 & ~n1771;
  assign n1789 = n1775 & n1788;
  assign n1790 = ~n1787 & ~n1789;
  assign n1791 = ~n1776 & n1790;
  assign n1792 = n1785 & ~n1791;
  assign n1793 = ~n1784 & ~n1792;
  assign n1794 = n1767 & ~n1768;
  assign n1795 = n1773 & ~n1774;
  assign n1796 = n1786 & n1795;
  assign n1797 = ~n1773 & ~n1774;
  assign n1798 = n1779 & n1797;
  assign n1799 = ~n1796 & ~n1798;
  assign n1800 = n1772 & n1795;
  assign n1801 = n1786 & n1797;
  assign n1802 = ~n1800 & ~n1801;
  assign n1803 = n1799 & n1802;
  assign n1804 = n1794 & ~n1803;
  assign n1805 = n1788 & n1795;
  assign n1806 = n1769 & n1805;
  assign n1807 = ~n1790 & n1794;
  assign n1808 = ~n1806 & ~n1807;
  assign n1809 = ~n1778 & ~n1785;
  assign n1810 = ~n1796 & ~n1805;
  assign n1811 = ~n1809 & ~n1810;
  assign n1812 = n1779 & n1781;
  assign n1813 = ~n1776 & ~n1812;
  assign n1814 = n1794 & ~n1813;
  assign n1815 = ~n1811 & ~n1814;
  assign n1816 = ~n1769 & ~n1785;
  assign n1817 = n1779 & n1795;
  assign n1818 = n1772 & n1797;
  assign n1819 = ~n1817 & ~n1818;
  assign n1820 = ~n1816 & ~n1819;
  assign n1821 = n1798 ^ n1778;
  assign n1822 = n1798 ^ n1769;
  assign n1823 = n1822 ^ n1769;
  assign n1824 = n1788 & n1797;
  assign n1825 = n1775 & n1786;
  assign n1826 = ~n1824 & ~n1825;
  assign n1827 = ~n1812 & n1826;
  assign n1828 = n1827 ^ n1769;
  assign n1829 = ~n1823 & n1828;
  assign n1830 = n1829 ^ n1769;
  assign n1831 = n1821 & n1830;
  assign n1832 = n1831 ^ n1778;
  assign n1833 = ~n1820 & ~n1832;
  assign n1834 = n1815 & n1833;
  assign n1835 = n1808 & n1834;
  assign n1836 = ~n1804 & n1835;
  assign n1837 = n1793 & n1836;
  assign n1838 = n1782 ^ n1769;
  assign n1839 = n1785 ^ n1782;
  assign n1840 = n1839 ^ n1785;
  assign n1841 = n1781 & n1788;
  assign n1842 = ~n1825 & ~n1841;
  assign n1843 = n1842 ^ n1785;
  assign n1844 = ~n1840 & n1843;
  assign n1845 = n1844 ^ n1785;
  assign n1846 = n1838 & n1845;
  assign n1847 = n1846 ^ n1769;
  assign n1848 = n1837 & ~n1847;
  assign n1849 = ~n1777 & n1848;
  assign n1850 = n1849 ^ x25;
  assign n1851 = n1850 ^ x119;
  assign n1852 = n1766 & n1851;
  assign n1853 = n1004 ^ x122;
  assign n1854 = n1184 & n1567;
  assign n1855 = n1194 & n1207;
  assign n1856 = n1167 & n1171;
  assign n1857 = n1194 & n1856;
  assign n1858 = n1156 & n1171;
  assign n1859 = ~n1214 & ~n1858;
  assign n1860 = ~n1168 & n1859;
  assign n1861 = ~n1191 & n1860;
  assign n1862 = n1183 & ~n1861;
  assign n1863 = ~n1857 & ~n1862;
  assign n1864 = n1149 ^ n1148;
  assign n1867 = ~n1166 & ~n1174;
  assign n1868 = ~n1187 & n1867;
  assign n1865 = n1171 & ~n1213;
  assign n1866 = ~n1162 & ~n1865;
  assign n1869 = n1868 ^ n1866;
  assign n1870 = n1869 ^ n1868;
  assign n1871 = n1868 ^ n1149;
  assign n1872 = n1871 ^ n1868;
  assign n1873 = ~n1870 & n1872;
  assign n1874 = n1873 ^ n1868;
  assign n1875 = ~n1864 & ~n1874;
  assign n1876 = n1875 ^ n1868;
  assign n1877 = n1863 & n1876;
  assign n1878 = ~n1855 & n1877;
  assign n1879 = ~n1854 & n1878;
  assign n1880 = ~n1157 & ~n1208;
  assign n1881 = n1880 ^ n1148;
  assign n1882 = n1881 ^ n1880;
  assign n1883 = n1880 ^ n1212;
  assign n1884 = n1882 & n1883;
  assign n1885 = n1884 ^ n1880;
  assign n1886 = ~n1149 & ~n1885;
  assign n1887 = n1879 & ~n1886;
  assign n1888 = n1186 & n1887;
  assign n1889 = ~n1560 & n1888;
  assign n1890 = n1563 & n1889;
  assign n1891 = n1164 & n1890;
  assign n1892 = ~n1556 & n1891;
  assign n1893 = n1892 ^ x9;
  assign n1894 = n1893 ^ x121;
  assign n1895 = ~n1853 & ~n1894;
  assign n1896 = n1852 & n1895;
  assign n1897 = n1719 & n1896;
  assign n1898 = n1766 & ~n1851;
  assign n1899 = n1853 & ~n1894;
  assign n1900 = n1898 & n1899;
  assign n1901 = n1717 & n1718;
  assign n1902 = ~n1717 & ~n1718;
  assign n1903 = ~n1901 & ~n1902;
  assign n1904 = n1900 & ~n1903;
  assign n1905 = ~n1897 & ~n1904;
  assign n1906 = ~n1766 & n1851;
  assign n1907 = ~n1853 & n1894;
  assign n1908 = n1906 & n1907;
  assign n1909 = n1852 & n1899;
  assign n1910 = ~n1908 & ~n1909;
  assign n1911 = n1902 & ~n1910;
  assign n1912 = n1853 & n1894;
  assign n1913 = n1906 & n1912;
  assign n1914 = n1901 & n1913;
  assign n1915 = n1717 & ~n1718;
  assign n1916 = n1899 & n1906;
  assign n1917 = ~n1896 & ~n1916;
  assign n1918 = n1915 & ~n1917;
  assign n1919 = ~n1914 & ~n1918;
  assign n1920 = ~n1911 & n1919;
  assign n1921 = n1898 & n1907;
  assign n1922 = n1901 & n1921;
  assign n1923 = ~n1766 & ~n1851;
  assign n1924 = n1895 & n1923;
  assign n1925 = n1901 & n1924;
  assign n1926 = n1901 & ~n1917;
  assign n1927 = n1852 & n1907;
  assign n1928 = n1717 & n1927;
  assign n1929 = n1894 ^ n1851;
  assign n1930 = n1929 ^ n1766;
  assign n1931 = n1930 ^ n1929;
  assign n1932 = n1929 ^ n1894;
  assign n1933 = ~n1931 & ~n1932;
  assign n1934 = n1933 ^ n1929;
  assign n1935 = ~n1853 & ~n1934;
  assign n1936 = n1935 ^ n1929;
  assign n1937 = n1719 & ~n1936;
  assign n1938 = n1898 & n1912;
  assign n1939 = n1907 & n1923;
  assign n1940 = ~n1938 & ~n1939;
  assign n1941 = n1912 & n1923;
  assign n1942 = ~n1921 & ~n1941;
  assign n1943 = n1940 & n1942;
  assign n1944 = n1915 & ~n1943;
  assign n1945 = n1895 & n1906;
  assign n1946 = n1895 & n1898;
  assign n1947 = ~n1941 & ~n1946;
  assign n1948 = ~n1924 & n1947;
  assign n1949 = ~n1945 & n1948;
  assign n1950 = n1902 & ~n1949;
  assign n1951 = ~n1944 & ~n1950;
  assign n1952 = ~n1937 & n1951;
  assign n1953 = ~n1928 & n1952;
  assign n1954 = ~n1926 & n1953;
  assign n1955 = n1899 & n1923;
  assign n1956 = n1955 ^ n1927;
  assign n1957 = n1927 ^ n1717;
  assign n1958 = n1957 ^ n1927;
  assign n1959 = n1956 & n1958;
  assign n1960 = n1959 ^ n1927;
  assign n1961 = n1718 & n1960;
  assign n1962 = n1954 & ~n1961;
  assign n1963 = ~n1925 & n1962;
  assign n1964 = ~n1922 & n1963;
  assign n1965 = n1920 & n1964;
  assign n1966 = n1905 & n1965;
  assign n1967 = n1913 ^ n1717;
  assign n1968 = n1967 ^ n1913;
  assign n1969 = n1913 ^ n1909;
  assign n1970 = n1968 & n1969;
  assign n1971 = n1970 ^ n1913;
  assign n1972 = ~n1718 & n1971;
  assign n1973 = n1966 & ~n1972;
  assign n1974 = n1973 ^ x52;
  assign n1975 = n1974 ^ x186;
  assign n1976 = n1098 & ~n1524;
  assign n1977 = n1111 & n1513;
  assign n1978 = n1125 & ~n1977;
  assign n1979 = ~n1976 & ~n1978;
  assign n1980 = ~n1094 & n1507;
  assign n1981 = n1084 & ~n1980;
  assign n1982 = ~n1110 & n1533;
  assign n1983 = n1084 & ~n1982;
  assign n1984 = n1119 & ~n1122;
  assign n1985 = n1125 & ~n1984;
  assign n1986 = ~n1983 & ~n1985;
  assign n1987 = n1080 & ~n1102;
  assign n1988 = n1103 & ~n1117;
  assign n1989 = ~n1108 & n1988;
  assign n1990 = ~n1120 & ~n1989;
  assign n1991 = ~n1987 & ~n1990;
  assign n1992 = ~n1524 & ~n1991;
  assign n1993 = n1986 & ~n1992;
  assign n1994 = ~n1981 & n1993;
  assign n1995 = n1079 ^ n1078;
  assign n1996 = n1109 ^ n1079;
  assign n1997 = n1996 ^ n1109;
  assign n1998 = ~n1077 & ~n1091;
  assign n1999 = n1998 ^ n1109;
  assign n2000 = ~n1997 & ~n1999;
  assign n2001 = n2000 ^ n1109;
  assign n2002 = ~n1995 & n2001;
  assign n2003 = n1994 & ~n2002;
  assign n2004 = n1979 & n2003;
  assign n2005 = ~n1092 & n2004;
  assign n2006 = ~n1114 & n2005;
  assign n2007 = n1088 & n2006;
  assign n2008 = n2007 ^ x61;
  assign n2009 = n2008 ^ x135;
  assign n2048 = n921 & ~n936;
  assign n2049 = ~n941 & ~n972;
  assign n2050 = n965 & ~n2049;
  assign n2051 = ~n2048 & ~n2050;
  assign n2052 = ~n949 & ~n987;
  assign n2053 = ~n972 & n2052;
  assign n2054 = n921 & ~n2053;
  assign n2055 = ~n943 & n960;
  assign n2056 = n952 & n2055;
  assign n2057 = n965 & ~n2056;
  assign n2058 = ~n2054 & ~n2057;
  assign n2059 = n920 & n956;
  assign n2060 = ~n921 & ~n955;
  assign n2061 = n964 & ~n2060;
  assign n2062 = ~n2059 & ~n2061;
  assign n2063 = ~n928 & ~n958;
  assign n2064 = ~n944 & ~n970;
  assign n2065 = ~n987 & n2064;
  assign n2066 = n2063 & n2065;
  assign n2067 = n955 & ~n2066;
  assign n2068 = n957 & n975;
  assign n2069 = n930 & ~n2068;
  assign n2070 = ~n2067 & ~n2069;
  assign n2071 = n2062 & n2070;
  assign n2072 = n2058 & n2071;
  assign n2073 = n2051 & n2072;
  assign n2074 = ~n1002 & n2073;
  assign n2075 = ~n929 & n2074;
  assign n2076 = n2075 ^ x19;
  assign n2077 = n2076 ^ x132;
  assign n2010 = n1469 & n1482;
  assign n2011 = n1446 & n1477;
  assign n2012 = ~n2010 & ~n2011;
  assign n2013 = n1461 & ~n1470;
  assign n2014 = ~n1442 & n1494;
  assign n2015 = ~n1478 & ~n1748;
  assign n2016 = ~n1446 & ~n2015;
  assign n2017 = n1436 ^ n1433;
  assign n2018 = n2017 ^ n1437;
  assign n2019 = n1436 ^ n1434;
  assign n2020 = n1437 ^ n1436;
  assign n2021 = n2020 ^ n1436;
  assign n2022 = ~n2019 & ~n2021;
  assign n2023 = n2022 ^ n1436;
  assign n2024 = ~n2018 & n2023;
  assign n2025 = n1444 & n2024;
  assign n2026 = ~n2016 & ~n2025;
  assign n2027 = ~n1483 & n1739;
  assign n2028 = n1445 & ~n2027;
  assign n2029 = ~n1439 & ~n1441;
  assign n2030 = ~n1482 & n2029;
  assign n2031 = ~n1463 & ~n1489;
  assign n2032 = ~n1461 & n2031;
  assign n2033 = ~n2030 & ~n2032;
  assign n2034 = ~n1475 & ~n2033;
  assign n2035 = ~n1484 & n2034;
  assign n2036 = n1446 & ~n2035;
  assign n2037 = ~n2028 & ~n2036;
  assign n2038 = n2026 & n2037;
  assign n2039 = ~n2014 & n2038;
  assign n2040 = ~n2013 & n2039;
  assign n2041 = n2012 & n2040;
  assign n2042 = ~n1459 & n2041;
  assign n2043 = ~n1762 & n2042;
  assign n2044 = n2043 ^ x3;
  assign n2045 = n2044 ^ x134;
  assign n2079 = ~n1798 & ~n1800;
  assign n2080 = n1769 & ~n2079;
  assign n2081 = n1769 & n1824;
  assign n2082 = ~n1782 & ~n1841;
  assign n2083 = n1794 & ~n2082;
  assign n2084 = ~n2081 & ~n2083;
  assign n2085 = n1802 & n1819;
  assign n2086 = n1785 & ~n2085;
  assign n2087 = ~n1801 & ~n1817;
  assign n2088 = n1799 & n2087;
  assign n2089 = n1778 & ~n2088;
  assign n2090 = n1794 & ~n2085;
  assign n2091 = n1785 & n1841;
  assign n2092 = ~n1780 & ~n1825;
  assign n2093 = n1769 & ~n2092;
  assign n2094 = ~n2091 & ~n2093;
  assign n2095 = ~n1787 & n2094;
  assign n2096 = ~n1816 & ~n2095;
  assign n2097 = ~n1778 & ~n1780;
  assign n2098 = n1780 & n1785;
  assign n2099 = n1813 & ~n2098;
  assign n2100 = ~n1782 & n2099;
  assign n2101 = ~n2097 & ~n2100;
  assign n2102 = ~n1789 & ~n2101;
  assign n2103 = ~n1809 & ~n2102;
  assign n2104 = ~n2096 & ~n2103;
  assign n2105 = ~n2090 & n2104;
  assign n2106 = ~n1777 & n2105;
  assign n2107 = ~n2089 & n2106;
  assign n2108 = ~n2086 & n2107;
  assign n2109 = n2084 & n2108;
  assign n2110 = n1808 & n2109;
  assign n2111 = ~n2080 & n2110;
  assign n2112 = n2111 ^ x11;
  assign n2113 = n2112 ^ x133;
  assign n2122 = ~n2045 & n2113;
  assign n2046 = n1226 ^ x130;
  assign n2047 = n917 ^ x131;
  assign n2151 = n2046 & ~n2047;
  assign n2152 = ~n2122 & n2151;
  assign n2153 = ~n2077 & n2152;
  assign n2125 = n2113 ^ n2045;
  assign n2126 = n2047 & ~n2125;
  assign n2121 = ~n2047 & n2077;
  assign n2154 = n2121 & n2122;
  assign n2155 = ~n2126 & ~n2154;
  assign n2156 = n2046 & ~n2155;
  assign n2078 = n2047 & n2077;
  assign n2157 = n2078 & n2125;
  assign n2123 = ~n2046 & n2122;
  assign n2158 = n2045 & n2121;
  assign n2159 = n2047 & ~n2113;
  assign n2160 = ~n2158 & ~n2159;
  assign n2161 = ~n2046 & ~n2160;
  assign n2162 = ~n2123 & ~n2161;
  assign n2163 = ~n2157 & ~n2162;
  assign n2164 = ~n2156 & ~n2163;
  assign n2165 = ~n2153 & n2164;
  assign n2115 = n2047 & ~n2077;
  assign n2116 = n2113 & n2115;
  assign n2114 = n2078 & ~n2113;
  assign n2117 = n2116 ^ n2114;
  assign n2118 = n2046 & n2117;
  assign n2119 = n2118 ^ n2116;
  assign n2120 = ~n2045 & n2119;
  assign n2124 = n2121 & n2123;
  assign n2127 = ~n2077 & n2126;
  assign n2128 = ~n2115 & ~n2121;
  assign n2129 = n2045 & ~n2113;
  assign n2130 = n2128 & n2129;
  assign n2131 = ~n2127 & ~n2130;
  assign n2132 = ~n2045 & ~n2113;
  assign n2133 = n2132 ^ n2129;
  assign n2134 = ~n2077 & n2133;
  assign n2135 = n2134 ^ n2129;
  assign n2136 = n2131 & ~n2135;
  assign n2137 = n2136 ^ n2046;
  assign n2138 = n2137 ^ n2136;
  assign n2139 = n2115 & n2129;
  assign n2140 = n2045 & n2113;
  assign n2141 = n2077 & n2140;
  assign n2142 = n2129 ^ n2077;
  assign n2143 = ~n2047 & ~n2142;
  assign n2144 = ~n2141 & ~n2143;
  assign n2145 = ~n2139 & n2144;
  assign n2146 = n2145 ^ n2136;
  assign n2147 = n2138 & n2146;
  assign n2148 = n2147 ^ n2136;
  assign n2149 = ~n2124 & n2148;
  assign n2150 = ~n2120 & n2149;
  assign n2166 = n2165 ^ n2150;
  assign n2167 = n2009 & ~n2166;
  assign n2168 = n2167 ^ n2165;
  assign n2169 = n2168 ^ x36;
  assign n2170 = n2169 ^ x188;
  assign n2171 = n1850 ^ x117;
  assign n2172 = n1579 ^ x112;
  assign n2173 = n2171 & n2172;
  assign n2174 = n1396 ^ x113;
  assign n2175 = n1716 ^ x116;
  assign n2176 = n2174 & n2175;
  assign n2177 = n835 & n870;
  assign n2178 = n869 & ~n886;
  assign n2179 = ~n2177 & ~n2178;
  assign n2180 = ~n863 & n869;
  assign n2181 = ~n885 & ~n1406;
  assign n2182 = n834 & ~n2181;
  assign n2183 = ~n873 & ~n880;
  assign n2184 = ~n877 & n2183;
  assign n2185 = ~n860 & n2184;
  assign n2186 = n835 & ~n2185;
  assign n2187 = ~n884 & ~n895;
  assign n2188 = ~n842 & n2187;
  assign n2189 = n887 & n1414;
  assign n2190 = n2188 & n2189;
  assign n2191 = n872 & ~n2190;
  assign n2192 = ~n2186 & ~n2191;
  assign n2193 = n1410 ^ n869;
  assign n2194 = n1410 ^ n844;
  assign n2195 = n2194 ^ n844;
  assign n2196 = n844 ^ n842;
  assign n2197 = n2195 & ~n2196;
  assign n2198 = n2197 ^ n844;
  assign n2199 = ~n2193 & n2198;
  assign n2200 = n2199 ^ n869;
  assign n2201 = n2192 & ~n2200;
  assign n2202 = ~n852 & n2201;
  assign n2203 = ~n2182 & n2202;
  assign n2204 = ~n2180 & n2203;
  assign n2205 = ~n1404 & n2204;
  assign n2206 = n2179 & n2205;
  assign n2207 = n2206 ^ x49;
  assign n2208 = n2207 ^ x114;
  assign n2209 = ~n971 & ~n2060;
  assign n2210 = n955 & ~n2056;
  assign n2211 = ~n2209 & ~n2210;
  assign n2215 = ~n959 & n998;
  assign n2212 = ~n935 & n2053;
  assign n2213 = ~n951 & n2212;
  assign n2214 = n957 & n2213;
  assign n2216 = n2215 ^ n2214;
  assign n2217 = n2215 ^ n919;
  assign n2218 = n2217 ^ n2215;
  assign n2219 = n2216 & ~n2218;
  assign n2220 = n2219 ^ n2215;
  assign n2221 = n920 & ~n2220;
  assign n2222 = n964 ^ n930;
  assign n2223 = n2222 ^ n964;
  assign n2224 = n926 ^ n922;
  assign n2225 = n2224 ^ n925;
  assign n2226 = n2225 ^ n926;
  assign n2227 = n926 ^ n925;
  assign n2228 = n2227 ^ n926;
  assign n2229 = n926 ^ n923;
  assign n2230 = n2229 ^ n926;
  assign n2231 = n2228 & n2230;
  assign n2232 = n2231 ^ n926;
  assign n2233 = ~n2226 & ~n2232;
  assign n2234 = n2233 ^ n2224;
  assign n2235 = n2234 ^ n964;
  assign n2236 = n2223 & ~n2235;
  assign n2237 = n2236 ^ n964;
  assign n2238 = ~n2221 & ~n2237;
  assign n2239 = n2211 & n2238;
  assign n2240 = n947 & n2239;
  assign n2241 = ~n929 & n2240;
  assign n2242 = n2241 ^ x41;
  assign n2243 = n2242 ^ x115;
  assign n2244 = n2208 & n2243;
  assign n2245 = n2176 & n2244;
  assign n2246 = n2173 & n2245;
  assign n2247 = n2171 & ~n2172;
  assign n2248 = ~n2208 & n2243;
  assign n2249 = ~n2174 & ~n2175;
  assign n2250 = n2248 & n2249;
  assign n2251 = n2247 & n2250;
  assign n2252 = ~n2246 & ~n2251;
  assign n2253 = n2174 & ~n2175;
  assign n2254 = ~n2208 & ~n2243;
  assign n2255 = n2253 & n2254;
  assign n2256 = n2173 & n2255;
  assign n2257 = n2244 & n2253;
  assign n2258 = n2208 & ~n2243;
  assign n2259 = n2253 & n2258;
  assign n2260 = n2176 & n2254;
  assign n2261 = ~n2259 & ~n2260;
  assign n2262 = ~n2257 & n2261;
  assign n2263 = n2247 & ~n2262;
  assign n2264 = ~n2256 & ~n2263;
  assign n2265 = n2249 & n2258;
  assign n2266 = n2173 & n2265;
  assign n2267 = ~n2171 & n2172;
  assign n2268 = ~n2174 & n2175;
  assign n2269 = n2254 & n2268;
  assign n2270 = n2267 & n2269;
  assign n2271 = ~n2266 & ~n2270;
  assign n2272 = ~n2171 & ~n2172;
  assign n2273 = n2244 & n2249;
  assign n2274 = n2272 & n2273;
  assign n2275 = n2176 & n2248;
  assign n2276 = n2244 & n2268;
  assign n2277 = n2249 & n2254;
  assign n2278 = ~n2276 & ~n2277;
  assign n2279 = ~n2275 & n2278;
  assign n2280 = ~n2257 & n2279;
  assign n2281 = n2173 & ~n2280;
  assign n2282 = ~n2274 & ~n2281;
  assign n2283 = n2258 & n2268;
  assign n2284 = ~n2265 & ~n2283;
  assign n2285 = ~n2171 & ~n2284;
  assign n2286 = n2248 & n2253;
  assign n2287 = n2176 & n2258;
  assign n2288 = ~n2276 & ~n2287;
  assign n2289 = ~n2286 & n2288;
  assign n2290 = n2247 & ~n2289;
  assign n2291 = n2272 & n2286;
  assign n2292 = ~n2259 & ~n2275;
  assign n2293 = ~n2245 & n2292;
  assign n2294 = n2272 & ~n2293;
  assign n2295 = ~n2255 & ~n2287;
  assign n2296 = ~n2257 & n2295;
  assign n2297 = ~n2245 & n2296;
  assign n2298 = n2267 & ~n2297;
  assign n2299 = ~n2294 & ~n2298;
  assign n2300 = ~n2291 & n2299;
  assign n2301 = ~n2290 & n2300;
  assign n2302 = ~n2285 & n2301;
  assign n2303 = n2282 & n2302;
  assign n2304 = n2283 ^ n2171;
  assign n2305 = n2304 ^ n2283;
  assign n2306 = n2283 ^ n2269;
  assign n2307 = ~n2305 & n2306;
  assign n2308 = n2307 ^ n2283;
  assign n2309 = ~n2172 & n2308;
  assign n2310 = n2303 & ~n2309;
  assign n2311 = n2248 & n2268;
  assign n2312 = n2311 ^ n2171;
  assign n2313 = n2312 ^ n2311;
  assign n2314 = n2311 ^ n2269;
  assign n2315 = n2313 & n2314;
  assign n2316 = n2315 ^ n2311;
  assign n2317 = n2172 & n2316;
  assign n2318 = n2310 & ~n2317;
  assign n2319 = n2271 & n2318;
  assign n2320 = n2264 & n2319;
  assign n2321 = n2252 & n2320;
  assign n2322 = n2321 ^ x60;
  assign n2323 = n2322 ^ x185;
  assign n2324 = n2170 & ~n2323;
  assign n2325 = ~n1975 & n2324;
  assign n2326 = n1689 & n2325;
  assign n2327 = n1383 & ~n1688;
  assign n2328 = n1028 ^ n1015;
  assign n2329 = n2328 ^ n1028;
  assign n2330 = n1060 ^ n1028;
  assign n2331 = ~n2329 & ~n2330;
  assign n2332 = n2331 ^ n1028;
  assign n2333 = ~n1047 & ~n2332;
  assign n2334 = ~n1048 & n2333;
  assign n2335 = n1045 & ~n2334;
  assign n2336 = ~n1036 & n1038;
  assign n2337 = ~n1029 & ~n1036;
  assign n2338 = n1034 & ~n2337;
  assign n2339 = ~n2336 & ~n2338;
  assign n2340 = ~n1027 & n2339;
  assign n2341 = ~n1046 & n2340;
  assign n2342 = n1055 & ~n2341;
  assign n2343 = ~n2335 & ~n2342;
  assign n2344 = n1038 & ~n2337;
  assign n2345 = ~n1035 & ~n2344;
  assign n2346 = ~n1026 & n2345;
  assign n2347 = ~n1046 & n2346;
  assign n2348 = n2347 ^ n1008;
  assign n2349 = n2348 ^ n2347;
  assign n2350 = n1012 & ~n1015;
  assign n2351 = n2350 ^ n1011;
  assign n2352 = n2351 ^ n2350;
  assign n2353 = n2350 ^ n1034;
  assign n2354 = ~n2352 & n2353;
  assign n2355 = n2354 ^ n2350;
  assign n2356 = ~n2344 & ~n2355;
  assign n2357 = n1031 & n2356;
  assign n2358 = n2357 ^ n2347;
  assign n2359 = n2349 & ~n2358;
  assign n2360 = n2359 ^ n2347;
  assign n2361 = ~n1387 & n2360;
  assign n2362 = n2343 & ~n2361;
  assign n2363 = n2362 ^ x37;
  assign n2364 = n2363 ^ x142;
  assign n2365 = n920 & ~n952;
  assign n2366 = ~n935 & n960;
  assign n2367 = ~n964 & n2366;
  assign n2368 = n955 & ~n2367;
  assign n2369 = n969 & n971;
  assign n2370 = n957 & n2369;
  assign n2371 = n930 & ~n2370;
  assign n2372 = ~n932 & n969;
  assign n2373 = ~n987 & n2372;
  assign n2374 = n965 & ~n2373;
  assign n2375 = ~n2371 & ~n2374;
  assign n2376 = n944 & n955;
  assign n2377 = ~n955 & n2065;
  assign n2378 = ~n956 & n2052;
  assign n2379 = ~n921 & n2378;
  assign n2380 = ~n2377 & ~n2379;
  assign n2381 = ~n2060 & n2380;
  assign n2382 = ~n2376 & ~n2381;
  assign n2383 = n2375 & n2382;
  assign n2384 = n938 & n2383;
  assign n2385 = ~n2368 & n2384;
  assign n2386 = ~n2365 & n2385;
  assign n2387 = n2051 & n2386;
  assign n2388 = n2387 ^ x63;
  assign n2389 = n2388 ^ x147;
  assign n2390 = ~n2364 & n2389;
  assign n2391 = ~n1776 & ~n1818;
  assign n2392 = n1794 & ~n2391;
  assign n2393 = n1768 & n1812;
  assign n2394 = ~n1816 & ~n1842;
  assign n2395 = ~n2393 & ~n2394;
  assign n2396 = n1801 ^ n1767;
  assign n2397 = n2396 ^ n1801;
  assign n2398 = ~n1796 & ~n1824;
  assign n2399 = n1802 & n2398;
  assign n2400 = n1790 & n2399;
  assign n2401 = ~n1780 & n2400;
  assign n2402 = n2401 ^ n1801;
  assign n2403 = ~n2397 & ~n2402;
  assign n2404 = n2403 ^ n1801;
  assign n2405 = n1768 & n2404;
  assign n2406 = n2395 & ~n2405;
  assign n2407 = n1794 & ~n1810;
  assign n2408 = ~n1785 & ~n1794;
  assign n2409 = ~n1783 & ~n2408;
  assign n2410 = ~n1816 & n1824;
  assign n2411 = n1769 & n1818;
  assign n2412 = ~n1805 & n1819;
  assign n2413 = n1785 & ~n2412;
  assign n2414 = ~n2411 & ~n2413;
  assign n2415 = ~n2410 & n2414;
  assign n2416 = ~n2080 & n2415;
  assign n2417 = ~n2409 & n2416;
  assign n2418 = ~n2407 & n2417;
  assign n2419 = n2406 & n2418;
  assign n2420 = ~n1807 & n2419;
  assign n2421 = ~n2392 & n2420;
  assign n2422 = n2421 ^ x29;
  assign n2423 = n2422 ^ x143;
  assign n2424 = n1079 & ~n1123;
  assign n2425 = ~n1097 & ~n1099;
  assign n2426 = n1125 & ~n2425;
  assign n2427 = ~n1110 & ~n1117;
  assign n2428 = n1080 & ~n2427;
  assign n2429 = n1512 & n1530;
  assign n2430 = ~n1086 & n2429;
  assign n2431 = n1108 & ~n2430;
  assign n2432 = ~n2428 & ~n2431;
  assign n2433 = ~n1077 & n1111;
  assign n2434 = ~n1098 & n2433;
  assign n2435 = n1125 & ~n2434;
  assign n2436 = n1119 & n1977;
  assign n2437 = ~n1097 & n2436;
  assign n2438 = n1084 & ~n2437;
  assign n2439 = ~n2435 & ~n2438;
  assign n2440 = n2432 & n2439;
  assign n2441 = ~n2426 & n2440;
  assign n2442 = ~n2424 & n2441;
  assign n2443 = ~n1987 & n2442;
  assign n2444 = n1529 & n2443;
  assign n2445 = ~n1092 & n2444;
  assign n2446 = ~n1115 & n2445;
  assign n2447 = n2446 ^ x13;
  assign n2448 = n2447 ^ x145;
  assign n2449 = n2423 & ~n2448;
  assign n2450 = n1439 & n1445;
  assign n2451 = n1451 & n1482;
  assign n2452 = ~n2450 & ~n2451;
  assign n2453 = ~n1442 & n1483;
  assign n2454 = n1446 & n1475;
  assign n2455 = ~n2453 & ~n2454;
  assign n2456 = n2452 & n2455;
  assign n2457 = ~n1446 & n1489;
  assign n2458 = ~n1439 & ~n1483;
  assign n2459 = n1444 & ~n2458;
  assign n2460 = ~n2457 & ~n2459;
  assign n2461 = n1446 & n1748;
  assign n2462 = n1470 & n1479;
  assign n2463 = n1445 & ~n2462;
  assign n2464 = ~n2461 & ~n2463;
  assign n2465 = n2460 & n2464;
  assign n2466 = n1722 & n2465;
  assign n2467 = n1460 & n2466;
  assign n2468 = n1444 ^ n1441;
  assign n2469 = n2468 ^ n1441;
  assign n2470 = n1484 ^ n1441;
  assign n2471 = ~n2469 & n2470;
  assign n2472 = n2471 ^ n1441;
  assign n2473 = n2467 & ~n2472;
  assign n2474 = n2456 & n2473;
  assign n2475 = n1472 & n2474;
  assign n2476 = n2475 ^ x5;
  assign n2477 = n2476 ^ x146;
  assign n2478 = ~n1191 & ~n1567;
  assign n2479 = n1150 & ~n2478;
  assign n2480 = ~n1166 & ~n1214;
  assign n2481 = n1194 & ~n2480;
  assign n2482 = ~n1168 & ~n1183;
  assign n2483 = ~n1182 & ~n1187;
  assign n2484 = ~n1150 & n2483;
  assign n2485 = ~n2482 & ~n2484;
  assign n2486 = ~n1865 & ~n2485;
  assign n2487 = ~n1184 & ~n2486;
  assign n2488 = ~n2481 & ~n2487;
  assign n2489 = ~n2479 & n2488;
  assign n2490 = ~n1162 & ~n1207;
  assign n2491 = n2490 ^ n1150;
  assign n2492 = n2491 ^ n2490;
  assign n2493 = ~n1182 & ~n1191;
  assign n2494 = n2493 ^ n2490;
  assign n2495 = n2494 ^ n2490;
  assign n2496 = ~n2492 & ~n2495;
  assign n2497 = n2496 ^ n2490;
  assign n2498 = ~n1183 & ~n2497;
  assign n2499 = n2498 ^ n2490;
  assign n2500 = n2489 & n2499;
  assign n2501 = n1174 ^ n1149;
  assign n2502 = n2501 ^ n1174;
  assign n2503 = n1187 ^ n1174;
  assign n2504 = n2503 ^ n1174;
  assign n2505 = n2502 & n2504;
  assign n2506 = n2505 ^ n1174;
  assign n2507 = ~n1148 & n2506;
  assign n2508 = n2507 ^ n1174;
  assign n2509 = n2500 & ~n2508;
  assign n2510 = ~n1170 & n2509;
  assign n2511 = n1558 & n2510;
  assign n2512 = ~n1886 & n2511;
  assign n2513 = ~n1556 & n2512;
  assign n2514 = n1164 & n2513;
  assign n2515 = n2514 ^ x21;
  assign n2516 = n2515 ^ x144;
  assign n2517 = n2477 & ~n2516;
  assign n2518 = n2449 & n2517;
  assign n2519 = n2423 & n2448;
  assign n2520 = ~n2477 & ~n2516;
  assign n2521 = n2519 & n2520;
  assign n2522 = ~n2518 & ~n2521;
  assign n2523 = n2390 & ~n2522;
  assign n2524 = ~n2423 & n2448;
  assign n2525 = n2520 & n2524;
  assign n2526 = n2390 & n2525;
  assign n2527 = n2364 & ~n2389;
  assign n2528 = ~n2423 & ~n2448;
  assign n2529 = ~n2477 & n2516;
  assign n2530 = n2528 & n2529;
  assign n2531 = n2527 & n2530;
  assign n2532 = n2364 & n2389;
  assign n2533 = ~n2364 & ~n2389;
  assign n2534 = ~n2532 & ~n2533;
  assign n2535 = n2520 & n2528;
  assign n2536 = ~n2534 & n2535;
  assign n2537 = ~n2531 & ~n2536;
  assign n2538 = ~n2526 & n2537;
  assign n2539 = n2519 & n2529;
  assign n2540 = ~n2518 & ~n2539;
  assign n2541 = n2533 & ~n2540;
  assign n2542 = n2477 & n2516;
  assign n2543 = n2449 & n2542;
  assign n2544 = n2390 & n2543;
  assign n2545 = n2533 & n2543;
  assign n2546 = n2528 & n2542;
  assign n2547 = n2517 & n2524;
  assign n2548 = ~n2535 & ~n2547;
  assign n2549 = ~n2546 & n2548;
  assign n2550 = ~n2539 & n2549;
  assign n2551 = n2390 & ~n2550;
  assign n2552 = ~n2545 & ~n2551;
  assign n2553 = n2524 & n2542;
  assign n2554 = ~n2389 & n2553;
  assign n2555 = n2524 & n2529;
  assign n2556 = ~n2547 & ~n2555;
  assign n2557 = n2449 & n2529;
  assign n2558 = n2449 & n2520;
  assign n2559 = ~n2557 & ~n2558;
  assign n2560 = n2522 & n2559;
  assign n2561 = n2556 & n2560;
  assign n2562 = n2527 & ~n2561;
  assign n2563 = n2517 & n2528;
  assign n2564 = ~n2525 & ~n2563;
  assign n2565 = ~n2557 & n2564;
  assign n2566 = n2532 & ~n2565;
  assign n2567 = n2517 & n2519;
  assign n2568 = n2519 & n2542;
  assign n2569 = n2532 & n2568;
  assign n2570 = n2521 & n2533;
  assign n2571 = ~n2569 & ~n2570;
  assign n2572 = ~n2567 & n2571;
  assign n2573 = ~n2534 & ~n2572;
  assign n2574 = ~n2566 & ~n2573;
  assign n2575 = ~n2562 & n2574;
  assign n2576 = ~n2554 & n2575;
  assign n2577 = n2552 & n2576;
  assign n2578 = ~n2544 & n2577;
  assign n2579 = ~n2541 & n2578;
  assign n2580 = n2546 ^ n2532;
  assign n2581 = n2546 ^ n2533;
  assign n2582 = n2581 ^ n2533;
  assign n2583 = n2539 ^ n2533;
  assign n2584 = ~n2582 & ~n2583;
  assign n2585 = n2584 ^ n2533;
  assign n2586 = n2580 & n2585;
  assign n2587 = n2586 ^ n2532;
  assign n2588 = n2579 & ~n2587;
  assign n2589 = n2538 & n2588;
  assign n2590 = ~n2523 & n2589;
  assign n2591 = n2590 ^ x44;
  assign n2592 = n2591 ^ x187;
  assign n2593 = ~n1975 & n2323;
  assign n2594 = n2170 & n2593;
  assign n2595 = n2592 & n2594;
  assign n2596 = ~n2323 & n2592;
  assign n2597 = ~n2170 & n2596;
  assign n2598 = n1975 & n2597;
  assign n2599 = n1975 & n2170;
  assign n2600 = ~n2323 & n2599;
  assign n2601 = ~n2592 & n2600;
  assign n2602 = ~n2598 & ~n2601;
  assign n2603 = ~n2595 & n2602;
  assign n2604 = n2327 & ~n2603;
  assign n2605 = ~n2326 & ~n2604;
  assign n2606 = ~n1975 & n2597;
  assign n2607 = ~n1689 & ~n2327;
  assign n2608 = n2606 & ~n2607;
  assign n2609 = n1383 & n1688;
  assign n2610 = ~n2592 & n2594;
  assign n2611 = ~n2170 & ~n2592;
  assign n2612 = n2593 & n2611;
  assign n2613 = ~n2170 & n2323;
  assign n2614 = n1975 & n2613;
  assign n2615 = n2592 & n2614;
  assign n2616 = n2323 & n2599;
  assign n2617 = ~n2592 & n2616;
  assign n2618 = ~n2615 & ~n2617;
  assign n2619 = ~n2612 & n2618;
  assign n2620 = ~n2610 & n2619;
  assign n2621 = n2609 & ~n2620;
  assign n2622 = ~n2608 & ~n2621;
  assign n2623 = n2605 & n2622;
  assign n2624 = ~n1383 & n2598;
  assign n2625 = ~n1383 & ~n1688;
  assign n2626 = ~n2323 & n2611;
  assign n2627 = n1975 & n2626;
  assign n2628 = n2596 & n2599;
  assign n2629 = ~n1975 & n2626;
  assign n2630 = ~n2628 & ~n2629;
  assign n2631 = ~n2627 & n2630;
  assign n2632 = n2625 & ~n2631;
  assign n2633 = n1689 & n2627;
  assign n2634 = ~n2609 & ~n2633;
  assign n2635 = n2170 & n2596;
  assign n2636 = ~n1975 & n2635;
  assign n2637 = ~n2606 & ~n2629;
  assign n2638 = ~n2633 & n2637;
  assign n2639 = ~n2636 & n2638;
  assign n2640 = ~n2601 & n2639;
  assign n2641 = ~n2634 & ~n2640;
  assign n2642 = ~n2170 & n2593;
  assign n2643 = n2592 & n2642;
  assign n2644 = n2592 & n2616;
  assign n2645 = ~n2612 & ~n2644;
  assign n2646 = ~n2643 & n2645;
  assign n2647 = n1689 & ~n2646;
  assign n2648 = n2625 ^ n2327;
  assign n2649 = n2323 & n2611;
  assign n2650 = n1975 & n2649;
  assign n2654 = n2645 & ~n2650;
  assign n2655 = ~n2617 & n2654;
  assign n2651 = ~n2610 & ~n2650;
  assign n2652 = ~n2595 & n2651;
  assign n2653 = ~n2643 & n2652;
  assign n2656 = n2655 ^ n2653;
  assign n2657 = n2655 ^ n2327;
  assign n2658 = n2657 ^ n2655;
  assign n2659 = ~n2656 & ~n2658;
  assign n2660 = n2659 ^ n2655;
  assign n2661 = n2648 & ~n2660;
  assign n2662 = n2661 ^ n2625;
  assign n2663 = ~n2647 & ~n2662;
  assign n2664 = ~n2641 & n2663;
  assign n2665 = ~n2632 & n2664;
  assign n2666 = ~n2624 & n2665;
  assign n2667 = n2623 & n2666;
  assign n2668 = n2667 ^ n1004;
  assign n2669 = n2668 ^ x220;
  assign n2670 = n2245 & n2247;
  assign n2671 = n2257 & n2267;
  assign n2672 = n2173 & ~n2284;
  assign n2673 = ~n2671 & ~n2672;
  assign n2674 = ~n2670 & n2673;
  assign n2675 = n2257 & n2272;
  assign n2676 = n2260 & n2267;
  assign n2677 = ~n2675 & ~n2676;
  assign n2678 = n2250 & n2267;
  assign n2679 = n2173 & n2286;
  assign n2680 = ~n2309 & ~n2679;
  assign n2681 = ~n2678 & n2680;
  assign n2682 = n2173 & n2273;
  assign n2683 = ~n2273 & ~n2311;
  assign n2684 = n2295 & n2683;
  assign n2685 = n2272 & ~n2684;
  assign n2686 = ~n2682 & ~n2685;
  assign n2687 = ~n2265 & n2288;
  assign n2688 = n2267 & ~n2687;
  assign n2689 = ~n2269 & n2279;
  assign n2690 = n2247 & ~n2689;
  assign n2691 = ~n2688 & ~n2690;
  assign n2692 = n2686 & n2691;
  assign n2693 = ~n2256 & n2692;
  assign n2694 = ~n2317 & n2693;
  assign n2695 = n2681 & n2694;
  assign n2696 = n2677 & n2695;
  assign n2697 = n2674 & n2696;
  assign n2698 = ~n2291 & n2697;
  assign n2699 = n2252 & n2698;
  assign n2700 = ~n2259 & n2699;
  assign n2701 = n2700 ^ x58;
  assign n2702 = n2701 ^ x171;
  assign n2703 = n2527 & n2543;
  assign n2704 = ~n2544 & ~n2703;
  assign n2705 = n2390 & n2535;
  assign n2706 = ~n2541 & ~n2705;
  assign n2707 = n2527 & n2567;
  assign n2708 = n2518 & n2532;
  assign n2709 = ~n2707 & ~n2708;
  assign n2710 = ~n2539 & ~n2558;
  assign n2711 = n2364 & ~n2710;
  assign n2712 = ~n2390 & ~n2527;
  assign n2713 = ~n2553 & ~n2557;
  assign n2714 = ~n2390 & n2713;
  assign n2715 = ~n2712 & ~n2714;
  assign n2716 = n2715 ^ n2527;
  assign n2717 = n2715 ^ n2548;
  assign n2718 = n2717 ^ n2548;
  assign n2719 = ~n2521 & n2559;
  assign n2720 = n2719 ^ n2548;
  assign n2721 = n2718 & ~n2720;
  assign n2722 = n2721 ^ n2548;
  assign n2723 = n2716 & n2722;
  assign n2724 = n2723 ^ n2527;
  assign n2725 = ~n2711 & ~n2724;
  assign n2726 = ~n2553 & n2556;
  assign n2727 = n2390 & ~n2726;
  assign n2728 = n2516 ^ n2477;
  assign n2729 = n2528 & n2728;
  assign n2730 = ~n2555 & ~n2729;
  assign n2731 = n2730 ^ n2565;
  assign n2732 = n2389 ^ n2364;
  assign n2733 = n2565 ^ n2389;
  assign n2734 = n2732 & ~n2733;
  assign n2735 = n2734 ^ n2389;
  assign n2736 = n2731 & ~n2735;
  assign n2737 = n2736 ^ n2730;
  assign n2738 = ~n2546 & n2737;
  assign n2739 = ~n2568 & n2738;
  assign n2740 = ~n2534 & ~n2739;
  assign n2741 = ~n2727 & ~n2740;
  assign n2742 = n2725 & n2741;
  assign n2743 = n2709 & n2742;
  assign n2744 = ~n2570 & n2743;
  assign n2745 = n2706 & n2744;
  assign n2746 = n2704 & n2745;
  assign n2747 = n2746 ^ x32;
  assign n2748 = n2747 ^ x166;
  assign n2749 = n2702 & ~n2748;
  assign n2750 = n2422 ^ x141;
  assign n2751 = n2044 ^ x136;
  assign n2752 = ~n2750 & ~n2751;
  assign n2753 = n2363 ^ x140;
  assign n2754 = n855 & ~n1407;
  assign n2755 = n834 & n847;
  assign n2756 = ~n2754 & ~n2755;
  assign n2757 = n863 & ~n877;
  assign n2758 = n835 & ~n2757;
  assign n2759 = n881 & ~n1406;
  assign n2760 = n869 & ~n2759;
  assign n2761 = ~n2758 & ~n2760;
  assign n2762 = n851 & ~n853;
  assign n2763 = n872 & ~n2762;
  assign n2764 = ~n860 & n2188;
  assign n2765 = n844 & ~n2764;
  assign n2766 = ~n2763 & ~n2765;
  assign n2767 = n2761 & n2766;
  assign n2768 = n2756 & n2767;
  assign n2769 = n2179 & n2768;
  assign n2770 = n1405 & n2769;
  assign n2771 = n868 & n2770;
  assign n2772 = ~n843 & n2771;
  assign n2773 = n2772 ^ x53;
  assign n2774 = n2773 ^ x138;
  assign n2775 = n2753 & n2774;
  assign n2776 = ~n1229 & n1245;
  assign n2777 = n1230 & ~n1588;
  assign n2778 = ~n2776 & ~n2777;
  assign n2779 = n1250 & n1257;
  assign n2780 = ~n1251 & ~n1259;
  assign n2781 = n1260 & ~n2780;
  assign n2782 = ~n1270 & n1695;
  assign n2783 = ~n1253 & n2782;
  assign n2784 = n1247 & n2783;
  assign n2785 = n1261 & n2784;
  assign n2786 = ~n1266 & n2785;
  assign n2787 = ~n1278 & n1287;
  assign n2788 = ~n1705 & ~n2787;
  assign n2789 = n1277 & ~n2788;
  assign n2790 = ~n2786 & ~n2789;
  assign n2791 = ~n2781 & ~n2790;
  assign n2792 = ~n2779 & n2791;
  assign n2793 = n2778 & n2792;
  assign n2794 = ~n1249 & n2793;
  assign n2795 = n1583 & n2794;
  assign n2796 = n2795 ^ x45;
  assign n2797 = n2796 ^ x139;
  assign n2798 = n2008 ^ x137;
  assign n2799 = ~n2797 & n2798;
  assign n2800 = n2775 & n2799;
  assign n2801 = ~n2753 & ~n2774;
  assign n2802 = n2799 & n2801;
  assign n2803 = ~n2800 & ~n2802;
  assign n2804 = n2752 & ~n2803;
  assign n2805 = ~n2750 & n2751;
  assign n2806 = ~n2753 & n2774;
  assign n2807 = n2799 & n2806;
  assign n2808 = n2753 & ~n2774;
  assign n2809 = n2799 & n2808;
  assign n2810 = ~n2807 & ~n2809;
  assign n2811 = n2805 & ~n2810;
  assign n2812 = ~n2804 & ~n2811;
  assign n2813 = n2750 & ~n2751;
  assign n2814 = ~n2797 & ~n2798;
  assign n2815 = n2801 & n2814;
  assign n2816 = n2797 & ~n2798;
  assign n2817 = n2808 & n2816;
  assign n2818 = ~n2815 & ~n2817;
  assign n2819 = n2813 & ~n2818;
  assign n2820 = n2750 & n2751;
  assign n2821 = n2806 & n2814;
  assign n2822 = n2820 & n2821;
  assign n2823 = n2797 & n2798;
  assign n2824 = n2808 & n2823;
  assign n2825 = n2752 & n2824;
  assign n2826 = n2806 & n2823;
  assign n2827 = ~n2800 & ~n2826;
  assign n2828 = n2805 & ~n2827;
  assign n2829 = ~n2825 & ~n2828;
  assign n2830 = ~n2822 & n2829;
  assign n2831 = ~n2819 & n2830;
  assign n2832 = n2813 & n2824;
  assign n2833 = n2817 & n2820;
  assign n2834 = ~n2832 & ~n2833;
  assign n2835 = n2806 & n2816;
  assign n2836 = n2808 & n2814;
  assign n2837 = ~n2835 & ~n2836;
  assign n2838 = n2752 & ~n2837;
  assign n2839 = n2775 & n2816;
  assign n2840 = n2801 & n2816;
  assign n2841 = ~n2839 & ~n2840;
  assign n2842 = ~n2809 & n2841;
  assign n2843 = ~n2826 & n2842;
  assign n2844 = n2813 & ~n2843;
  assign n2845 = ~n2838 & ~n2844;
  assign n2846 = n2801 & n2823;
  assign n2847 = ~n2750 & n2846;
  assign n2848 = ~n2821 & ~n2839;
  assign n2849 = ~n2817 & n2848;
  assign n2850 = n2805 & ~n2849;
  assign n2851 = n2775 & n2823;
  assign n2852 = n2810 & ~n2851;
  assign n2853 = ~n2802 & n2852;
  assign n2854 = ~n2840 & n2853;
  assign n2855 = ~n2836 & n2854;
  assign n2856 = n2820 & ~n2855;
  assign n2857 = ~n2850 & ~n2856;
  assign n2858 = ~n2847 & n2857;
  assign n2859 = n2845 & n2858;
  assign n2860 = n2834 & n2859;
  assign n2861 = n2775 & n2814;
  assign n2862 = n2861 ^ n2752;
  assign n2863 = n2861 ^ n2813;
  assign n2864 = n2863 ^ n2813;
  assign n2865 = n2839 ^ n2813;
  assign n2866 = ~n2864 & ~n2865;
  assign n2867 = n2866 ^ n2813;
  assign n2868 = n2862 & n2867;
  assign n2869 = n2868 ^ n2752;
  assign n2870 = n2860 & ~n2869;
  assign n2871 = n2831 & n2870;
  assign n2872 = n2812 & n2871;
  assign n2873 = n2872 ^ x0;
  assign n2874 = n2873 ^ x170;
  assign n2875 = n1622 & n1642;
  assign n2876 = n1629 ^ n1619;
  assign n2877 = n2876 ^ n1619;
  assign n2878 = n1619 ^ n1431;
  assign n2879 = n2878 ^ n1619;
  assign n2880 = n2877 & ~n2879;
  assign n2881 = n2880 ^ n1619;
  assign n2882 = n1397 & n2881;
  assign n2883 = n2882 ^ n1619;
  assign n2884 = ~n2875 & ~n2883;
  assign n2885 = ~n1651 & ~n1664;
  assign n2886 = n1625 & ~n2885;
  assign n2887 = n1432 & n1629;
  assign n2888 = n1642 & ~n1674;
  assign n2889 = ~n2887 & ~n2888;
  assign n2890 = ~n1397 & ~n1669;
  assign n2891 = ~n1629 & ~n1668;
  assign n2892 = ~n1619 & n2891;
  assign n2893 = n1674 & n2892;
  assign n2894 = n1625 & ~n2893;
  assign n2895 = ~n1615 & n1660;
  assign n2896 = ~n1622 & n2895;
  assign n2897 = n1617 & ~n2896;
  assign n2898 = ~n2894 & ~n2897;
  assign n2899 = ~n2890 & n2898;
  assign n2900 = n1652 ^ n1397;
  assign n2901 = n2900 ^ n1652;
  assign n2902 = n1664 ^ n1652;
  assign n2903 = n2902 ^ n1652;
  assign n2904 = ~n2901 & n2903;
  assign n2905 = n2904 ^ n1652;
  assign n2906 = n1431 & ~n2905;
  assign n2907 = n2906 ^ n1652;
  assign n2908 = n2899 & n2907;
  assign n2909 = n2889 & n2908;
  assign n2910 = ~n2886 & n2909;
  assign n2911 = n1641 & n2910;
  assign n2912 = n2884 & n2911;
  assign n2913 = ~n1616 & n2912;
  assign n2914 = n2913 ^ x24;
  assign n2915 = n2914 ^ x167;
  assign n2916 = ~n2874 & n2915;
  assign n2917 = n1055 & ~n2357;
  assign n2918 = n1009 & ~n2334;
  assign n2919 = ~n2917 & ~n2918;
  assign n2920 = n1033 & n2341;
  assign n2921 = n1045 & ~n2347;
  assign n2922 = ~n2920 & ~n2921;
  assign n2923 = n2919 & n2922;
  assign n2924 = n2923 ^ x55;
  assign n2925 = n2924 ^ x150;
  assign n2926 = n1430 ^ x152;
  assign n2927 = n2925 & ~n2926;
  assign n2928 = n2388 ^ x149;
  assign n2929 = n1785 & ~n2398;
  assign n2930 = n1774 ^ n1770;
  assign n2931 = n2930 ^ n1773;
  assign n2932 = n2931 ^ n1770;
  assign n2933 = n2932 ^ n1771;
  assign n2934 = n2930 ^ n1771;
  assign n2935 = n2930 ^ n1770;
  assign n2936 = n2935 ^ n2930;
  assign n2937 = n2934 & n2936;
  assign n2938 = n2937 ^ n2930;
  assign n2939 = n2933 & ~n2938;
  assign n2940 = n2939 ^ n2930;
  assign n2941 = n1794 & ~n2940;
  assign n2942 = ~n2929 & ~n2941;
  assign n2943 = ~n1816 & ~n2087;
  assign n2944 = n1810 & n1819;
  assign n2945 = n1778 & ~n2944;
  assign n2946 = n1769 & n1841;
  assign n2947 = ~n1784 & ~n2946;
  assign n2948 = n1790 & n2947;
  assign n2949 = n2948 ^ n1767;
  assign n2950 = n2949 ^ n2948;
  assign n2951 = n1783 & ~n1789;
  assign n2952 = ~n1812 & n2951;
  assign n2953 = n2952 ^ n2948;
  assign n2954 = n2953 ^ n2948;
  assign n2955 = ~n2950 & ~n2954;
  assign n2956 = n2955 ^ n2948;
  assign n2957 = ~n1768 & ~n2956;
  assign n2958 = n2957 ^ n2948;
  assign n2959 = ~n2945 & n2958;
  assign n2960 = ~n2943 & n2959;
  assign n2961 = n2942 & n2960;
  assign n2962 = ~n2392 & n2961;
  assign n2963 = ~n1777 & n2962;
  assign n2964 = ~n2080 & n2963;
  assign n2965 = n2964 ^ x47;
  assign n2966 = n2965 ^ x151;
  assign n2967 = n2928 & ~n2966;
  assign n2968 = n2927 & n2967;
  assign n2969 = n2476 ^ x148;
  assign n2970 = n1612 ^ x153;
  assign n2971 = n2969 & n2970;
  assign n2972 = n2968 & n2971;
  assign n2973 = ~n2928 & n2966;
  assign n2974 = ~n2925 & ~n2926;
  assign n2975 = n2973 & n2974;
  assign n2976 = ~n2969 & n2970;
  assign n2977 = n2975 & n2976;
  assign n2978 = ~n2972 & ~n2977;
  assign n2979 = ~n2925 & n2926;
  assign n2980 = n2967 & n2979;
  assign n2981 = n2928 & n2966;
  assign n2982 = n2927 & n2981;
  assign n2983 = ~n2980 & ~n2982;
  assign n2984 = n2976 & ~n2983;
  assign n2985 = n2974 & n2981;
  assign n2986 = ~n2980 & ~n2985;
  assign n2987 = ~n2975 & n2986;
  assign n2988 = n2969 & ~n2970;
  assign n2989 = ~n2987 & n2988;
  assign n2990 = ~n2984 & ~n2989;
  assign n2991 = ~n2976 & ~n2988;
  assign n2992 = n2966 ^ n2925;
  assign n2993 = n2992 ^ n2925;
  assign n2994 = n2926 ^ n2925;
  assign n2995 = n2994 ^ n2925;
  assign n2996 = ~n2993 & n2995;
  assign n2997 = n2996 ^ n2925;
  assign n2998 = ~n2928 & n2997;
  assign n2999 = ~n2991 & n2998;
  assign n3000 = n2925 & n2926;
  assign n3001 = n2981 & n3000;
  assign n3002 = n2967 & n2974;
  assign n3003 = ~n3001 & ~n3002;
  assign n3004 = n2979 & n2981;
  assign n3005 = ~n2982 & ~n3004;
  assign n3006 = n3003 & n3005;
  assign n3007 = ~n2969 & ~n2970;
  assign n3008 = ~n3006 & n3007;
  assign n3009 = n2973 & n2979;
  assign n3010 = ~n2928 & ~n2966;
  assign n3011 = n2974 & n3010;
  assign n3012 = ~n3009 & ~n3011;
  assign n3013 = n2927 & n2973;
  assign n3014 = n3000 & n3010;
  assign n3015 = ~n3013 & ~n3014;
  assign n3016 = ~n2985 & n3015;
  assign n3017 = ~n3001 & n3016;
  assign n3018 = n3012 & n3017;
  assign n3019 = n2971 & ~n3018;
  assign n3020 = ~n3008 & ~n3019;
  assign n3021 = ~n2999 & n3020;
  assign n3022 = n3012 & ~n3014;
  assign n3023 = ~n2968 & n3022;
  assign n3024 = n3023 ^ n3007;
  assign n3025 = n3024 ^ n3023;
  assign n3026 = n2967 & n3000;
  assign n3027 = n3026 ^ n3023;
  assign n3028 = ~n3025 & ~n3027;
  assign n3029 = n3028 ^ n3023;
  assign n3030 = n3021 & n3029;
  assign n3031 = n2990 & n3030;
  assign n3032 = n2978 & n3031;
  assign n3033 = n3032 ^ x8;
  assign n3034 = n3033 ^ x169;
  assign n3035 = n1006 & n1369;
  assign n3036 = n1316 & n1321;
  assign n3037 = n1006 & n1362;
  assign n3038 = ~n1330 & ~n1343;
  assign n3039 = n1317 & ~n3038;
  assign n3040 = ~n3037 & ~n3039;
  assign n3041 = ~n3036 & n3040;
  assign n3042 = ~n3035 & n3041;
  assign n3043 = n1321 & n1338;
  assign n3044 = ~n1312 & ~n1349;
  assign n3045 = n1318 & ~n3044;
  assign n3046 = ~n3043 & ~n3045;
  assign n3047 = n1006 & ~n1350;
  assign n3048 = ~n1347 & n1365;
  assign n3049 = ~n1323 & n3048;
  assign n3050 = n1317 & ~n3049;
  assign n3051 = n1321 & ~n3044;
  assign n3052 = ~n1355 & ~n1369;
  assign n3053 = ~n1346 & ~n1364;
  assign n3054 = n3052 & n3053;
  assign n3055 = n1318 & ~n3054;
  assign n3056 = ~n1355 & ~n1360;
  assign n3057 = ~n1321 & n3056;
  assign n3058 = ~n1371 & ~n3057;
  assign n3059 = ~n1346 & ~n3058;
  assign n3060 = n1319 & ~n3059;
  assign n3061 = ~n3055 & ~n3060;
  assign n3062 = ~n3051 & n3061;
  assign n3063 = ~n3050 & n3062;
  assign n3064 = ~n3047 & n3063;
  assign n3065 = n3046 & n3064;
  assign n3066 = n1336 & n3065;
  assign n3067 = n3042 & n3066;
  assign n3068 = ~n1313 & n3067;
  assign n3069 = n3068 ^ x16;
  assign n3070 = n3069 ^ x168;
  assign n3071 = n3034 & n3070;
  assign n3072 = n2916 & n3071;
  assign n3073 = n2749 & n3072;
  assign n3074 = ~n2702 & ~n2748;
  assign n3075 = ~n2874 & ~n2915;
  assign n3076 = n3071 & n3075;
  assign n3077 = n3074 & n3076;
  assign n3078 = n2702 & n2748;
  assign n3079 = ~n3034 & ~n3070;
  assign n3080 = n3075 & n3079;
  assign n3081 = n3078 & n3080;
  assign n3082 = ~n3077 & ~n3081;
  assign n3083 = ~n3073 & n3082;
  assign n3084 = ~n3034 & n3070;
  assign n3085 = n3075 & n3084;
  assign n3086 = n3078 & n3085;
  assign n3087 = n2916 & n3079;
  assign n3088 = n2749 & n3087;
  assign n3089 = ~n3086 & ~n3088;
  assign n3090 = n2874 & n2915;
  assign n3091 = n3034 & ~n3070;
  assign n3092 = n3090 & n3091;
  assign n3093 = n2749 & n3092;
  assign n3094 = ~n2702 & n2748;
  assign n3095 = n2874 & ~n2915;
  assign n3096 = n3071 & n3095;
  assign n3097 = n3075 & n3091;
  assign n3098 = ~n3096 & ~n3097;
  assign n3099 = n3094 & ~n3098;
  assign n3100 = ~n3093 & ~n3099;
  assign n3101 = n2915 & n3084;
  assign n3102 = n2874 & n3101;
  assign n3103 = n2749 & n3102;
  assign n3104 = n3074 & n3080;
  assign n3105 = ~n3103 & ~n3104;
  assign n3106 = n3084 & n3095;
  assign n3107 = ~n3080 & ~n3106;
  assign n3108 = n3094 & ~n3107;
  assign n3109 = n3079 & n3090;
  assign n3110 = n3094 & n3109;
  assign n3111 = n3074 & n3109;
  assign n3112 = n3078 & n3092;
  assign n3113 = ~n3111 & ~n3112;
  assign n3114 = ~n3074 & ~n3078;
  assign n3115 = n3091 & n3095;
  assign n3116 = n3079 & n3095;
  assign n3117 = n2916 & n3091;
  assign n3118 = ~n3102 & ~n3117;
  assign n3119 = ~n3116 & n3118;
  assign n3120 = ~n3115 & n3119;
  assign n3121 = ~n3072 & n3120;
  assign n3122 = ~n3114 & ~n3121;
  assign n3123 = ~n2874 & n3101;
  assign n3124 = ~n3117 & ~n3123;
  assign n3125 = n3094 & ~n3124;
  assign n3126 = ~n3085 & n3098;
  assign n3127 = n2749 & ~n3126;
  assign n3128 = ~n3125 & ~n3127;
  assign n3129 = n2748 ^ n2702;
  assign n3130 = n3071 & n3090;
  assign n3131 = n3130 ^ n2748;
  assign n3132 = n3131 ^ n3130;
  assign n3133 = n3130 ^ n3106;
  assign n3134 = ~n3132 & n3133;
  assign n3135 = n3134 ^ n3130;
  assign n3136 = n3129 & n3135;
  assign n3137 = n3128 & ~n3136;
  assign n3138 = ~n3122 & n3137;
  assign n3139 = n3113 & n3138;
  assign n3140 = ~n3110 & n3139;
  assign n3141 = ~n3108 & n3140;
  assign n3142 = n3105 & n3141;
  assign n3143 = n3100 & n3142;
  assign n3144 = n3089 & n3143;
  assign n3145 = n3083 & n3144;
  assign n3146 = n3145 ^ n917;
  assign n3147 = n3146 ^ x225;
  assign n3148 = n2669 & n3147;
  assign n3149 = n2521 & n2527;
  assign n3150 = n2527 & ~n2548;
  assign n3151 = ~n3149 & ~n3150;
  assign n3152 = n2532 & n2557;
  assign n3153 = ~n2530 & ~n2553;
  assign n3154 = n2390 & ~n3153;
  assign n3155 = ~n3152 & ~n3154;
  assign n3156 = ~n2389 & n2563;
  assign n3157 = ~n2534 & ~n2556;
  assign n3158 = ~n2522 & n2532;
  assign n3159 = ~n3157 & ~n3158;
  assign n3160 = ~n3156 & n3159;
  assign n3161 = n2527 & n2568;
  assign n3162 = ~n2539 & ~n2567;
  assign n3163 = ~n2557 & n3162;
  assign n3164 = n2533 & ~n3163;
  assign n3165 = ~n3161 & ~n3164;
  assign n3166 = n3160 & n3165;
  assign n3167 = n2558 ^ n2390;
  assign n3168 = n2558 ^ n2527;
  assign n3169 = n3168 ^ n2527;
  assign n3170 = n2567 ^ n2527;
  assign n3171 = ~n3169 & ~n3170;
  assign n3172 = n3171 ^ n2527;
  assign n3173 = n3167 & n3172;
  assign n3174 = n3173 ^ n2390;
  assign n3175 = n3166 & ~n3174;
  assign n3176 = ~n2587 & n3175;
  assign n3177 = n3155 & n3176;
  assign n3178 = n2704 & n3177;
  assign n3179 = n3151 & n3178;
  assign n3180 = n2538 & n3179;
  assign n3181 = ~n2523 & n3180;
  assign n3182 = n3181 ^ x30;
  assign n3183 = n3182 ^ x201;
  assign n3184 = ~n1318 & n1369;
  assign n3185 = ~n1319 & ~n3056;
  assign n3186 = ~n3184 & ~n3185;
  assign n3187 = ~n1346 & ~n1363;
  assign n3188 = n1317 & ~n3187;
  assign n3189 = ~n1311 & ~n1348;
  assign n3190 = ~n1321 & n3189;
  assign n3191 = ~n1326 & ~n1346;
  assign n3192 = n1006 & ~n3191;
  assign n3193 = n1366 & ~n3192;
  assign n3194 = ~n3190 & ~n3193;
  assign n3195 = n1319 & n3194;
  assign n3196 = ~n3188 & ~n3195;
  assign n3197 = ~n1343 & ~n1362;
  assign n3198 = n3197 ^ n1317;
  assign n3199 = n3198 ^ n3197;
  assign n3200 = n3197 ^ n1347;
  assign n3201 = n3200 ^ n3197;
  assign n3202 = ~n3199 & n3201;
  assign n3203 = n3202 ^ n3197;
  assign n3204 = ~n1318 & ~n3203;
  assign n3205 = n3204 ^ n3197;
  assign n3206 = n3196 & n3205;
  assign n3207 = n3186 & n3206;
  assign n3208 = n1341 & n3207;
  assign n3209 = n3046 & n3208;
  assign n3210 = n1335 & n3209;
  assign n3211 = n3041 & n3210;
  assign n3212 = n3211 ^ x4;
  assign n3213 = n3212 ^ x196;
  assign n3214 = n3183 & n3213;
  assign n3215 = n2805 & n2824;
  assign n3216 = n2820 & ~n2837;
  assign n3217 = ~n3215 & ~n3216;
  assign n3218 = ~n2835 & n2853;
  assign n3219 = n2813 & ~n3218;
  assign n3220 = ~n2846 & ~n2851;
  assign n3221 = ~n2807 & n3220;
  assign n3222 = ~n2824 & n3221;
  assign n3223 = ~n2861 & n3222;
  assign n3224 = n2820 & ~n3223;
  assign n3225 = ~n3219 & ~n3224;
  assign n3226 = n2810 & ~n2840;
  assign n3227 = ~n2815 & n3226;
  assign n3228 = ~n2802 & n3227;
  assign n3229 = n2752 & ~n3228;
  assign n3230 = n2818 & n3220;
  assign n3231 = ~n2836 & n3230;
  assign n3232 = n2805 & ~n3231;
  assign n3233 = ~n3229 & ~n3232;
  assign n3234 = n3225 & n3233;
  assign n3235 = n3217 & n3234;
  assign n3236 = ~n2869 & n3235;
  assign n3237 = n2831 & n3236;
  assign n3238 = n3237 ^ x62;
  assign n3239 = n3238 ^ x197;
  assign n3240 = n1554 ^ n1506;
  assign n3241 = n3240 ^ n1580;
  assign n3242 = n1580 ^ n1554;
  assign n3243 = n1613 ^ n1554;
  assign n3244 = n3243 ^ n1554;
  assign n3245 = ~n3242 & ~n3244;
  assign n3246 = n3245 ^ n1554;
  assign n3247 = n3241 & ~n3246;
  assign n3248 = n1617 & n3247;
  assign n3249 = ~n1615 & ~n1634;
  assign n3250 = ~n1658 & n3249;
  assign n3251 = n1642 & ~n3250;
  assign n3252 = ~n3248 & ~n3251;
  assign n3253 = n1649 & ~n1651;
  assign n3254 = n1625 & ~n3253;
  assign n3255 = ~n1657 & ~n1673;
  assign n3256 = ~n1663 & ~n3255;
  assign n3257 = n1669 & n1674;
  assign n3258 = n1432 & ~n3257;
  assign n3259 = ~n3256 & ~n3258;
  assign n3260 = ~n3254 & n3259;
  assign n3261 = n3252 & n3260;
  assign n3262 = n1640 & n3261;
  assign n3263 = n1654 & n3262;
  assign n3264 = ~n1631 & n3263;
  assign n3265 = n1646 & n3264;
  assign n3266 = n2884 & n3265;
  assign n3267 = n3266 ^ x46;
  assign n3268 = n3267 ^ x199;
  assign n3269 = n3239 & n3268;
  assign n3270 = ~n2009 & n2166;
  assign n3271 = n3270 ^ n2165;
  assign n3272 = n3271 ^ x54;
  assign n3273 = n3272 ^ x198;
  assign n3274 = n1719 & ~n1910;
  assign n3275 = ~n1922 & ~n3274;
  assign n3276 = ~n1921 & ~n1955;
  assign n3277 = n1902 & ~n3276;
  assign n3278 = ~n1925 & ~n3277;
  assign n3279 = n1717 & n1913;
  assign n3280 = n1915 & n1927;
  assign n3281 = ~n3279 & ~n3280;
  assign n3282 = n1901 & ~n1947;
  assign n3283 = n1910 & ~n1939;
  assign n3284 = n1902 & ~n3283;
  assign n3285 = n1852 & n1912;
  assign n3286 = ~n1945 & ~n3285;
  assign n3287 = ~n1903 & ~n3286;
  assign n3288 = n1940 & ~n1955;
  assign n3289 = ~n1927 & n3288;
  assign n3290 = n1719 & ~n3289;
  assign n3291 = ~n3287 & ~n3290;
  assign n3292 = ~n3284 & n3291;
  assign n3293 = n1903 & n1916;
  assign n3294 = ~n1938 & n1948;
  assign n3295 = ~n1908 & n3294;
  assign n3296 = n1915 & ~n3295;
  assign n3297 = ~n3293 & ~n3296;
  assign n3298 = n3292 & n3297;
  assign n3299 = n1905 & n3298;
  assign n3300 = ~n3282 & n3299;
  assign n3301 = n3281 & n3300;
  assign n3302 = n3278 & n3301;
  assign n3303 = n3275 & n3302;
  assign n3304 = n3303 ^ x38;
  assign n3305 = n3304 ^ x200;
  assign n3306 = ~n3273 & ~n3305;
  assign n3307 = n3269 & n3306;
  assign n3308 = ~n3273 & n3305;
  assign n3309 = n3239 & ~n3268;
  assign n3310 = n3308 & n3309;
  assign n3311 = ~n3307 & ~n3310;
  assign n3312 = n3214 & ~n3311;
  assign n3313 = n3183 & ~n3213;
  assign n3314 = n3306 & n3309;
  assign n3315 = n3273 & n3305;
  assign n3316 = n3309 & n3315;
  assign n3317 = ~n3314 & ~n3316;
  assign n3318 = n3313 & ~n3317;
  assign n3319 = ~n3312 & ~n3318;
  assign n3320 = n3273 & ~n3305;
  assign n3321 = n3309 & n3320;
  assign n3322 = ~n3183 & ~n3213;
  assign n3323 = n3321 & n3322;
  assign n3324 = ~n3239 & ~n3268;
  assign n3325 = n3306 & n3324;
  assign n3326 = n3214 & n3325;
  assign n3327 = n3305 ^ n3273;
  assign n3328 = n3269 & n3327;
  assign n3329 = n3322 & n3328;
  assign n3330 = ~n3326 & ~n3329;
  assign n3331 = ~n3239 & n3268;
  assign n3332 = n3308 & n3331;
  assign n3333 = n3313 & n3332;
  assign n3334 = n3310 & n3322;
  assign n3335 = ~n3333 & ~n3334;
  assign n3336 = n3307 & n3313;
  assign n3337 = ~n3183 & n3213;
  assign n3338 = n3306 & n3331;
  assign n3339 = n3315 & n3324;
  assign n3340 = n3315 & n3331;
  assign n3341 = ~n3325 & ~n3340;
  assign n3342 = ~n3339 & n3341;
  assign n3343 = n3269 & n3320;
  assign n3344 = ~n3316 & ~n3343;
  assign n3345 = ~n3332 & n3344;
  assign n3346 = n3342 & n3345;
  assign n3347 = ~n3310 & n3346;
  assign n3348 = ~n3338 & n3347;
  assign n3349 = n3337 & n3348;
  assign n3350 = ~n3336 & ~n3349;
  assign n3351 = ~n3338 & ~n3339;
  assign n3355 = n3320 & n3331;
  assign n3356 = n3308 & n3324;
  assign n3357 = ~n3355 & ~n3356;
  assign n3358 = n3351 & n3357;
  assign n3352 = ~n3321 & ~n3340;
  assign n3353 = n3351 & n3352;
  assign n3354 = ~n3343 & n3353;
  assign n3359 = n3358 ^ n3354;
  assign n3360 = n3359 ^ n3358;
  assign n3361 = n3358 ^ n3183;
  assign n3362 = n3361 ^ n3358;
  assign n3363 = ~n3360 & n3362;
  assign n3364 = n3363 ^ n3358;
  assign n3365 = n3213 & ~n3364;
  assign n3366 = n3365 ^ n3358;
  assign n3367 = n3350 & n3366;
  assign n3368 = n3335 & n3367;
  assign n3369 = n3330 & n3368;
  assign n3370 = ~n3323 & n3369;
  assign n3371 = n3319 & n3370;
  assign n3372 = n3371 ^ n1226;
  assign n3373 = n3372 ^ x224;
  assign n3374 = n2971 & n2982;
  assign n3375 = ~n3002 & ~n3026;
  assign n3376 = n2976 & ~n3375;
  assign n3377 = n2971 & ~n2986;
  assign n3378 = ~n3376 & ~n3377;
  assign n3379 = ~n3374 & n3378;
  assign n3380 = n2973 & n3000;
  assign n3381 = ~n3011 & ~n3380;
  assign n3382 = n2971 & ~n3381;
  assign n3383 = ~n2975 & ~n3014;
  assign n3384 = n3012 & ~n3026;
  assign n3385 = n3383 & n3384;
  assign n3386 = n2983 & n3385;
  assign n3387 = ~n3380 & n3386;
  assign n3388 = n2988 & n3387;
  assign n3389 = ~n3382 & ~n3388;
  assign n3390 = n2979 & n3010;
  assign n3391 = ~n3009 & n3016;
  assign n3392 = ~n3390 & n3391;
  assign n3393 = n2976 & ~n3392;
  assign n3394 = n2983 & ~n3004;
  assign n3395 = ~n3390 & n3394;
  assign n3396 = ~n2975 & n3395;
  assign n3397 = n3007 & ~n3396;
  assign n3398 = ~n3393 & ~n3397;
  assign n3399 = n3389 & n3398;
  assign n3400 = n2978 & n3399;
  assign n3401 = n2970 ^ n2969;
  assign n3402 = n3383 ^ n2970;
  assign n3403 = n3402 ^ n3383;
  assign n3404 = ~n2968 & n3015;
  assign n3405 = n3404 ^ n3383;
  assign n3406 = ~n3403 & n3405;
  assign n3407 = n3406 ^ n3383;
  assign n3408 = ~n3401 & ~n3407;
  assign n3409 = n3400 & ~n3408;
  assign n3410 = n3379 & n3409;
  assign n3411 = n3410 ^ x34;
  assign n3412 = n3411 ^ x178;
  assign n3413 = n2322 ^ x183;
  assign n3414 = n3412 & n3413;
  assign n3415 = n1382 ^ x182;
  assign n3416 = ~n2803 & n2820;
  assign n3417 = n2813 & ~n3222;
  assign n3418 = ~n3416 & ~n3417;
  assign n3419 = n2752 & n2809;
  assign n3420 = ~n2750 & n2826;
  assign n3421 = ~n3419 & ~n3420;
  assign n3422 = n2751 ^ n2750;
  assign n3423 = n2841 & ~n2846;
  assign n3424 = ~n2821 & n3423;
  assign n3425 = ~n3422 & ~n3424;
  assign n3426 = ~n2839 & ~n2861;
  assign n3427 = ~n2815 & ~n2836;
  assign n3428 = ~n2805 & n3427;
  assign n3429 = n3426 & n3428;
  assign n3430 = n2797 ^ n2774;
  assign n3431 = n3430 ^ n2753;
  assign n3432 = ~n2798 & ~n3431;
  assign n3433 = n2805 & n3432;
  assign n3434 = ~n2813 & ~n3433;
  assign n3435 = ~n3429 & ~n3434;
  assign n3436 = ~n3425 & ~n3435;
  assign n3437 = n3421 & n3436;
  assign n3438 = n3418 & n3437;
  assign n3439 = n3217 & n3438;
  assign n3440 = n2812 & n3439;
  assign n3441 = n3440 ^ x18;
  assign n3442 = n3441 ^ x180;
  assign n3443 = n3415 & n3442;
  assign n3444 = n1901 & n1909;
  assign n3445 = n1902 & n1916;
  assign n3446 = ~n3444 & ~n3445;
  assign n3447 = n1717 & n1908;
  assign n3448 = ~n1903 & n1927;
  assign n3449 = ~n3447 & ~n3448;
  assign n3450 = n3446 & n3449;
  assign n3451 = n1915 & n3285;
  assign n3452 = n1940 & ~n1946;
  assign n3453 = ~n1900 & n3452;
  assign n3454 = n1719 & ~n3453;
  assign n3455 = ~n1902 & ~n1915;
  assign n3456 = n1924 & ~n3455;
  assign n3457 = ~n1961 & ~n3456;
  assign n3458 = n1719 & n1945;
  assign n3459 = n1915 & ~n1940;
  assign n3460 = ~n3458 & ~n3459;
  assign n3461 = n1900 & n1915;
  assign n3462 = n1902 & n1941;
  assign n3463 = ~n1909 & ~n1913;
  assign n3464 = n1719 & ~n3463;
  assign n3465 = ~n3462 & ~n3464;
  assign n3466 = ~n3461 & n3465;
  assign n3467 = ~n3282 & n3466;
  assign n3468 = n3278 & n3467;
  assign n3469 = n3460 & n3468;
  assign n3470 = n3457 & n3469;
  assign n3471 = ~n3454 & n3470;
  assign n3472 = ~n3451 & n3471;
  assign n3473 = n3450 & n3472;
  assign n3474 = n1920 & n3473;
  assign n3475 = n3474 ^ x26;
  assign n3476 = n3475 ^ x179;
  assign n3477 = ~n1431 & n1627;
  assign n3478 = n1625 & n1633;
  assign n3479 = ~n1397 & n1657;
  assign n3480 = n1623 & ~n1673;
  assign n3481 = ~n1651 & n3480;
  assign n3482 = ~n1658 & n3481;
  assign n3483 = n1432 & ~n3482;
  assign n3484 = ~n3479 & ~n3483;
  assign n3485 = ~n1554 & n1614;
  assign n3486 = ~n1657 & ~n3485;
  assign n3487 = n1674 & n3486;
  assign n3488 = n1617 & ~n3487;
  assign n3489 = n1652 & ~n1664;
  assign n3490 = ~n1642 & n3489;
  assign n3491 = ~n1636 & ~n2886;
  assign n3492 = n1649 & n3491;
  assign n3493 = ~n3490 & ~n3492;
  assign n3494 = ~n1638 & ~n3493;
  assign n3495 = ~n1663 & ~n3494;
  assign n3496 = ~n3488 & ~n3495;
  assign n3497 = n3484 & n3496;
  assign n3498 = ~n3478 & n3497;
  assign n3499 = ~n3477 & n3498;
  assign n3500 = n1632 & n3499;
  assign n3501 = n2889 & n3500;
  assign n3502 = ~n1616 & n3501;
  assign n3503 = n3502 ^ x10;
  assign n3504 = n3503 ^ x181;
  assign n3505 = ~n3476 & n3504;
  assign n3506 = n3443 & n3505;
  assign n3507 = n3414 & n3506;
  assign n3508 = ~n3412 & n3413;
  assign n3509 = ~n3415 & ~n3442;
  assign n3510 = n3476 & n3504;
  assign n3511 = n3509 & n3510;
  assign n3512 = ~n3476 & ~n3504;
  assign n3513 = n3443 & n3512;
  assign n3514 = ~n3511 & ~n3513;
  assign n3515 = n3508 & ~n3514;
  assign n3516 = ~n3507 & ~n3515;
  assign n3517 = n3476 & ~n3504;
  assign n3518 = ~n3415 & n3517;
  assign n3519 = ~n3415 & n3442;
  assign n3520 = ~n3476 & n3519;
  assign n3521 = ~n3511 & ~n3520;
  assign n3522 = ~n3518 & n3521;
  assign n3523 = n3414 & ~n3522;
  assign n3524 = ~n3476 & n3509;
  assign n3525 = n3510 & n3519;
  assign n3526 = ~n3524 & ~n3525;
  assign n3527 = n3415 & ~n3442;
  assign n3528 = n3505 & n3527;
  assign n3529 = n3517 & n3527;
  assign n3530 = ~n3528 & ~n3529;
  assign n3531 = n3526 & n3530;
  assign n3532 = n3508 & ~n3531;
  assign n3533 = ~n3523 & ~n3532;
  assign n3534 = n3412 & ~n3413;
  assign n3535 = ~n3415 & n3512;
  assign n3536 = n3442 ^ n3415;
  assign n3537 = n3510 ^ n3442;
  assign n3538 = n3537 ^ n3510;
  assign n3539 = n3510 ^ n3504;
  assign n3540 = n3539 ^ n3510;
  assign n3541 = ~n3538 & ~n3540;
  assign n3542 = n3541 ^ n3510;
  assign n3543 = ~n3536 & n3542;
  assign n3544 = n3543 ^ n3510;
  assign n3545 = ~n3535 & ~n3544;
  assign n3546 = ~n3513 & n3545;
  assign n3547 = n3534 & n3546;
  assign n3548 = n3530 & n3547;
  assign n3549 = ~n3412 & ~n3413;
  assign n3550 = ~n3513 & ~n3524;
  assign n3551 = ~n3506 & n3545;
  assign n3552 = n3550 & n3551;
  assign n3553 = n3549 & ~n3552;
  assign n3554 = ~n3548 & ~n3553;
  assign n3555 = n3533 & n3554;
  assign n3556 = n3516 & n3555;
  assign n3557 = n3443 & n3517;
  assign n3558 = n3557 ^ n3412;
  assign n3559 = n3558 ^ n3557;
  assign n3560 = n3557 ^ n3530;
  assign n3561 = n3559 & ~n3560;
  assign n3562 = n3561 ^ n3557;
  assign n3563 = n3413 & n3562;
  assign n3564 = n3556 & ~n3563;
  assign n3565 = n3564 ^ n1069;
  assign n3566 = n3565 ^ x222;
  assign n3567 = n3373 & n3566;
  assign n3568 = ~n2800 & n3226;
  assign n3569 = n2837 & n3568;
  assign n3570 = ~n2861 & n3569;
  assign n3571 = n3570 ^ n2809;
  assign n3572 = n3571 ^ n2809;
  assign n3573 = n2809 ^ n2751;
  assign n3574 = n3573 ^ n2809;
  assign n3575 = ~n3572 & ~n3574;
  assign n3576 = n3575 ^ n2809;
  assign n3577 = n2750 & n3576;
  assign n3578 = n3577 ^ n2809;
  assign n3579 = n2848 & n3428;
  assign n3580 = ~n2821 & n2837;
  assign n3581 = ~n2824 & n3580;
  assign n3582 = ~n2752 & n3581;
  assign n3583 = ~n3579 & ~n3582;
  assign n3584 = n3583 ^ n2751;
  assign n3585 = n3584 ^ n3583;
  assign n3586 = ~n2826 & n3426;
  assign n3587 = ~n2802 & n3586;
  assign n3588 = n3587 ^ n3583;
  assign n3589 = n3588 ^ n3583;
  assign n3590 = n3585 & ~n3589;
  assign n3591 = n3590 ^ n3583;
  assign n3592 = n2750 & n3591;
  assign n3593 = n3592 ^ n3583;
  assign n3594 = ~n3578 & ~n3593;
  assign n3595 = n3220 ^ n2751;
  assign n3596 = n3595 ^ n3220;
  assign n3597 = n3220 ^ n2802;
  assign n3598 = n3597 ^ n3220;
  assign n3599 = n3596 & n3598;
  assign n3600 = n3599 ^ n3220;
  assign n3601 = n3422 & ~n3600;
  assign n3602 = n3601 ^ n3220;
  assign n3603 = n3594 & n3602;
  assign n3604 = n2834 & n3603;
  assign n3605 = n2830 & n3604;
  assign n3606 = n3605 ^ x40;
  assign n3607 = n3606 ^ x163;
  assign n3608 = ~n1896 & ~n1945;
  assign n3609 = n1901 & ~n3608;
  assign n3610 = ~n1900 & n3276;
  assign n3611 = n1719 & ~n3610;
  assign n3612 = ~n3609 & ~n3611;
  assign n3613 = n1903 & n3285;
  assign n3614 = n1915 & n1955;
  assign n3615 = ~n1921 & ~n3285;
  assign n3616 = ~n1900 & n3615;
  assign n3617 = n1902 & ~n3616;
  assign n3618 = ~n1938 & ~n1946;
  assign n3619 = n1901 & ~n3618;
  assign n3620 = ~n3617 & ~n3619;
  assign n3621 = ~n3614 & n3620;
  assign n3622 = n3275 & n3621;
  assign n3623 = n3460 & n3622;
  assign n3624 = n3457 & n3623;
  assign n3625 = ~n3613 & n3624;
  assign n3626 = n3612 & n3625;
  assign n3627 = n1908 ^ n1902;
  assign n3628 = n1902 ^ n1901;
  assign n3629 = n3628 ^ n1901;
  assign n3630 = n1917 ^ n1901;
  assign n3631 = n3629 & n3630;
  assign n3632 = n3631 ^ n1901;
  assign n3633 = n3627 & ~n3632;
  assign n3634 = n3633 ^ n1908;
  assign n3635 = n3626 & ~n3634;
  assign n3636 = n3281 & n3635;
  assign n3637 = ~n1972 & n3636;
  assign n3638 = n3637 ^ x48;
  assign n3639 = n3638 ^ x162;
  assign n3640 = ~n3607 & n3639;
  assign n3651 = n2123 & ~n2128;
  assign n3652 = n2045 & n2128;
  assign n3653 = ~n2114 & ~n3652;
  assign n3654 = ~n2046 & ~n3653;
  assign n3655 = ~n3651 & ~n3654;
  assign n3656 = n2135 & n2151;
  assign n3657 = n2078 & n2122;
  assign n3658 = n2113 ^ n2077;
  assign n3659 = n3658 ^ n2077;
  assign n3660 = n2128 ^ n2077;
  assign n3661 = ~n3659 & n3660;
  assign n3662 = n3661 ^ n2077;
  assign n3663 = ~n2125 & ~n3662;
  assign n3664 = ~n3657 & ~n3663;
  assign n3665 = n2046 & ~n3664;
  assign n3666 = ~n3656 & ~n3665;
  assign n3667 = n3655 & n3666;
  assign n3668 = ~n2139 & n3667;
  assign n3641 = n2140 & n2151;
  assign n3642 = ~n2045 & ~n2128;
  assign n3643 = n3642 ^ n2046;
  assign n3644 = n3643 ^ n3642;
  assign n3645 = ~n2143 & ~n2157;
  assign n3646 = n3645 ^ n3642;
  assign n3647 = ~n3644 & ~n3646;
  assign n3648 = n3647 ^ n3642;
  assign n3649 = ~n3641 & ~n3648;
  assign n3650 = ~n2120 & n3649;
  assign n3669 = n3668 ^ n3650;
  assign n3670 = ~n2009 & n3669;
  assign n3671 = n3670 ^ n3668;
  assign n3672 = ~n2139 & n3671;
  assign n3673 = n3672 ^ x56;
  assign n3674 = n3673 ^ x161;
  assign n3675 = n2747 ^ x164;
  assign n3676 = n3674 & ~n3675;
  assign n3677 = n3640 & n3676;
  assign n3678 = n2927 & n3010;
  assign n3679 = n2971 & n3678;
  assign n3680 = n2975 & n2988;
  assign n3681 = ~n3679 & ~n3680;
  assign n3682 = n3007 & n3387;
  assign n3683 = n3384 & ~n3390;
  assign n3684 = n2971 & ~n3683;
  assign n3685 = n3005 & ~n3011;
  assign n3686 = ~n2975 & n3685;
  assign n3687 = n2976 & ~n3686;
  assign n3688 = ~n3684 & ~n3687;
  assign n3689 = ~n3682 & n3688;
  assign n3690 = n3014 ^ n2988;
  assign n3691 = n2988 ^ n2976;
  assign n3692 = n3691 ^ n2976;
  assign n3693 = ~n3002 & ~n3678;
  assign n3694 = n3394 & n3693;
  assign n3695 = n3694 ^ n2976;
  assign n3696 = n3692 & n3695;
  assign n3697 = n3696 ^ n2976;
  assign n3698 = n3690 & ~n3697;
  assign n3699 = n3698 ^ n3014;
  assign n3700 = n3689 & ~n3699;
  assign n3701 = n3681 & n3700;
  assign n3702 = n3380 ^ n2970;
  assign n3703 = n3702 ^ n3380;
  assign n3704 = n3390 ^ n3380;
  assign n3705 = ~n3703 & n3704;
  assign n3706 = n3705 ^ n3380;
  assign n3707 = n3401 & n3706;
  assign n3708 = n3701 & ~n3707;
  assign n3709 = n3379 & n3708;
  assign n3710 = n3709 ^ x6;
  assign n3711 = n3710 ^ x160;
  assign n3712 = n2914 ^ x165;
  assign n3713 = n3711 & n3712;
  assign n3714 = n3607 & ~n3639;
  assign n3715 = n3676 & n3714;
  assign n3716 = n3713 & n3715;
  assign n3717 = ~n3711 & n3712;
  assign n3718 = n3607 & n3639;
  assign n3719 = ~n3674 & n3675;
  assign n3720 = n3718 & n3719;
  assign n3721 = n3717 & n3720;
  assign n3722 = ~n3711 & ~n3712;
  assign n3723 = n3715 & n3722;
  assign n3724 = ~n3721 & ~n3723;
  assign n3725 = n3640 & n3719;
  assign n3726 = ~n3674 & ~n3675;
  assign n3727 = n3714 & n3726;
  assign n3728 = ~n3725 & ~n3727;
  assign n3729 = n3717 & ~n3728;
  assign n3730 = n3724 & ~n3729;
  assign n3731 = ~n3607 & ~n3639;
  assign n3732 = n3719 & n3731;
  assign n3733 = n3717 & n3732;
  assign n3734 = n3711 & ~n3712;
  assign n3735 = n3727 & n3734;
  assign n3736 = ~n3733 & ~n3735;
  assign n3737 = n3674 & n3675;
  assign n3738 = n3718 & n3737;
  assign n3739 = n3717 & n3738;
  assign n3740 = n3640 & n3726;
  assign n3741 = ~n3725 & ~n3740;
  assign n3742 = n3713 & ~n3741;
  assign n3743 = ~n3739 & ~n3742;
  assign n3744 = ~n3720 & ~n3740;
  assign n3745 = n3734 & ~n3744;
  assign n3746 = n3712 ^ n3711;
  assign n3747 = n3718 & n3726;
  assign n3748 = ~n3732 & ~n3747;
  assign n3749 = ~n3746 & ~n3748;
  assign n3750 = n3714 & n3719;
  assign n3751 = ~n3712 & n3750;
  assign n3752 = n3674 & n3731;
  assign n3753 = ~n3675 & n3752;
  assign n3754 = ~n3738 & ~n3753;
  assign n3755 = n3713 & ~n3754;
  assign n3756 = ~n3751 & ~n3755;
  assign n3757 = ~n3749 & n3756;
  assign n3758 = ~n3745 & n3757;
  assign n3759 = n3640 & n3737;
  assign n3760 = n3676 & n3718;
  assign n3761 = ~n3759 & ~n3760;
  assign n3762 = n3734 ^ n3722;
  assign n3763 = ~n3675 & n3762;
  assign n3764 = n3763 ^ n3734;
  assign n3765 = n3752 & n3764;
  assign n3766 = n3761 & ~n3765;
  assign n3767 = n3766 ^ n3711;
  assign n3768 = n3767 ^ n3766;
  assign n3769 = n3714 & n3737;
  assign n3770 = n3726 & n3731;
  assign n3771 = ~n3769 & ~n3770;
  assign n3772 = n3771 ^ n3766;
  assign n3773 = n3772 ^ n3766;
  assign n3774 = ~n3768 & ~n3773;
  assign n3775 = n3774 ^ n3766;
  assign n3776 = n3712 & ~n3775;
  assign n3777 = n3776 ^ n3766;
  assign n3778 = n3758 & n3777;
  assign n3779 = n3743 & n3778;
  assign n3780 = n3736 & n3779;
  assign n3781 = n3730 & n3780;
  assign n3782 = ~n3716 & n3781;
  assign n3783 = ~n3677 & n3782;
  assign n3784 = n3783 ^ n1145;
  assign n3785 = n3784 ^ x221;
  assign n3786 = n3238 ^ x195;
  assign n3787 = n2169 ^ x190;
  assign n3788 = n3786 & ~n3787;
  assign n3789 = n1687 ^ x191;
  assign n3790 = n3212 ^ x194;
  assign n3791 = n3789 & ~n3790;
  assign n3792 = n2245 & n2272;
  assign n3793 = n2247 & n2265;
  assign n3794 = ~n2259 & n2683;
  assign n3795 = n2267 & ~n3794;
  assign n3796 = ~n3793 & ~n3795;
  assign n3797 = ~n3792 & n3796;
  assign n3798 = n2173 & n2287;
  assign n3799 = ~n2262 & n2272;
  assign n3800 = ~n3798 & ~n3799;
  assign n3801 = ~n2275 & n2295;
  assign n3802 = n2267 & ~n3801;
  assign n3803 = n2272 & n2283;
  assign n3804 = ~n2269 & n2297;
  assign n3805 = n2247 & ~n3804;
  assign n3806 = n2278 & n2683;
  assign n3807 = ~n2277 & ~n2311;
  assign n3808 = n2272 & ~n3807;
  assign n3809 = ~n2173 & ~n3808;
  assign n3810 = ~n3806 & ~n3809;
  assign n3811 = ~n3805 & ~n3810;
  assign n3812 = ~n3803 & n3811;
  assign n3813 = ~n3802 & n3812;
  assign n3814 = n3800 & n3813;
  assign n3815 = n3797 & n3814;
  assign n3816 = n2681 & n3815;
  assign n3817 = n2271 & n3816;
  assign n3818 = n2252 & n3817;
  assign n3819 = n3818 ^ x12;
  assign n3820 = n3819 ^ x193;
  assign n3821 = n2968 & n2976;
  assign n3822 = n2971 & ~n3003;
  assign n3823 = ~n3821 & ~n3822;
  assign n3824 = ~n2968 & ~n3026;
  assign n3825 = n3005 & n3824;
  assign n3826 = ~n2976 & n3825;
  assign n3827 = n3394 ^ n2988;
  assign n3828 = n3824 ^ n2988;
  assign n3829 = n3828 ^ n3824;
  assign n3830 = n3824 ^ n2979;
  assign n3831 = ~n3829 & n3830;
  assign n3832 = n3831 ^ n3824;
  assign n3833 = ~n3827 & ~n3832;
  assign n3834 = n3833 ^ n3394;
  assign n3835 = ~n3826 & ~n3834;
  assign n3836 = ~n3013 & ~n3835;
  assign n3837 = ~n2991 & ~n3836;
  assign n3838 = ~n3001 & n3381;
  assign n3839 = n2986 & n3838;
  assign n3840 = n3839 ^ n3007;
  assign n3841 = n3840 ^ n3839;
  assign n3842 = n3839 ^ n3009;
  assign n3843 = ~n3841 & ~n3842;
  assign n3844 = n3843 ^ n3839;
  assign n3845 = ~n3837 & n3844;
  assign n3846 = n3823 & n3845;
  assign n3847 = n3681 & n3846;
  assign n3848 = ~n3707 & n3847;
  assign n3849 = n3378 & n3848;
  assign n3850 = ~n3408 & n3849;
  assign n3851 = n3850 ^ x20;
  assign n3852 = n3851 ^ x192;
  assign n3853 = ~n3820 & n3852;
  assign n3854 = n3791 & n3853;
  assign n3855 = n3788 & n3854;
  assign n3856 = n3789 & n3790;
  assign n3857 = n3820 & n3852;
  assign n3858 = n3856 & n3857;
  assign n3859 = n3788 & n3858;
  assign n3860 = ~n3786 & n3787;
  assign n3861 = ~n3789 & n3790;
  assign n3862 = ~n3820 & ~n3852;
  assign n3863 = n3861 & n3862;
  assign n3864 = n3860 & n3863;
  assign n3865 = ~n3789 & ~n3790;
  assign n3866 = n3857 & n3865;
  assign n3867 = n3853 & n3861;
  assign n3868 = ~n3866 & ~n3867;
  assign n3869 = n3788 & ~n3868;
  assign n3870 = ~n3864 & ~n3869;
  assign n3871 = n3820 & ~n3852;
  assign n3872 = n3865 & n3871;
  assign n3873 = n3788 & n3872;
  assign n3874 = ~n3786 & ~n3787;
  assign n3875 = n3861 & n3871;
  assign n3876 = n3874 & n3875;
  assign n3877 = ~n3873 & ~n3876;
  assign n3878 = n3787 ^ n3786;
  assign n3879 = n3862 & n3865;
  assign n3880 = ~n3867 & ~n3879;
  assign n3881 = ~n3878 & ~n3880;
  assign n3882 = n3853 & n3856;
  assign n3883 = n3791 & n3862;
  assign n3884 = ~n3882 & ~n3883;
  assign n3885 = ~n3875 & n3884;
  assign n3886 = n3788 & ~n3885;
  assign n3887 = n3857 & n3861;
  assign n3888 = ~n3872 & ~n3887;
  assign n3889 = n3860 & ~n3888;
  assign n3890 = n3791 & n3871;
  assign n3891 = ~n3854 & ~n3858;
  assign n3892 = ~n3890 & n3891;
  assign n3893 = n3874 & ~n3892;
  assign n3894 = n3856 & n3862;
  assign n3895 = ~n3883 & ~n3894;
  assign n3896 = n3791 & n3857;
  assign n3897 = n3856 & n3871;
  assign n3898 = ~n3896 & ~n3897;
  assign n3899 = n3895 & n3898;
  assign n3900 = n3892 & ~n3897;
  assign n3901 = ~n3860 & n3900;
  assign n3902 = ~n3899 & ~n3901;
  assign n3903 = ~n3893 & ~n3902;
  assign n3904 = ~n3786 & ~n3903;
  assign n3905 = ~n3889 & ~n3904;
  assign n3906 = ~n3886 & n3905;
  assign n3907 = ~n3881 & n3906;
  assign n3908 = n3820 ^ n3790;
  assign n3909 = n3908 ^ n3852;
  assign n3910 = ~n3789 & ~n3852;
  assign n3911 = n3909 & n3910;
  assign n3912 = n3911 ^ n3909;
  assign n3913 = n3912 ^ n3866;
  assign n3914 = n3913 ^ n3866;
  assign n3915 = n3866 ^ n3787;
  assign n3916 = n3915 ^ n3866;
  assign n3917 = n3914 & n3916;
  assign n3918 = n3917 ^ n3866;
  assign n3919 = n3786 & n3918;
  assign n3920 = n3919 ^ n3866;
  assign n3921 = n3907 & ~n3920;
  assign n3922 = n3877 & n3921;
  assign n3923 = n3870 & n3922;
  assign n3924 = ~n3859 & n3923;
  assign n3925 = ~n3855 & n3924;
  assign n3926 = n3925 ^ n1309;
  assign n3927 = n3926 ^ x223;
  assign n3928 = ~n3785 & n3927;
  assign n3929 = n3567 & n3928;
  assign n3930 = n3148 & n3929;
  assign n3931 = ~n3373 & ~n3566;
  assign n3932 = ~n3785 & ~n3927;
  assign n3933 = n3931 & n3932;
  assign n3934 = n3148 & n3933;
  assign n3935 = ~n2669 & n3147;
  assign n3936 = n3785 & n3927;
  assign n3937 = n3567 & n3936;
  assign n3938 = n3931 & n3936;
  assign n3939 = ~n3937 & ~n3938;
  assign n3940 = n3935 & ~n3939;
  assign n3941 = ~n3934 & ~n3940;
  assign n3942 = ~n3930 & n3941;
  assign n3943 = n3373 & ~n3566;
  assign n3944 = n3928 & n3943;
  assign n3945 = n3148 & n3944;
  assign n3946 = n3785 & ~n3927;
  assign n3947 = n3931 & n3946;
  assign n3948 = n3935 & n3947;
  assign n3949 = ~n3945 & ~n3948;
  assign n3950 = n2669 & ~n3147;
  assign n3951 = n3928 & n3931;
  assign n3952 = n3950 & n3951;
  assign n3953 = ~n2669 & ~n3147;
  assign n3954 = n3567 & n3932;
  assign n3955 = n3953 & n3954;
  assign n3956 = ~n3952 & ~n3955;
  assign n3957 = n3949 & n3956;
  assign n3958 = n3567 & n3946;
  assign n3959 = n3953 & n3958;
  assign n3960 = ~n3951 & ~n3954;
  assign n3961 = n3935 & ~n3960;
  assign n3962 = ~n3373 & n3566;
  assign n3963 = n3946 & n3962;
  assign n3964 = n3943 & n3946;
  assign n3965 = ~n3963 & ~n3964;
  assign n3966 = n3950 & ~n3965;
  assign n3967 = ~n3961 & ~n3966;
  assign n3968 = n3932 & n3962;
  assign n3969 = n3935 & n3968;
  assign n3970 = n3932 & n3943;
  assign n3971 = n3935 & n3970;
  assign n3972 = n3148 & n3958;
  assign n3973 = ~n3971 & ~n3972;
  assign n3974 = ~n3969 & n3973;
  assign n3975 = ~n3939 & n3950;
  assign n3976 = ~n3935 & ~n3950;
  assign n3977 = n3936 & n3962;
  assign n3978 = n3936 & n3943;
  assign n3979 = ~n3977 & ~n3978;
  assign n3980 = ~n3947 & n3979;
  assign n3981 = n3976 & ~n3980;
  assign n3982 = ~n3929 & ~n3970;
  assign n3983 = ~n3147 & ~n3982;
  assign n3984 = ~n3981 & ~n3983;
  assign n3985 = ~n3975 & n3984;
  assign n3986 = n3974 & n3985;
  assign n3987 = n3967 & n3986;
  assign n3988 = ~n3959 & n3987;
  assign n3989 = n3976 ^ n3968;
  assign n3990 = n3989 ^ n3968;
  assign n3991 = n3928 & n3962;
  assign n3992 = n3991 ^ n3968;
  assign n3993 = ~n3990 & n3992;
  assign n3994 = n3993 ^ n3968;
  assign n3995 = n3988 & ~n3994;
  assign n3996 = n3957 & n3995;
  assign n3997 = n3942 & n3996;
  assign n3998 = n3997 ^ n3212;
  assign n3999 = n3998 ^ x292;
  assign n4000 = ~n1383 & n2610;
  assign n4001 = n1689 & ~n2618;
  assign n4002 = ~n4000 & ~n4001;
  assign n4003 = ~n2327 & ~n2625;
  assign n4004 = n2643 & ~n4003;
  assign n4005 = n2609 & ~n2630;
  assign n4006 = ~n4004 & ~n4005;
  assign n4007 = n4002 & n4006;
  assign n4008 = n2617 & n2625;
  assign n4009 = ~n2615 & ~n2644;
  assign n4010 = ~n2650 & n4009;
  assign n4011 = n2327 & ~n4010;
  assign n4012 = n2325 & ~n2592;
  assign n4013 = ~n2598 & ~n2636;
  assign n4014 = ~n4012 & n4013;
  assign n4015 = ~n2627 & n4014;
  assign n4016 = n2625 & ~n4015;
  assign n4017 = ~n2595 & n2618;
  assign n4018 = ~n2643 & n4017;
  assign n4019 = n2609 & ~n4018;
  assign n4020 = ~n4016 & ~n4019;
  assign n4021 = ~n2327 & ~n2633;
  assign n4022 = ~n2638 & ~n4021;
  assign n4023 = ~n2606 & ~n2628;
  assign n4024 = n4023 ^ n2595;
  assign n4025 = n2327 ^ n1689;
  assign n4026 = n4023 ^ n2327;
  assign n4027 = n4026 ^ n2327;
  assign n4028 = ~n4025 & ~n4027;
  assign n4029 = n4028 ^ n2327;
  assign n4030 = ~n4024 & ~n4029;
  assign n4031 = n4030 ^ n2595;
  assign n4032 = ~n4012 & ~n4031;
  assign n4033 = ~n2607 & ~n4032;
  assign n4034 = ~n4022 & ~n4033;
  assign n4035 = n4020 & n4034;
  assign n4036 = ~n4011 & n4035;
  assign n4037 = ~n4008 & n4036;
  assign n4038 = n4007 & n4037;
  assign n4039 = ~n2601 & ~n2627;
  assign n4040 = n4039 ^ n2612;
  assign n4041 = n4040 ^ n2612;
  assign n4042 = n2612 ^ n1688;
  assign n4043 = n4042 ^ n2612;
  assign n4044 = ~n4041 & n4043;
  assign n4045 = n4044 ^ n2612;
  assign n4046 = n1383 & n4045;
  assign n4047 = n4046 ^ n2612;
  assign n4048 = n4038 & ~n4047;
  assign n4049 = n4048 ^ n2388;
  assign n4050 = n4049 ^ x243;
  assign n4051 = n3304 ^ x202;
  assign n4052 = n3673 ^ x207;
  assign n4053 = ~n4051 & n4052;
  assign n4054 = ~n2255 & ~n2283;
  assign n4055 = ~n2286 & n4054;
  assign n4056 = n2267 & ~n4055;
  assign n4057 = ~n2265 & n2278;
  assign n4058 = n2272 & ~n4057;
  assign n4059 = n2272 & n2287;
  assign n4060 = n2247 & ~n3807;
  assign n4061 = ~n2250 & n2288;
  assign n4062 = ~n2275 & n4061;
  assign n4063 = n2173 & ~n4062;
  assign n4064 = ~n4060 & ~n4063;
  assign n4065 = ~n4059 & n4064;
  assign n4066 = ~n2291 & n4065;
  assign n4067 = ~n4058 & n4066;
  assign n4068 = ~n4056 & n4067;
  assign n4069 = n3797 & n4068;
  assign n4070 = n2680 & n4069;
  assign n4071 = n2677 & n4070;
  assign n4072 = n2264 & n4071;
  assign n4073 = n2674 & n4072;
  assign n4074 = n4073 ^ x14;
  assign n4075 = n4074 ^ x205;
  assign n4076 = n3182 ^ x203;
  assign n4077 = n4075 & n4076;
  assign n4078 = n3710 ^ x206;
  assign n4079 = ~n1319 & ~n3044;
  assign n4080 = n1321 & ~n3053;
  assign n4081 = ~n4079 & ~n4080;
  assign n4082 = n1006 & n1326;
  assign n4083 = ~n1316 & n1366;
  assign n4084 = ~n1338 & n4083;
  assign n4085 = n1318 & ~n4084;
  assign n4086 = ~n4082 & ~n4085;
  assign n4087 = n1311 ^ n1070;
  assign n4088 = ~n1146 & n4087;
  assign n4089 = n1317 & n4088;
  assign n4090 = n3052 ^ n1343;
  assign n4091 = n3052 ^ n1005;
  assign n4092 = ~n1325 & ~n4091;
  assign n4093 = n4092 ^ n1005;
  assign n4094 = ~n4090 & ~n4093;
  assign n4095 = n4094 ^ n1343;
  assign n4096 = ~n1330 & ~n4095;
  assign n4097 = ~n1323 & n4096;
  assign n4098 = n1319 & ~n4097;
  assign n4099 = ~n4089 & ~n4098;
  assign n4100 = n4086 & n4099;
  assign n4101 = n4081 & n4100;
  assign n4102 = n3042 & n4101;
  assign n4103 = ~n1313 & n4102;
  assign n4104 = ~n1360 & n4103;
  assign n4105 = n4104 ^ x22;
  assign n4106 = n4105 ^ x204;
  assign n4107 = ~n4078 & n4106;
  assign n4108 = n4077 & n4107;
  assign n4109 = ~n4075 & n4076;
  assign n4110 = n4078 & n4106;
  assign n4111 = n4109 & n4110;
  assign n4112 = ~n4078 & ~n4106;
  assign n4113 = n4109 & n4112;
  assign n4114 = ~n4111 & ~n4113;
  assign n4115 = ~n4108 & n4114;
  assign n4116 = n4053 & ~n4115;
  assign n4117 = n4051 & n4052;
  assign n4118 = n4078 & ~n4106;
  assign n4119 = n4109 & n4118;
  assign n4120 = n4117 & n4119;
  assign n4121 = n4051 & ~n4052;
  assign n4122 = ~n4114 & n4121;
  assign n4123 = ~n4120 & ~n4122;
  assign n4124 = n4052 ^ n4051;
  assign n4125 = n4075 & ~n4076;
  assign n4126 = n4107 & n4125;
  assign n4127 = ~n4124 & n4126;
  assign n4128 = ~n4075 & ~n4076;
  assign n4129 = n4110 & n4128;
  assign n4130 = n4112 & n4128;
  assign n4131 = ~n4129 & ~n4130;
  assign n4132 = n4121 & ~n4131;
  assign n4133 = ~n4127 & ~n4132;
  assign n4134 = n4077 & n4112;
  assign n4135 = n4121 & n4134;
  assign n4136 = n4077 & n4110;
  assign n4137 = n4118 & n4128;
  assign n4138 = ~n4134 & ~n4137;
  assign n4139 = ~n4136 & n4138;
  assign n4140 = ~n4126 & n4139;
  assign n4141 = ~n4129 & n4140;
  assign n4142 = n4053 & ~n4141;
  assign n4143 = ~n4135 & ~n4142;
  assign n4144 = n4110 & n4125;
  assign n4145 = n4107 & n4128;
  assign n4146 = n4077 & n4118;
  assign n4147 = ~n4145 & ~n4146;
  assign n4148 = ~n4144 & n4147;
  assign n4149 = n4051 & ~n4148;
  assign n4150 = n4107 & n4109;
  assign n4151 = ~n4130 & ~n4150;
  assign n4152 = ~n4124 & ~n4151;
  assign n4153 = ~n4051 & ~n4052;
  assign n4154 = ~n4119 & n4139;
  assign n4155 = n4153 & ~n4154;
  assign n4156 = ~n4152 & ~n4155;
  assign n4157 = ~n4149 & n4156;
  assign n4158 = n4143 & n4157;
  assign n4159 = n4133 & n4158;
  assign n4160 = n4123 & n4159;
  assign n4161 = ~n4116 & n4160;
  assign n4162 = n4118 & n4125;
  assign n4163 = n4162 ^ n4052;
  assign n4164 = n4163 ^ n4162;
  assign n4165 = n4112 & n4125;
  assign n4166 = n4165 ^ n4162;
  assign n4167 = n4164 & n4166;
  assign n4168 = n4167 ^ n4162;
  assign n4169 = ~n4124 & n4168;
  assign n4170 = n4161 & ~n4169;
  assign n4171 = n4170 ^ n2422;
  assign n4172 = n4171 ^ x239;
  assign n4173 = n2873 ^ x172;
  assign n4174 = n3475 ^ x177;
  assign n4175 = n4173 & ~n4174;
  assign n4176 = ~n4173 & n4174;
  assign n4177 = ~n4175 & ~n4176;
  assign n4178 = n2701 ^ x173;
  assign n4179 = ~n2139 & n3650;
  assign n4180 = n4179 ^ n3668;
  assign n4181 = n2009 & ~n4180;
  assign n4182 = n4181 ^ n3668;
  assign n4183 = n4182 ^ x50;
  assign n4184 = n4183 ^ x174;
  assign n4185 = n4178 & ~n4184;
  assign n4186 = n3411 ^ x176;
  assign n4187 = n2532 & n2543;
  assign n4188 = n2390 & n2546;
  assign n4189 = ~n4187 & ~n4188;
  assign n4190 = n2364 & n2568;
  assign n4191 = ~n2534 & n2558;
  assign n4192 = n2557 & ~n2712;
  assign n4193 = ~n2389 & n2567;
  assign n4194 = ~n2555 & n2564;
  assign n4195 = ~n2553 & n4194;
  assign n4196 = n2533 & ~n4195;
  assign n4197 = ~n4193 & ~n4196;
  assign n4198 = ~n4192 & n4197;
  assign n4199 = n2532 ^ n2516;
  assign n4200 = n4199 ^ n2532;
  assign n4201 = n2532 ^ n2477;
  assign n4202 = n4200 & ~n4201;
  assign n4203 = n4202 ^ n2532;
  assign n4204 = n2524 & n4203;
  assign n4205 = ~n2546 & ~n4204;
  assign n4206 = n4205 ^ n2389;
  assign n4207 = n4206 ^ n4205;
  assign n4208 = n4205 ^ n2568;
  assign n4209 = n4208 ^ n4205;
  assign n4210 = n4207 & n4209;
  assign n4211 = n4210 ^ n4205;
  assign n4212 = ~n2364 & ~n4211;
  assign n4213 = n4212 ^ n4205;
  assign n4214 = n4198 & n4213;
  assign n4215 = n3151 & n4214;
  assign n4216 = ~n2523 & n4215;
  assign n4217 = ~n4191 & n4216;
  assign n4218 = ~n4190 & n4217;
  assign n4219 = n4189 & n4218;
  assign n4220 = n3155 & n4219;
  assign n4221 = n2706 & n4220;
  assign n4222 = n4221 ^ x42;
  assign n4223 = n4222 ^ x175;
  assign n4224 = n4186 & ~n4223;
  assign n4225 = n4185 & n4224;
  assign n4226 = ~n4177 & n4225;
  assign n4227 = ~n4173 & ~n4174;
  assign n4228 = n4186 & n4223;
  assign n4229 = n4185 & n4228;
  assign n4230 = n4178 & n4184;
  assign n4231 = ~n4186 & n4223;
  assign n4232 = n4230 & n4231;
  assign n4233 = ~n4229 & ~n4232;
  assign n4234 = n4227 & ~n4233;
  assign n4235 = ~n4226 & ~n4234;
  assign n4236 = n4173 & n4174;
  assign n4237 = ~n4178 & n4184;
  assign n4238 = n4231 & n4237;
  assign n4239 = n4236 & n4238;
  assign n4240 = n4174 ^ n4173;
  assign n4241 = n4185 & n4231;
  assign n4242 = n4241 ^ n4174;
  assign n4243 = n4242 ^ n4241;
  assign n4244 = n4228 & n4230;
  assign n4245 = n4244 ^ n4241;
  assign n4246 = n4243 & n4245;
  assign n4247 = n4246 ^ n4241;
  assign n4248 = n4240 & n4247;
  assign n4249 = ~n4239 & ~n4248;
  assign n4250 = n4224 & n4230;
  assign n4251 = ~n4186 & ~n4223;
  assign n4252 = n4185 & n4251;
  assign n4253 = ~n4250 & ~n4252;
  assign n4254 = n4227 & ~n4253;
  assign n4255 = n4175 & n4244;
  assign n4256 = n4176 & n4241;
  assign n4257 = n4228 & n4237;
  assign n4258 = ~n4178 & ~n4184;
  assign n4259 = n4228 & n4258;
  assign n4260 = n4251 & n4258;
  assign n4261 = ~n4259 & ~n4260;
  assign n4262 = ~n4257 & n4261;
  assign n4263 = n4236 & ~n4262;
  assign n4264 = n4230 & n4251;
  assign n4271 = ~n4257 & ~n4259;
  assign n4265 = n4224 & n4237;
  assign n4266 = ~n4238 & ~n4265;
  assign n4267 = n4231 & n4258;
  assign n4268 = n4224 & n4258;
  assign n4269 = ~n4267 & ~n4268;
  assign n4270 = n4266 & n4269;
  assign n4272 = n4271 ^ n4270;
  assign n4273 = n4270 ^ n4175;
  assign n4274 = n4273 ^ n4175;
  assign n4275 = ~n4176 & n4266;
  assign n4276 = n4275 ^ n4175;
  assign n4277 = ~n4274 & n4276;
  assign n4278 = n4277 ^ n4175;
  assign n4279 = n4272 & ~n4278;
  assign n4280 = n4279 ^ n4271;
  assign n4281 = ~n4264 & n4280;
  assign n4282 = n4281 ^ n4177;
  assign n4283 = n4282 ^ n4281;
  assign n4284 = n4237 & n4251;
  assign n4286 = n4261 & ~n4265;
  assign n4285 = ~n4241 & n4253;
  assign n4287 = n4286 ^ n4285;
  assign n4288 = n4285 ^ n4227;
  assign n4289 = n4288 ^ n4227;
  assign n4290 = n4236 ^ n4227;
  assign n4291 = ~n4289 & ~n4290;
  assign n4292 = n4291 ^ n4227;
  assign n4293 = n4287 & ~n4292;
  assign n4294 = n4293 ^ n4286;
  assign n4295 = ~n4284 & n4294;
  assign n4296 = n4295 ^ n4281;
  assign n4297 = n4283 & n4296;
  assign n4298 = n4297 ^ n4281;
  assign n4299 = ~n4263 & n4298;
  assign n4300 = ~n4256 & n4299;
  assign n4301 = ~n4255 & n4300;
  assign n4302 = ~n4254 & n4301;
  assign n4303 = n4249 & n4302;
  assign n4304 = n4235 & n4303;
  assign n4305 = n4304 ^ n2476;
  assign n4306 = n4305 ^ x242;
  assign n4307 = ~n4172 & n4306;
  assign n4308 = n3337 & ~n3357;
  assign n4309 = ~n3332 & ~n3338;
  assign n4310 = n3213 & ~n4309;
  assign n4311 = n3320 & n3324;
  assign n4312 = n3269 & n3315;
  assign n4313 = ~n3314 & ~n4312;
  assign n4314 = ~n4311 & n4313;
  assign n4315 = ~n3339 & n4314;
  assign n4316 = n3214 & ~n4315;
  assign n4317 = n3342 & ~n4312;
  assign n4318 = ~n3355 & n4317;
  assign n4319 = ~n3307 & n4318;
  assign n4320 = n3322 & ~n4319;
  assign n4321 = ~n4316 & ~n4320;
  assign n4322 = n3352 & ~n3355;
  assign n4323 = n3313 & ~n4322;
  assign n4324 = n3213 ^ n3183;
  assign n4325 = ~n3308 & ~n3337;
  assign n4326 = n3310 & n3313;
  assign n4327 = ~n3328 & ~n4326;
  assign n4328 = ~n3321 & n4327;
  assign n4329 = ~n3316 & n4328;
  assign n4330 = ~n4325 & ~n4329;
  assign n4331 = n4324 & n4330;
  assign n4332 = ~n4323 & ~n4331;
  assign n4333 = n4321 & n4332;
  assign n4334 = n3319 & n4333;
  assign n4335 = ~n4310 & n4334;
  assign n4336 = ~n4308 & n4335;
  assign n4337 = n3335 & n4336;
  assign n4338 = ~n3323 & n4337;
  assign n4339 = n4338 ^ n2515;
  assign n4340 = n4339 ^ x240;
  assign n4341 = n3722 & n3732;
  assign n4342 = n3717 & n3760;
  assign n4343 = ~n4341 & ~n4342;
  assign n4344 = n3717 & n3759;
  assign n4345 = n3713 & n3720;
  assign n4346 = ~n3725 & ~n3738;
  assign n4347 = n3722 & ~n4346;
  assign n4348 = ~n4345 & ~n4347;
  assign n4349 = ~n4344 & n4348;
  assign n4350 = ~n3747 & ~n3750;
  assign n4351 = n3734 & ~n4350;
  assign n4352 = n3732 & n3734;
  assign n4353 = n3675 & n3752;
  assign n4354 = ~n3677 & ~n4353;
  assign n4355 = ~n3760 & n4354;
  assign n4356 = n3722 & ~n4355;
  assign n4357 = ~n4352 & ~n4356;
  assign n4358 = n3713 & n3747;
  assign n4359 = ~n3740 & n3754;
  assign n4360 = n3717 & ~n4359;
  assign n4361 = ~n4358 & ~n4360;
  assign n4362 = ~n3750 & ~n3770;
  assign n4363 = ~n3746 & ~n4362;
  assign n4364 = n3759 ^ n3711;
  assign n4367 = ~n3738 & ~n3740;
  assign n4365 = ~n3677 & ~n3769;
  assign n4366 = ~n3753 & n4365;
  assign n4368 = n4367 ^ n4366;
  assign n4369 = n4367 ^ n3712;
  assign n4370 = n4369 ^ n4367;
  assign n4371 = n4368 & ~n4370;
  assign n4372 = n4371 ^ n4367;
  assign n4373 = n4372 ^ n3759;
  assign n4374 = ~n4364 & ~n4373;
  assign n4375 = n4374 ^ n4371;
  assign n4376 = n4375 ^ n4367;
  assign n4377 = n4376 ^ n3711;
  assign n4378 = ~n3759 & n4377;
  assign n4379 = n4378 ^ n3759;
  assign n4380 = n4379 ^ n3711;
  assign n4381 = ~n4363 & n4380;
  assign n4382 = n4361 & n4381;
  assign n4383 = n4357 & n4382;
  assign n4384 = ~n4351 & n4383;
  assign n4385 = n3736 & n4384;
  assign n4386 = ~n3729 & n4385;
  assign n4387 = n4349 & n4386;
  assign n4388 = ~n3716 & n4387;
  assign n4389 = n4343 & n4388;
  assign n4390 = n4389 ^ n2447;
  assign n4391 = n4390 ^ x241;
  assign n4392 = n4340 & ~n4391;
  assign n4393 = n4307 & n4392;
  assign n4394 = ~n4050 & n4393;
  assign n4395 = ~n3509 & n3510;
  assign n4396 = ~n3443 & n3512;
  assign n4397 = ~n4395 & ~n4396;
  assign n4398 = ~n3528 & n4397;
  assign n4399 = ~n3557 & n4398;
  assign n4400 = n3549 & ~n4399;
  assign n4401 = n3443 & n3510;
  assign n4402 = n3517 & n3519;
  assign n4403 = ~n4401 & ~n4402;
  assign n4404 = ~n3528 & n4403;
  assign n4405 = n3504 ^ n3442;
  assign n4410 = n4405 ^ n3442;
  assign n4407 = n4405 ^ n3476;
  assign n4406 = n4405 ^ n3415;
  assign n4408 = n4407 ^ n4406;
  assign n4409 = n4408 ^ n3442;
  assign n4411 = n4410 ^ n4409;
  assign n4412 = n4407 ^ n4405;
  assign n4413 = n4412 ^ n3442;
  assign n4414 = n4413 ^ n3442;
  assign n4415 = ~n4408 & n4414;
  assign n4416 = n4415 ^ n4408;
  assign n4417 = n4413 & ~n4416;
  assign n4418 = n4417 ^ n3442;
  assign n4419 = n4411 & n4418;
  assign n4420 = n4419 ^ n4415;
  assign n4421 = n4420 ^ n3442;
  assign n4422 = n4421 ^ n4410;
  assign n4423 = n4404 & n4422;
  assign n4424 = n3534 & n4423;
  assign n4425 = ~n4400 & ~n4424;
  assign n4426 = n3550 & n4403;
  assign n4427 = n3414 & ~n4426;
  assign n4428 = n3508 & ~n4422;
  assign n4429 = ~n4427 & ~n4428;
  assign n4430 = n4425 & n4429;
  assign n4431 = n3516 & n4430;
  assign n4432 = ~n3563 & n4431;
  assign n4433 = n4432 ^ n2363;
  assign n4434 = n4433 ^ x238;
  assign n4435 = ~n4050 & ~n4434;
  assign n4436 = ~n4340 & ~n4391;
  assign n4437 = n4307 & n4436;
  assign n4438 = ~n4172 & ~n4306;
  assign n4439 = n4392 & n4438;
  assign n4440 = ~n4437 & ~n4439;
  assign n4441 = n4435 & ~n4440;
  assign n4442 = ~n4394 & ~n4441;
  assign n4443 = n4050 & n4434;
  assign n4444 = ~n4435 & ~n4443;
  assign n4445 = ~n4340 & n4391;
  assign n4446 = n4438 & n4445;
  assign n4447 = ~n4444 & n4446;
  assign n4448 = n4050 & ~n4434;
  assign n4449 = n4340 & n4391;
  assign n4450 = n4172 & n4306;
  assign n4451 = n4449 & n4450;
  assign n4452 = n4392 & n4450;
  assign n4453 = n4172 & ~n4306;
  assign n4454 = n4340 & n4453;
  assign n4455 = ~n4452 & ~n4454;
  assign n4456 = ~n4451 & n4455;
  assign n4457 = n4448 & ~n4456;
  assign n4458 = ~n4447 & ~n4457;
  assign n4459 = n4442 & n4458;
  assign n4460 = n4307 & n4449;
  assign n4461 = ~n4439 & ~n4460;
  assign n4462 = ~n4437 & n4461;
  assign n4463 = n4443 & ~n4462;
  assign n4464 = ~n4050 & n4434;
  assign n4465 = n4436 & n4438;
  assign n4466 = n4461 & ~n4465;
  assign n4467 = n4464 & ~n4466;
  assign n4468 = n4436 & n4453;
  assign n4469 = n4445 & n4453;
  assign n4470 = ~n4451 & ~n4469;
  assign n4471 = ~n4460 & n4470;
  assign n4472 = ~n4468 & n4471;
  assign n4473 = n4435 & ~n4472;
  assign n4474 = n4436 & n4450;
  assign n4475 = n4438 & n4449;
  assign n4476 = n4307 & n4445;
  assign n4477 = ~n4465 & ~n4476;
  assign n4478 = ~n4475 & n4477;
  assign n4479 = ~n4474 & n4478;
  assign n4480 = n4448 & ~n4479;
  assign n4481 = n4464 ^ n4443;
  assign n4486 = n4445 & n4450;
  assign n4487 = ~n4454 & ~n4486;
  assign n4488 = ~n4474 & n4487;
  assign n4482 = n4449 & n4453;
  assign n4483 = ~n4452 & ~n4469;
  assign n4484 = ~n4482 & n4483;
  assign n4485 = ~n4468 & n4484;
  assign n4489 = n4488 ^ n4485;
  assign n4490 = n4488 ^ n4464;
  assign n4491 = n4490 ^ n4488;
  assign n4492 = ~n4489 & ~n4491;
  assign n4493 = n4492 ^ n4488;
  assign n4494 = n4481 & ~n4493;
  assign n4495 = n4494 ^ n4443;
  assign n4496 = ~n4480 & ~n4495;
  assign n4497 = ~n4473 & n4496;
  assign n4498 = ~n4467 & n4497;
  assign n4499 = ~n4463 & n4498;
  assign n4500 = n4459 & n4499;
  assign n4501 = n4500 ^ n3182;
  assign n4502 = n4501 ^ x297;
  assign n4503 = n3999 & n4502;
  assign n4504 = n3508 & n3552;
  assign n4505 = n3414 & ~n3546;
  assign n4506 = ~n4504 & ~n4505;
  assign n4507 = ~n3522 & n3534;
  assign n4508 = ~n3415 & n3510;
  assign n4509 = n3550 & ~n4508;
  assign n4510 = n3549 & ~n4509;
  assign n4511 = ~n4507 & ~n4510;
  assign n4512 = n4506 & n4511;
  assign n4513 = n3506 ^ n3412;
  assign n4514 = n4513 ^ n3506;
  assign n4515 = n3557 ^ n3506;
  assign n4516 = ~n4514 & n4515;
  assign n4517 = n4516 ^ n3506;
  assign n4518 = ~n3413 & n4517;
  assign n4519 = n4512 & ~n4518;
  assign n4520 = n3530 & n4519;
  assign n4521 = n4520 ^ n1396;
  assign n4522 = n4521 ^ x255;
  assign n4523 = n3072 & n3094;
  assign n4524 = n2749 & n3116;
  assign n4525 = ~n4523 & ~n4524;
  assign n4526 = n2749 & n3123;
  assign n4527 = n3076 ^ n2748;
  assign n4528 = n4527 ^ n3076;
  assign n4529 = n3106 ^ n3076;
  assign n4530 = ~n4528 & n4529;
  assign n4531 = n4530 ^ n3076;
  assign n4532 = ~n3129 & n4531;
  assign n4533 = ~n4526 & ~n4532;
  assign n4534 = ~n3087 & ~n3130;
  assign n4535 = ~n3114 & ~n4534;
  assign n4536 = n3098 & n3118;
  assign n4537 = ~n3109 & n4536;
  assign n4538 = n2749 & ~n4537;
  assign n4539 = ~n3097 & n3119;
  assign n4540 = n3074 & ~n4539;
  assign n4541 = ~n4538 & ~n4540;
  assign n4542 = ~n4535 & n4541;
  assign n4543 = ~n3085 & ~n3115;
  assign n4544 = ~n3106 & n4543;
  assign n4545 = n3078 & ~n4544;
  assign n4546 = n3034 ^ n2874;
  assign n4547 = n4546 ^ n2874;
  assign n4548 = n3070 ^ n2874;
  assign n4549 = n4548 ^ n2874;
  assign n4550 = n4547 & n4549;
  assign n4551 = n4550 ^ n2874;
  assign n4552 = n2915 & ~n4551;
  assign n4553 = n4552 ^ n4546;
  assign n4554 = n3094 & ~n4553;
  assign n4555 = ~n4545 & ~n4554;
  assign n4556 = n4542 & n4555;
  assign n4557 = n3083 & n4556;
  assign n4558 = n4533 & n4557;
  assign n4559 = ~n3110 & n4558;
  assign n4560 = ~n3112 & n4559;
  assign n4561 = n4525 & n4560;
  assign n4562 = n4561 ^ n1430;
  assign n4563 = n4562 ^ x250;
  assign n4564 = n4522 & n4563;
  assign n4565 = n3324 & n3327;
  assign n4566 = n3213 & n4565;
  assign n4567 = n3328 & n4324;
  assign n4568 = ~n4566 & ~n4567;
  assign n4569 = ~n3314 & n3351;
  assign n4570 = n3337 & ~n4569;
  assign n4571 = n3313 & ~n3342;
  assign n4572 = ~n4570 & ~n4571;
  assign n4573 = n4568 & n4572;
  assign n4574 = n3214 & ~n3345;
  assign n4575 = n3322 & n3348;
  assign n4576 = ~n4574 & ~n4575;
  assign n4577 = n4573 & n4576;
  assign n4578 = ~n3326 & n4577;
  assign n4579 = n3338 ^ n3213;
  assign n4580 = n4579 ^ n3338;
  assign n4581 = n3338 ^ n3310;
  assign n4582 = n4580 & n4581;
  assign n4583 = n4582 ^ n3338;
  assign n4584 = n4324 & n4583;
  assign n4585 = n4578 & ~n4584;
  assign n4586 = n3319 & n4585;
  assign n4587 = n4586 ^ n1579;
  assign n4588 = n4587 ^ x254;
  assign n4589 = ~n3875 & ~n3879;
  assign n4590 = n3874 & ~n4589;
  assign n4591 = n3870 & ~n4590;
  assign n4592 = ~n3854 & ~n3866;
  assign n4593 = n3898 & n4592;
  assign n4594 = ~n3875 & n4593;
  assign n4595 = n3860 & ~n4594;
  assign n4596 = ~n3863 & n3884;
  assign n4597 = ~n3858 & n4596;
  assign n4598 = n3874 & ~n4597;
  assign n4599 = ~n4595 & ~n4598;
  assign n4600 = ~n3878 & n3890;
  assign n4601 = ~n3894 & ~n3896;
  assign n4602 = ~n3890 & n4601;
  assign n4603 = n4589 & n4602;
  assign n4604 = n3788 & ~n4603;
  assign n4605 = n3786 & n3787;
  assign n4606 = n3853 & n3865;
  assign n4607 = n3895 & ~n4606;
  assign n4608 = ~n3882 & ~n3897;
  assign n4609 = ~n3887 & n4608;
  assign n4610 = n4607 & n4609;
  assign n4611 = ~n3872 & n4610;
  assign n4612 = n4605 & ~n4611;
  assign n4613 = ~n4604 & ~n4612;
  assign n4614 = ~n4600 & n4613;
  assign n4615 = n4599 & n4614;
  assign n4616 = n4606 ^ n3787;
  assign n4617 = n4616 ^ n4606;
  assign n4618 = n4606 ^ n3880;
  assign n4619 = n4617 & ~n4618;
  assign n4620 = n4619 ^ n4606;
  assign n4621 = ~n3786 & n4620;
  assign n4622 = n4615 & ~n4621;
  assign n4623 = n4591 & n4622;
  assign n4624 = ~n3855 & n4623;
  assign n4625 = n4624 ^ n1612;
  assign n4626 = n4625 ^ x251;
  assign n4627 = n4588 & ~n4626;
  assign n4628 = n4176 & n4260;
  assign n4629 = n4175 & n4265;
  assign n4630 = ~n4628 & ~n4629;
  assign n4631 = n4236 & ~n4269;
  assign n4632 = n4630 & ~n4631;
  assign n4633 = ~n4229 & ~n4244;
  assign n4634 = ~n4252 & n4633;
  assign n4635 = n4175 & ~n4634;
  assign n4636 = n4175 & ~n4261;
  assign n4637 = n4253 & ~n4257;
  assign n4638 = n4236 & ~n4637;
  assign n4639 = ~n4636 & ~n4638;
  assign n4640 = n4233 & ~n4260;
  assign n4641 = n4177 & ~n4640;
  assign n4642 = ~n4225 & n4270;
  assign n4643 = n4227 & ~n4642;
  assign n4644 = ~n4641 & ~n4643;
  assign n4645 = n4639 & n4644;
  assign n4646 = n4250 ^ n4176;
  assign n4647 = n4250 ^ n4175;
  assign n4648 = n4647 ^ n4175;
  assign n4649 = n4269 & ~n4284;
  assign n4650 = ~n4241 & n4649;
  assign n4651 = ~n4257 & n4650;
  assign n4652 = n4651 ^ n4175;
  assign n4653 = ~n4648 & n4652;
  assign n4654 = n4653 ^ n4175;
  assign n4655 = n4646 & n4654;
  assign n4656 = n4655 ^ n4176;
  assign n4657 = n4645 & ~n4656;
  assign n4658 = ~n4248 & n4657;
  assign n4659 = ~n4635 & n4658;
  assign n4660 = n4632 & n4659;
  assign n4661 = n4660 ^ n1505;
  assign n4662 = n4661 ^ x252;
  assign n4663 = n3725 & n3734;
  assign n4664 = n3717 & ~n4354;
  assign n4665 = ~n4663 & ~n4664;
  assign n4666 = ~n3712 & n3715;
  assign n4667 = n3734 & ~n4355;
  assign n4668 = ~n4666 & ~n4667;
  assign n4669 = n3711 & n3753;
  assign n4670 = n3720 & ~n3746;
  assign n4671 = ~n4669 & ~n4670;
  assign n4672 = ~n3740 & ~n3770;
  assign n4673 = ~n3725 & n4672;
  assign n4674 = ~n3750 & n4673;
  assign n4675 = n3717 & ~n4674;
  assign n4676 = ~n3727 & ~n3759;
  assign n4677 = ~n3769 & n4676;
  assign n4678 = n3713 & ~n4677;
  assign n4679 = ~n3738 & n3761;
  assign n4680 = n4672 & n4679;
  assign n4681 = n3722 & ~n4680;
  assign n4682 = ~n4678 & ~n4681;
  assign n4683 = ~n4675 & n4682;
  assign n4684 = n4671 & n4683;
  assign n4685 = n4668 & n4684;
  assign n4686 = n3743 & n4685;
  assign n4687 = n4665 & n4686;
  assign n4688 = ~n4351 & n4687;
  assign n4689 = ~n3716 & n4688;
  assign n4690 = n4343 & n4689;
  assign n4691 = n4690 ^ n1553;
  assign n4692 = n4691 ^ x253;
  assign n4693 = n4662 & ~n4692;
  assign n4694 = n4627 & n4693;
  assign n4695 = ~n4588 & ~n4626;
  assign n4696 = ~n4662 & ~n4692;
  assign n4697 = n4695 & n4696;
  assign n4698 = ~n4694 & ~n4697;
  assign n4699 = n4564 & ~n4698;
  assign n4700 = n4522 & ~n4563;
  assign n4701 = ~n4588 & n4626;
  assign n4702 = n4693 & n4701;
  assign n4703 = n4700 & n4702;
  assign n4704 = ~n4522 & n4563;
  assign n4705 = ~n4662 & n4692;
  assign n4706 = n4627 & n4705;
  assign n4707 = n4662 & n4692;
  assign n4708 = n4627 & n4707;
  assign n4709 = ~n4706 & ~n4708;
  assign n4710 = n4704 & ~n4709;
  assign n4711 = ~n4703 & ~n4710;
  assign n4712 = n4588 & n4626;
  assign n4713 = n4707 & n4712;
  assign n4714 = n4705 & n4712;
  assign n4715 = n4701 & n4707;
  assign n4716 = ~n4714 & ~n4715;
  assign n4717 = ~n4713 & n4716;
  assign n4718 = n4700 & ~n4717;
  assign n4719 = n4627 & n4696;
  assign n4720 = n4693 & n4695;
  assign n4721 = ~n4719 & ~n4720;
  assign n4722 = n4704 & ~n4721;
  assign n4723 = ~n4718 & ~n4722;
  assign n4724 = n4695 & n4707;
  assign n4725 = ~n4719 & ~n4724;
  assign n4726 = n4564 & ~n4725;
  assign n4727 = ~n4522 & ~n4563;
  assign n4728 = n4695 & n4705;
  assign n4729 = ~n4708 & n4725;
  assign n4730 = ~n4728 & n4729;
  assign n4731 = n4727 & ~n4730;
  assign n4732 = n4696 & n4701;
  assign n4733 = n4704 & n4732;
  assign n4734 = n4701 & n4705;
  assign n4735 = ~n4713 & ~n4734;
  assign n4736 = n4704 & ~n4735;
  assign n4737 = ~n4733 & ~n4736;
  assign n4738 = n4564 & n4702;
  assign n4739 = n4694 & n4700;
  assign n4740 = ~n4738 & ~n4739;
  assign n4741 = n4693 & n4712;
  assign n4742 = ~n4732 & ~n4741;
  assign n4743 = n4727 & ~n4742;
  assign n4744 = n4704 & n4741;
  assign n4745 = ~n4714 & n4735;
  assign n4746 = n4564 & ~n4745;
  assign n4747 = ~n4744 & ~n4746;
  assign n4748 = n4696 & n4712;
  assign n4749 = ~n4734 & ~n4748;
  assign n4750 = n4727 & ~n4749;
  assign n4751 = ~n4697 & ~n4706;
  assign n4752 = ~n4720 & n4751;
  assign n4753 = n4700 & ~n4752;
  assign n4754 = ~n4750 & ~n4753;
  assign n4755 = n4747 & n4754;
  assign n4756 = ~n4743 & n4755;
  assign n4757 = n4740 & n4756;
  assign n4758 = n4737 & n4757;
  assign n4759 = ~n4731 & n4758;
  assign n4760 = ~n4726 & n4759;
  assign n4761 = n4723 & n4760;
  assign n4762 = n4711 & n4761;
  assign n4763 = ~n4699 & n4762;
  assign n4764 = n4763 ^ n3267;
  assign n4765 = n4764 ^ x295;
  assign n4766 = n4171 ^ x237;
  assign n4767 = n4176 & n4265;
  assign n4768 = n4175 & n4284;
  assign n4769 = ~n4252 & ~n4264;
  assign n4770 = n4236 & ~n4769;
  assign n4771 = ~n4768 & ~n4770;
  assign n4772 = ~n4767 & n4771;
  assign n4773 = ~n4177 & n4238;
  assign n4774 = ~n4256 & ~n4773;
  assign n4775 = n4262 & ~n4267;
  assign n4776 = n4227 & ~n4775;
  assign n4777 = ~n4225 & ~n4268;
  assign n4778 = n4175 & ~n4777;
  assign n4779 = n4253 & n4633;
  assign n4780 = n4176 & ~n4779;
  assign n4781 = ~n4778 & ~n4780;
  assign n4782 = ~n4225 & ~n4232;
  assign n4783 = ~n4264 & n4782;
  assign n4784 = ~n4250 & n4783;
  assign n4785 = n4784 ^ n4174;
  assign n4786 = n4785 ^ n4784;
  assign n4787 = n4186 ^ n4178;
  assign n4788 = n4787 ^ n4223;
  assign n4789 = n4788 ^ n4178;
  assign n4790 = n4789 ^ n4184;
  assign n4791 = n4790 ^ n4223;
  assign n4792 = n4223 ^ n4184;
  assign n4793 = n4792 ^ n4184;
  assign n4794 = n4184 ^ n4178;
  assign n4795 = n4794 ^ n4184;
  assign n4796 = ~n4793 & n4795;
  assign n4797 = n4796 ^ n4184;
  assign n4798 = ~n4791 & ~n4797;
  assign n4799 = n4798 ^ n4788;
  assign n4800 = n4799 ^ n4784;
  assign n4801 = n4786 & n4800;
  assign n4802 = n4801 ^ n4784;
  assign n4803 = ~n4240 & ~n4802;
  assign n4804 = n4781 & ~n4803;
  assign n4805 = ~n4635 & n4804;
  assign n4806 = ~n4776 & n4805;
  assign n4807 = n4774 & n4806;
  assign n4808 = n4772 & n4807;
  assign n4809 = n4630 & n4808;
  assign n4810 = n4809 ^ n2044;
  assign n4811 = n4810 ^ x232;
  assign n4812 = ~n4766 & n4811;
  assign n4813 = n4433 ^ x236;
  assign n4814 = n3078 & n3116;
  assign n4815 = ~n3073 & ~n4814;
  assign n4816 = n2749 & n3130;
  assign n4817 = n3078 & ~n3107;
  assign n4818 = ~n4816 & ~n4817;
  assign n4819 = ~n3080 & n4543;
  assign n4820 = n3074 & ~n4819;
  assign n4821 = ~n3076 & ~n3115;
  assign n4822 = n3094 & ~n4821;
  assign n4823 = ~n3072 & ~n3123;
  assign n4824 = ~n3109 & n4823;
  assign n4825 = n3078 & ~n4824;
  assign n4826 = ~n3097 & n3107;
  assign n4827 = n2749 & ~n4826;
  assign n4828 = ~n4825 & ~n4827;
  assign n4829 = n3094 & n3101;
  assign n4830 = ~n3087 & n3118;
  assign n4831 = ~n3092 & n4830;
  assign n4832 = n3074 & ~n4831;
  assign n4833 = ~n4829 & ~n4832;
  assign n4834 = n4828 & n4833;
  assign n4835 = ~n3110 & n4834;
  assign n4836 = ~n3112 & n4835;
  assign n4837 = n4525 & n4836;
  assign n4838 = ~n4822 & n4837;
  assign n4839 = ~n4820 & n4838;
  assign n4840 = n4818 & n4839;
  assign n4841 = n4815 & n4840;
  assign n4842 = n4533 & n4841;
  assign n4843 = n3100 & n4842;
  assign n4844 = n4843 ^ n2773;
  assign n4845 = n4844 ^ x234;
  assign n4846 = n4813 & n4845;
  assign n4847 = ~n4589 & n4605;
  assign n4848 = ~n3863 & ~n3896;
  assign n4849 = n3788 & ~n4848;
  assign n4850 = ~n4847 & ~n4849;
  assign n4851 = n3880 & ~n3897;
  assign n4852 = n3788 & ~n4851;
  assign n4853 = n4602 & n4609;
  assign n4854 = n3860 & ~n4853;
  assign n4855 = ~n4852 & ~n4854;
  assign n4856 = ~n3890 & n4592;
  assign n4857 = ~n3887 & n4856;
  assign n4858 = n3895 & n4857;
  assign n4859 = n3874 & ~n4858;
  assign n4860 = ~n3867 & n4602;
  assign n4861 = ~n3872 & n4860;
  assign n4862 = ~n3882 & n4861;
  assign n4863 = n4605 & ~n4862;
  assign n4864 = ~n4859 & ~n4863;
  assign n4865 = n4855 & n4864;
  assign n4866 = n3877 & n4865;
  assign n4867 = n4850 & n4866;
  assign n4868 = ~n4621 & n4867;
  assign n4869 = ~n3859 & n4868;
  assign n4870 = ~n3855 & n4869;
  assign n4871 = n4870 ^ n2796;
  assign n4872 = n4871 ^ x235;
  assign n4873 = n3734 & n3750;
  assign n4874 = n3711 & n3732;
  assign n4875 = ~n4873 & ~n4874;
  assign n4876 = n3740 ^ n3713;
  assign n4877 = n3740 ^ n3712;
  assign n4878 = n4877 ^ n3712;
  assign n4879 = n3770 ^ n3712;
  assign n4880 = ~n4878 & n4879;
  assign n4881 = n4880 ^ n3712;
  assign n4882 = n4876 & ~n4881;
  assign n4883 = n4882 ^ n3713;
  assign n4884 = n4875 & ~n4883;
  assign n4885 = n3715 & n3717;
  assign n4886 = n3754 & ~n3769;
  assign n4887 = ~n3760 & n4886;
  assign n4888 = ~n3734 & n4887;
  assign n4889 = n3713 & ~n4886;
  assign n4890 = n4679 & ~n4889;
  assign n4891 = ~n3753 & n4890;
  assign n4892 = ~n4888 & ~n4891;
  assign n4893 = n4892 ^ n3712;
  assign n4894 = n4893 ^ n4892;
  assign n4895 = ~n3747 & n4365;
  assign n4896 = n4895 ^ n4892;
  assign n4897 = n4896 ^ n4892;
  assign n4898 = ~n4894 & ~n4897;
  assign n4899 = n4898 ^ n4892;
  assign n4900 = ~n3711 & n4899;
  assign n4901 = n4900 ^ n4892;
  assign n4902 = ~n4885 & ~n4901;
  assign n4903 = n4884 & n4902;
  assign n4904 = n4665 & n4903;
  assign n4905 = n4349 & n4904;
  assign n4906 = n3730 & n4905;
  assign n4907 = n4343 & n4906;
  assign n4908 = n4907 ^ n2008;
  assign n4909 = n4908 ^ x233;
  assign n4910 = ~n4872 & ~n4909;
  assign n4911 = n4846 & n4910;
  assign n4912 = ~n4813 & ~n4845;
  assign n4913 = n4910 & n4912;
  assign n4914 = ~n4911 & ~n4913;
  assign n4915 = n4812 & ~n4914;
  assign n4916 = n4811 ^ n4766;
  assign n4917 = n4813 & ~n4845;
  assign n4918 = n4910 & n4917;
  assign n4919 = n4918 ^ n4811;
  assign n4920 = n4919 ^ n4918;
  assign n4921 = n4872 & ~n4909;
  assign n4922 = n4846 & n4921;
  assign n4923 = n4912 & n4921;
  assign n4924 = ~n4922 & ~n4923;
  assign n4925 = n4924 ^ n4918;
  assign n4926 = n4920 & ~n4925;
  assign n4927 = n4926 ^ n4918;
  assign n4928 = ~n4916 & n4927;
  assign n4929 = ~n4915 & ~n4928;
  assign n4930 = n4812 & n4922;
  assign n4931 = n4766 & ~n4811;
  assign n4932 = n4872 & n4909;
  assign n4933 = ~n4813 & n4845;
  assign n4934 = n4932 & n4933;
  assign n4935 = ~n4872 & n4909;
  assign n4936 = n4846 & n4935;
  assign n4937 = n4912 & n4935;
  assign n4938 = n4917 & n4935;
  assign n4939 = ~n4937 & ~n4938;
  assign n4940 = ~n4936 & n4939;
  assign n4941 = ~n4934 & n4940;
  assign n4942 = n4931 & ~n4941;
  assign n4943 = ~n4930 & ~n4942;
  assign n4944 = ~n4766 & n4923;
  assign n4945 = ~n4766 & ~n4811;
  assign n4946 = n4917 & n4921;
  assign n4947 = ~n4937 & ~n4946;
  assign n4948 = n4945 & ~n4947;
  assign n4949 = ~n4944 & ~n4948;
  assign n4950 = n4766 & n4811;
  assign n4951 = n4910 & n4933;
  assign n4952 = ~n4918 & ~n4951;
  assign n4953 = n4950 & ~n4952;
  assign n4954 = n4938 & n4945;
  assign n4955 = n4921 & n4933;
  assign n4956 = n4931 & n4955;
  assign n4957 = n4933 & n4935;
  assign n4958 = n4945 & n4957;
  assign n4959 = ~n4956 & ~n4958;
  assign n4960 = n4846 & n4932;
  assign n4961 = ~n4936 & ~n4960;
  assign n4962 = n4945 & ~n4961;
  assign n4963 = n4912 & n4932;
  assign n4964 = ~n4936 & ~n4963;
  assign n4965 = n4917 & n4932;
  assign n4966 = ~n4934 & ~n4965;
  assign n4967 = n4964 & n4966;
  assign n4968 = n4950 & ~n4967;
  assign n4969 = ~n4962 & ~n4968;
  assign n4970 = ~n4922 & ~n4951;
  assign n4971 = ~n4946 & n4970;
  assign n4972 = n4931 & ~n4971;
  assign n4973 = ~n4938 & n4966;
  assign n4974 = ~n4963 & n4973;
  assign n4975 = n4812 & ~n4974;
  assign n4976 = ~n4972 & ~n4975;
  assign n4977 = n4969 & n4976;
  assign n4978 = n4959 & n4977;
  assign n4979 = ~n4954 & n4978;
  assign n4980 = ~n4953 & n4979;
  assign n4981 = n4949 & n4980;
  assign n4982 = n4943 & n4981;
  assign n4983 = n4929 & n4982;
  assign n4984 = n4983 ^ n3238;
  assign n4985 = n4984 ^ x293;
  assign n4986 = n4765 & n4985;
  assign n4987 = n3146 ^ x227;
  assign n4988 = n4117 & n4150;
  assign n4989 = ~n4114 & n4153;
  assign n4990 = ~n4988 & ~n4989;
  assign n4991 = n4053 & n4126;
  assign n4992 = ~n4108 & ~n4111;
  assign n4993 = n4117 & ~n4992;
  assign n4994 = ~n4991 & ~n4993;
  assign n4995 = n4119 & n4153;
  assign n4998 = n4076 ^ n4075;
  assign n4999 = n4998 ^ n4106;
  assign n4996 = n4076 & ~n4106;
  assign n4997 = n4078 & n4996;
  assign n5000 = n4999 ^ n4997;
  assign n5001 = n4121 & n5000;
  assign n5002 = n4114 & ~n4136;
  assign n5003 = ~n4119 & n5002;
  assign n5004 = n4053 & ~n5003;
  assign n5005 = ~n4145 & ~n4162;
  assign n5006 = ~n4144 & n5005;
  assign n5007 = ~n4126 & n5006;
  assign n5008 = n4153 & ~n5007;
  assign n5009 = ~n4137 & ~n4165;
  assign n5010 = ~n4144 & n5009;
  assign n5011 = ~n4130 & n5010;
  assign n5012 = n4117 & ~n5011;
  assign n5013 = ~n5008 & ~n5012;
  assign n5014 = ~n5004 & n5013;
  assign n5015 = ~n5001 & n5014;
  assign n5016 = ~n4995 & n5015;
  assign n5017 = n5006 ^ n4134;
  assign n5018 = n5017 ^ n4134;
  assign n5019 = n4134 ^ n4052;
  assign n5020 = n5019 ^ n4134;
  assign n5021 = ~n5018 & n5020;
  assign n5022 = n5021 ^ n4134;
  assign n5023 = n4124 & n5022;
  assign n5024 = n5023 ^ n4134;
  assign n5025 = n5016 & ~n5024;
  assign n5026 = n4994 & n5025;
  assign n5027 = n4990 & n5026;
  assign n5028 = n5027 ^ n2112;
  assign n5029 = n5028 ^ x229;
  assign n5030 = n4810 ^ x230;
  assign n5031 = ~n5029 & ~n5030;
  assign n5032 = n3372 ^ x226;
  assign n5033 = n4908 ^ x231;
  assign n5034 = n5032 & ~n5033;
  assign n5035 = n5031 & n5034;
  assign n5036 = ~n4987 & n5035;
  assign n5037 = ~n5032 & ~n5033;
  assign n5038 = n2595 & n2609;
  assign n5039 = ~n2633 & ~n5038;
  assign n5040 = ~n2598 & ~n2629;
  assign n5041 = n1689 & ~n5040;
  assign n5042 = ~n2601 & n2651;
  assign n5043 = n2609 & ~n5042;
  assign n5044 = ~n2645 & ~n4003;
  assign n5045 = ~n2617 & ~n2643;
  assign n5046 = n2327 & ~n5045;
  assign n5047 = n2630 & n4013;
  assign n5048 = n2609 & ~n5047;
  assign n5049 = ~n5046 & ~n5048;
  assign n5050 = ~n5044 & n5049;
  assign n5051 = n1689 & ~n4018;
  assign n5052 = n2603 & n2651;
  assign n5053 = ~n2636 & n5052;
  assign n5054 = n2625 & ~n5053;
  assign n5055 = ~n5051 & ~n5054;
  assign n5056 = n5050 & n5055;
  assign n5057 = ~n5043 & n5056;
  assign n5058 = ~n5041 & n5057;
  assign n5059 = n4012 ^ n2327;
  assign n5060 = n4012 ^ n1689;
  assign n5061 = n5060 ^ n1689;
  assign n5062 = ~n2627 & n4023;
  assign n5063 = n5062 ^ n1689;
  assign n5064 = ~n5061 & n5063;
  assign n5065 = n5064 ^ n1689;
  assign n5066 = n5059 & n5065;
  assign n5067 = n5066 ^ n2327;
  assign n5068 = n5058 & ~n5067;
  assign n5069 = n5039 & n5068;
  assign n5070 = n5069 ^ n2076;
  assign n5071 = n5070 ^ x228;
  assign n5072 = ~n5029 & n5030;
  assign n5073 = n4987 & n5072;
  assign n5074 = n5071 & n5073;
  assign n5075 = n5029 & ~n5030;
  assign n5076 = ~n4987 & ~n5071;
  assign n5077 = n5075 & n5076;
  assign n5078 = n4987 & n5075;
  assign n5079 = ~n5071 & n5078;
  assign n5080 = ~n5077 & ~n5079;
  assign n5081 = ~n5074 & n5080;
  assign n5082 = n5037 & ~n5081;
  assign n5083 = ~n5036 & ~n5082;
  assign n5084 = ~n5032 & n5033;
  assign n5085 = n5071 ^ n4987;
  assign n5086 = n5085 ^ n5029;
  assign n5087 = n5086 ^ n4987;
  assign n5088 = n5030 ^ n4987;
  assign n5089 = n5088 ^ n5030;
  assign n5090 = n5030 ^ n5029;
  assign n5091 = n5090 ^ n5030;
  assign n5092 = n5089 & ~n5091;
  assign n5093 = n5092 ^ n5030;
  assign n5094 = n5087 & n5093;
  assign n5095 = n5094 ^ n5085;
  assign n5096 = n5084 & ~n5095;
  assign n5097 = ~n4987 & n5071;
  assign n5098 = ~n5075 & n5097;
  assign n5099 = n4987 & ~n5090;
  assign n5100 = ~n5071 & n5099;
  assign n5101 = n4987 & n5071;
  assign n5102 = ~n5076 & ~n5101;
  assign n5103 = n5075 & ~n5102;
  assign n5104 = ~n5100 & ~n5103;
  assign n5105 = ~n5098 & n5104;
  assign n5106 = n5034 & ~n5105;
  assign n5107 = ~n5096 & ~n5106;
  assign n5108 = n5033 ^ n5032;
  assign n5109 = ~n5076 & ~n5090;
  assign n5110 = n5072 & n5076;
  assign n5111 = n5075 & n5097;
  assign n5112 = ~n5110 & ~n5111;
  assign n5113 = ~n5109 & n5112;
  assign n5114 = n5113 ^ n5033;
  assign n5115 = n5114 ^ n5113;
  assign n5116 = n5031 & n5101;
  assign n5117 = n5029 & n5030;
  assign n5118 = n5071 & n5117;
  assign n5119 = n5112 & ~n5118;
  assign n5120 = ~n5116 & n5119;
  assign n5121 = n5120 ^ n5113;
  assign n5122 = ~n5115 & n5121;
  assign n5123 = n5122 ^ n5113;
  assign n5124 = ~n5108 & ~n5123;
  assign n5125 = n5107 & ~n5124;
  assign n5126 = n5083 & n5125;
  assign n5127 = n5126 ^ n3272;
  assign n5128 = n5127 ^ x294;
  assign n5129 = n3784 ^ x219;
  assign n5130 = n4605 & ~n4857;
  assign n5131 = n3788 & ~n4607;
  assign n5132 = ~n5130 & ~n5131;
  assign n5133 = ~n3786 & n3854;
  assign n5134 = ~n3878 & ~n3884;
  assign n5135 = ~n5133 & ~n5134;
  assign n5136 = ~n3887 & n3898;
  assign n5137 = n3874 & ~n5136;
  assign n5138 = ~n3858 & n4861;
  assign n5139 = n3860 & ~n5138;
  assign n5140 = ~n5137 & ~n5139;
  assign n5141 = n5135 & n5140;
  assign n5142 = n5132 & n5141;
  assign n5143 = n4850 & n5142;
  assign n5144 = n4591 & n5143;
  assign n5145 = ~n3859 & n5144;
  assign n5146 = n5145 ^ n1716;
  assign n5147 = n5146 ^ x214;
  assign n5148 = ~n5129 & n5147;
  assign n5149 = ~n4119 & ~n4162;
  assign n5150 = n4117 & ~n5149;
  assign n5151 = ~n4134 & ~n4146;
  assign n5152 = ~n4136 & n5151;
  assign n5153 = n5009 & n5152;
  assign n5154 = ~n4150 & n5153;
  assign n5155 = n4121 & ~n5154;
  assign n5156 = ~n5150 & ~n5155;
  assign n5157 = n4129 & n4153;
  assign n5158 = ~n4108 & ~n4136;
  assign n5159 = ~n4137 & n5158;
  assign n5160 = ~n4124 & ~n5159;
  assign n5161 = ~n4129 & ~n4165;
  assign n5162 = n4148 & n5161;
  assign n5163 = n4053 & ~n5162;
  assign n5164 = ~n5160 & ~n5163;
  assign n5165 = ~n5157 & n5164;
  assign n5166 = n5156 & n5165;
  assign n5167 = n4133 & n5166;
  assign n5168 = n4990 & n5167;
  assign n5169 = ~n4116 & n5168;
  assign n5170 = ~n4169 & n5169;
  assign n5171 = n5170 ^ n1850;
  assign n5172 = n5171 ^ x215;
  assign n5173 = n4176 & n4267;
  assign n5174 = n4175 & n4260;
  assign n5175 = ~n5173 & ~n5174;
  assign n5176 = n4177 & n4250;
  assign n5177 = ~n4244 & ~n4259;
  assign n5178 = n4236 & ~n5177;
  assign n5179 = ~n5176 & ~n5178;
  assign n5180 = n5175 & n5179;
  assign n5181 = n4233 & ~n4257;
  assign n5182 = ~n4177 & ~n5181;
  assign n5183 = n4227 & ~n4651;
  assign n5184 = ~n5182 & ~n5183;
  assign n5185 = n5180 & n5184;
  assign n5186 = n4772 & n5185;
  assign n5187 = n4235 & n5186;
  assign n5188 = n4249 & n5187;
  assign n5189 = n4632 & n5188;
  assign n5190 = n5189 ^ n1765;
  assign n5191 = n5190 ^ x216;
  assign n5192 = ~n5172 & ~n5191;
  assign n5193 = n2668 ^ x218;
  assign n5194 = n3337 & n3338;
  assign n5195 = ~n3332 & ~n3339;
  assign n5196 = ~n3325 & n5195;
  assign n5197 = n3322 & ~n5196;
  assign n5198 = ~n5194 & ~n5197;
  assign n5199 = n3313 & ~n3344;
  assign n5200 = ~n3307 & ~n3316;
  assign n5201 = n3213 & ~n5200;
  assign n5202 = ~n3321 & ~n4312;
  assign n5203 = n3214 & ~n5202;
  assign n5204 = n4313 ^ n3322;
  assign n5205 = n5204 ^ n4313;
  assign n5206 = ~n3340 & ~n4565;
  assign n5207 = n5206 ^ n5195;
  assign n5208 = n5195 ^ n3214;
  assign n5209 = n5208 ^ n3214;
  assign n5210 = n4324 ^ n3214;
  assign n5211 = n5209 & ~n5210;
  assign n5212 = n5211 ^ n3214;
  assign n5213 = n5207 & n5212;
  assign n5214 = n5213 ^ n5206;
  assign n5215 = ~n3355 & n5214;
  assign n5216 = n5215 ^ n4313;
  assign n5217 = ~n5205 & n5216;
  assign n5218 = n5217 ^ n4313;
  assign n5219 = ~n5203 & n5218;
  assign n5220 = n3330 & n5219;
  assign n5221 = ~n5201 & n5220;
  assign n5222 = ~n5199 & n5221;
  assign n5223 = n5198 & n5222;
  assign n5224 = ~n4584 & n5223;
  assign n5225 = ~n4326 & n5224;
  assign n5226 = ~n3323 & n5225;
  assign n5227 = n5226 ^ n1893;
  assign n5228 = n5227 ^ x217;
  assign n5229 = ~n5193 & ~n5228;
  assign n5230 = n5192 & n5229;
  assign n5231 = n5148 & n5230;
  assign n5232 = n5129 & n5147;
  assign n5233 = n5193 & n5228;
  assign n5234 = n5192 & n5233;
  assign n5235 = n5232 & n5234;
  assign n5236 = ~n5172 & n5191;
  assign n5237 = n5233 & n5236;
  assign n5238 = n5148 & n5237;
  assign n5239 = ~n5235 & ~n5238;
  assign n5240 = ~n5129 & ~n5147;
  assign n5241 = ~n5193 & n5228;
  assign n5242 = n5236 & n5241;
  assign n5243 = n5193 & ~n5228;
  assign n5244 = n5192 & n5243;
  assign n5245 = ~n5242 & ~n5244;
  assign n5246 = n5240 & ~n5245;
  assign n5247 = n5172 & n5191;
  assign n5248 = n5241 & n5247;
  assign n5249 = n5243 & n5247;
  assign n5250 = ~n5248 & ~n5249;
  assign n5251 = n5148 & ~n5250;
  assign n5252 = ~n5246 & ~n5251;
  assign n5253 = n5239 & n5252;
  assign n5254 = ~n5231 & n5253;
  assign n5255 = n5129 & ~n5147;
  assign n5256 = n5230 & n5255;
  assign n5257 = n5229 & n5247;
  assign n5258 = n5232 & n5257;
  assign n5259 = n5236 & n5243;
  assign n5260 = n5255 & n5259;
  assign n5261 = ~n5258 & ~n5260;
  assign n5262 = ~n5256 & n5261;
  assign n5263 = n5229 & n5236;
  assign n5264 = n5148 & n5263;
  assign n5265 = ~n5148 & ~n5255;
  assign n5266 = n5192 & n5241;
  assign n5267 = n5265 & n5266;
  assign n5268 = n5232 & n5244;
  assign n5269 = ~n5267 & ~n5268;
  assign n5270 = ~n5264 & n5269;
  assign n5271 = n5228 ^ n5193;
  assign n5272 = n5228 ^ n5191;
  assign n5273 = n5272 ^ n5191;
  assign n5274 = n5191 ^ n5172;
  assign n5275 = n5274 ^ n5191;
  assign n5276 = ~n5273 & n5275;
  assign n5277 = n5276 ^ n5191;
  assign n5278 = ~n5271 & n5277;
  assign n5279 = n5232 & n5278;
  assign n5280 = n5172 & ~n5191;
  assign n5281 = n5243 & n5280;
  assign n5282 = ~n5234 & ~n5257;
  assign n5283 = ~n5281 & n5282;
  assign n5284 = n5148 & ~n5283;
  assign n5285 = n5229 & n5280;
  assign n5286 = n5233 & n5247;
  assign n5287 = n5241 & n5280;
  assign n5288 = ~n5286 & ~n5287;
  assign n5289 = ~n5249 & n5288;
  assign n5290 = ~n5259 & n5289;
  assign n5291 = ~n5285 & n5290;
  assign n5292 = n5240 & ~n5291;
  assign n5293 = n5233 & n5280;
  assign n5294 = ~n5248 & ~n5281;
  assign n5295 = ~n5293 & n5294;
  assign n5296 = ~n5287 & n5295;
  assign n5297 = ~n5249 & n5296;
  assign n5298 = ~n5242 & n5297;
  assign n5299 = n5255 & ~n5298;
  assign n5300 = ~n5292 & ~n5299;
  assign n5301 = ~n5284 & n5300;
  assign n5302 = ~n5279 & n5301;
  assign n5303 = n5270 & n5302;
  assign n5304 = n5262 & n5303;
  assign n5305 = n5254 & n5304;
  assign n5306 = n5305 ^ n3304;
  assign n5307 = n5306 ^ x296;
  assign n5308 = n5128 & ~n5307;
  assign n5309 = n4986 & n5308;
  assign n5310 = n5128 & n5307;
  assign n5311 = ~n4765 & n4985;
  assign n5312 = n5310 & n5311;
  assign n5313 = ~n5309 & ~n5312;
  assign n5314 = n4503 & ~n5313;
  assign n5315 = ~n3999 & n4502;
  assign n5316 = n5308 & n5311;
  assign n5317 = ~n5128 & n5307;
  assign n5318 = n5311 & n5317;
  assign n5319 = ~n5316 & ~n5318;
  assign n5320 = n5315 & ~n5319;
  assign n5321 = ~n5314 & ~n5320;
  assign n5322 = n4765 & ~n4985;
  assign n5323 = n5308 & n5322;
  assign n5324 = n5315 & n5323;
  assign n5325 = ~n4765 & ~n4985;
  assign n5326 = n5308 & n5325;
  assign n5327 = n4503 & n5326;
  assign n5328 = ~n5324 & ~n5327;
  assign n5329 = n5317 & n5325;
  assign n5330 = n4503 & n5329;
  assign n5331 = ~n3999 & ~n4502;
  assign n5332 = ~n5312 & ~n5323;
  assign n5333 = n5331 & ~n5332;
  assign n5334 = ~n5128 & ~n5307;
  assign n5335 = n4986 & n5334;
  assign n5336 = n5317 & n5322;
  assign n5337 = ~n5335 & ~n5336;
  assign n5338 = ~n5323 & n5337;
  assign n5339 = n4503 & ~n5338;
  assign n5340 = ~n5333 & ~n5339;
  assign n5341 = n3999 & ~n4502;
  assign n5342 = n5310 & n5322;
  assign n5343 = ~n5318 & ~n5335;
  assign n5344 = ~n5342 & n5343;
  assign n5345 = ~n5326 & ~n5329;
  assign n5346 = ~n5336 & n5345;
  assign n5347 = n5344 & n5346;
  assign n5348 = n5332 & n5347;
  assign n5349 = n5341 & n5348;
  assign n5350 = ~n5309 & ~n5342;
  assign n5351 = n5315 & ~n5350;
  assign n5352 = n5310 & n5325;
  assign n5353 = n5322 & n5334;
  assign n5354 = ~n5352 & ~n5353;
  assign n5355 = ~n5329 & n5354;
  assign n5356 = ~n3999 & ~n5355;
  assign n5357 = ~n5351 & ~n5356;
  assign n5358 = ~n5349 & n5357;
  assign n5359 = n5340 & n5358;
  assign n5360 = n5311 & n5334;
  assign n5361 = n5360 ^ n5331;
  assign n5362 = n5331 ^ n4503;
  assign n5363 = n5362 ^ n4503;
  assign n5364 = n4986 & n5310;
  assign n5365 = ~n5335 & ~n5364;
  assign n5366 = n5365 ^ n4503;
  assign n5367 = n5363 & n5366;
  assign n5368 = n5367 ^ n4503;
  assign n5369 = n5361 & ~n5368;
  assign n5370 = n5369 ^ n5360;
  assign n5371 = n5359 & ~n5370;
  assign n5372 = ~n5330 & n5371;
  assign n5373 = n5328 & n5372;
  assign n5374 = n5321 & n5373;
  assign n5375 = n5374 ^ n3372;
  assign n5376 = n5375 ^ x322;
  assign n5377 = n4700 & ~n4735;
  assign n5378 = ~n4721 & n4727;
  assign n5379 = ~n5377 & ~n5378;
  assign n5380 = n4704 & n4728;
  assign n5381 = n4564 & ~n4716;
  assign n5382 = ~n5380 & ~n5381;
  assign n5383 = ~n4694 & ~n4724;
  assign n5384 = ~n4708 & n5383;
  assign n5385 = n4700 & ~n5384;
  assign n5386 = ~n4709 & n4727;
  assign n5387 = n4727 & ~n4735;
  assign n5388 = n4563 ^ n4522;
  assign n5389 = ~n4702 & ~n4741;
  assign n5390 = ~n5388 & ~n5389;
  assign n5391 = ~n5387 & ~n5390;
  assign n5392 = ~n4697 & ~n4748;
  assign n5393 = n4700 & ~n5392;
  assign n5394 = n4721 & n4751;
  assign n5395 = n4564 & ~n5394;
  assign n5396 = ~n4715 & n5392;
  assign n5397 = ~n4741 & n5396;
  assign n5398 = n4704 & ~n5397;
  assign n5399 = ~n5395 & ~n5398;
  assign n5400 = ~n5393 & n5399;
  assign n5401 = n5391 & n5400;
  assign n5402 = ~n5386 & n5401;
  assign n5403 = ~n5385 & n5402;
  assign n5404 = ~n4733 & n5403;
  assign n5405 = n4711 & n5404;
  assign n5406 = n5382 & n5405;
  assign n5407 = n5379 & n5406;
  assign n5408 = n5407 ^ n2914;
  assign n5409 = n5408 ^ x261;
  assign n5410 = n4131 & n5152;
  assign n5411 = n4153 & ~n5410;
  assign n5412 = ~n4117 & ~n4145;
  assign n5413 = ~n5006 & ~n5412;
  assign n5414 = ~n4124 & n5413;
  assign n5415 = ~n5411 & ~n5414;
  assign n5416 = n4141 & ~n4162;
  assign n5417 = n4121 & ~n5416;
  assign n5418 = n4113 & ~n4124;
  assign n5419 = n4992 & n5010;
  assign n5420 = ~n4150 & n5419;
  assign n5421 = ~n4119 & n5420;
  assign n5422 = n4053 & ~n5421;
  assign n5423 = ~n5418 & ~n5422;
  assign n5424 = ~n5417 & n5423;
  assign n5425 = n5415 & n5424;
  assign n5426 = n4994 & n5425;
  assign n5427 = n4123 & n5426;
  assign n5428 = ~n4169 & n5427;
  assign n5429 = n5428 ^ n2965;
  assign n5430 = n5429 ^ x247;
  assign n5431 = n4049 ^ x245;
  assign n5432 = ~n5430 & ~n5431;
  assign n5433 = n3530 & n4426;
  assign n5434 = n3534 & ~n5433;
  assign n5435 = n3514 & n4422;
  assign n5436 = n3549 & ~n5435;
  assign n5437 = ~n5434 & ~n5436;
  assign n5438 = n3508 & n4399;
  assign n5439 = n3414 & ~n4423;
  assign n5440 = ~n5438 & ~n5439;
  assign n5441 = n5437 & n5440;
  assign n5442 = ~n4518 & n5441;
  assign n5443 = n5442 ^ n2924;
  assign n5444 = n5443 ^ x246;
  assign n5445 = n4562 ^ x248;
  assign n5446 = ~n5444 & n5445;
  assign n5447 = n5432 & n5446;
  assign n5448 = n5430 & ~n5431;
  assign n5449 = n5444 & ~n5445;
  assign n5450 = n5448 & n5449;
  assign n5451 = ~n5447 & ~n5450;
  assign n5452 = n4625 ^ x249;
  assign n5453 = n4305 ^ x244;
  assign n5454 = n5452 & ~n5453;
  assign n5455 = ~n5451 & n5454;
  assign n5456 = ~n5430 & n5431;
  assign n5457 = n5444 & n5445;
  assign n5458 = n5456 & n5457;
  assign n5459 = n5430 & n5431;
  assign n5460 = n5449 & n5459;
  assign n5461 = ~n5458 & ~n5460;
  assign n5462 = n5461 ^ n5453;
  assign n5463 = n5462 ^ n5461;
  assign n5464 = n5446 & n5456;
  assign n5465 = n5449 & n5456;
  assign n5466 = ~n5464 & ~n5465;
  assign n5467 = n5466 ^ n5461;
  assign n5468 = ~n5463 & n5467;
  assign n5469 = n5468 ^ n5461;
  assign n5470 = n5452 & ~n5469;
  assign n5471 = ~n5455 & ~n5470;
  assign n5472 = n5446 & n5448;
  assign n5473 = n5454 & n5472;
  assign n5474 = ~n5452 & n5453;
  assign n5475 = n5445 ^ n5444;
  assign n5476 = n5432 & ~n5475;
  assign n5477 = n5451 & ~n5458;
  assign n5478 = n5459 & ~n5475;
  assign n5479 = n5477 & ~n5478;
  assign n5480 = ~n5476 & n5479;
  assign n5481 = ~n5465 & n5480;
  assign n5482 = n5474 & ~n5481;
  assign n5483 = ~n5473 & ~n5482;
  assign n5484 = ~n5452 & ~n5453;
  assign n5485 = n5448 & n5457;
  assign n5486 = ~n5444 & ~n5445;
  assign n5487 = n5459 & n5486;
  assign n5488 = n5432 & n5475;
  assign n5489 = ~n5472 & ~n5488;
  assign n5490 = ~n5450 & n5489;
  assign n5491 = ~n5487 & n5490;
  assign n5492 = ~n5458 & n5491;
  assign n5493 = ~n5464 & n5492;
  assign n5494 = ~n5485 & n5493;
  assign n5495 = n5484 & n5494;
  assign n5496 = n5452 & n5453;
  assign n5497 = ~n5476 & ~n5485;
  assign n5498 = n5496 & ~n5497;
  assign n5499 = n5432 & n5449;
  assign n5500 = ~n5454 & ~n5487;
  assign n5501 = n5478 & ~n5500;
  assign n5502 = ~n5499 & ~n5501;
  assign n5503 = ~n5464 & n5502;
  assign n5504 = n5452 & ~n5503;
  assign n5505 = ~n5498 & ~n5504;
  assign n5506 = ~n5495 & n5505;
  assign n5507 = n5483 & n5506;
  assign n5508 = n5471 & n5507;
  assign n5509 = n5508 ^ n3710;
  assign n5510 = n5509 ^ x256;
  assign n5511 = n5409 & n5510;
  assign n5512 = n4931 & ~n4964;
  assign n5513 = ~n4911 & ~n4946;
  assign n5514 = n4812 & ~n5513;
  assign n5515 = ~n5512 & ~n5514;
  assign n5516 = n4812 & n4923;
  assign n5517 = ~n4946 & ~n4951;
  assign n5518 = ~n4916 & ~n5517;
  assign n5519 = ~n4911 & ~n4922;
  assign n5520 = ~n4918 & n5519;
  assign n5521 = n4931 & ~n5520;
  assign n5522 = ~n4960 & ~n4963;
  assign n5523 = ~n4965 & n5522;
  assign n5524 = n4945 & ~n5523;
  assign n5525 = ~n5521 & ~n5524;
  assign n5526 = n4940 & ~n4965;
  assign n5527 = n4812 & ~n5526;
  assign n5529 = ~n4913 & ~n4922;
  assign n5528 = ~n4960 & n4973;
  assign n5530 = n5529 ^ n5528;
  assign n5531 = n5529 ^ n4950;
  assign n5532 = n5529 & n5531;
  assign n5533 = n5532 ^ n5529;
  assign n5534 = n5530 & n5533;
  assign n5535 = n5534 ^ n5532;
  assign n5536 = n5535 ^ n5529;
  assign n5537 = n5536 ^ n4950;
  assign n5538 = ~n5527 & n5537;
  assign n5539 = n5538 ^ n5527;
  assign n5540 = n5525 & ~n5539;
  assign n5541 = n4959 & n5540;
  assign n5542 = ~n5518 & n5541;
  assign n5543 = ~n5516 & n5542;
  assign n5544 = ~n4937 & ~n4957;
  assign n5545 = n5544 ^ n4955;
  assign n5546 = n5545 ^ n4955;
  assign n5547 = n4955 ^ n4811;
  assign n5548 = n5547 ^ n4955;
  assign n5549 = ~n5546 & ~n5548;
  assign n5550 = n5549 ^ n4955;
  assign n5551 = n4766 & n5550;
  assign n5552 = n5551 ^ n4955;
  assign n5553 = n5543 & ~n5552;
  assign n5554 = n5515 & n5553;
  assign n5555 = ~n4954 & n5554;
  assign n5556 = n5555 ^ n3606;
  assign n5557 = n5556 ^ x259;
  assign n5558 = n4448 & n4474;
  assign n5559 = n4393 & n4443;
  assign n5560 = ~n5558 & ~n5559;
  assign n5561 = ~n4393 & ~n4475;
  assign n5562 = n4435 & ~n5561;
  assign n5563 = ~n4437 & ~n4446;
  assign n5564 = n4443 & ~n5563;
  assign n5565 = ~n5562 & ~n5564;
  assign n5566 = n4443 & n4465;
  assign n5567 = n4435 & n4437;
  assign n5568 = ~n5566 & ~n5567;
  assign n5569 = ~n4050 & n4468;
  assign n5570 = n4461 & ~n4476;
  assign n5571 = n4444 & ~n5570;
  assign n5572 = ~n5569 & ~n5571;
  assign n5573 = ~n4454 & ~n4468;
  assign n5574 = ~n4446 & n5573;
  assign n5575 = n4448 & ~n5574;
  assign n5576 = n4392 & n4453;
  assign n5577 = ~n4474 & ~n5576;
  assign n5578 = n4470 & n5577;
  assign n5579 = n4464 & ~n5578;
  assign n5580 = ~n4443 & n4484;
  assign n5581 = n4483 & ~n5576;
  assign n5582 = ~n4435 & n5581;
  assign n5583 = ~n5580 & ~n5582;
  assign n5584 = ~n4486 & ~n5583;
  assign n5585 = ~n4444 & ~n5584;
  assign n5586 = ~n5579 & ~n5585;
  assign n5587 = ~n5575 & n5586;
  assign n5588 = n5572 & n5587;
  assign n5589 = n5568 & n5588;
  assign n5590 = n5565 & n5589;
  assign n5591 = n5560 & n5590;
  assign n5592 = n5591 ^ n2747;
  assign n5593 = n5592 ^ x260;
  assign n5594 = ~n5557 & n5593;
  assign n5595 = n5071 & n5078;
  assign n5596 = ~n5071 & n5073;
  assign n5597 = ~n5098 & ~n5596;
  assign n5598 = n5037 & ~n5597;
  assign n5599 = ~n5595 & ~n5598;
  assign n5600 = n5031 & n5097;
  assign n5601 = ~n5074 & ~n5600;
  assign n5602 = ~n5100 & n5601;
  assign n5603 = n5112 & n5602;
  assign n5604 = ~n5078 & n5603;
  assign n5605 = n5084 & ~n5604;
  assign n5606 = n5599 & ~n5605;
  assign n5607 = ~n5071 & n5117;
  assign n5608 = n5030 & ~n5102;
  assign n5609 = ~n5607 & ~n5608;
  assign n5610 = n5034 & ~n5609;
  assign n5611 = n5032 & n5033;
  assign n5612 = ~n4987 & n5117;
  assign n5613 = n5071 & ~n5090;
  assign n5614 = ~n5103 & ~n5613;
  assign n5615 = ~n5612 & n5614;
  assign n5616 = ~n5596 & n5615;
  assign n5617 = n5611 & ~n5616;
  assign n5618 = ~n5610 & ~n5617;
  assign n5619 = n5606 & n5618;
  assign n5620 = n5083 & n5619;
  assign n5621 = n5620 ^ n3673;
  assign n5622 = n5621 ^ x257;
  assign n5623 = n5232 & n5242;
  assign n5624 = n5148 & n5259;
  assign n5625 = ~n5623 & ~n5624;
  assign n5626 = n5237 & n5240;
  assign n5627 = n5255 & n5281;
  assign n5628 = ~n5626 & ~n5627;
  assign n5629 = n5625 & n5628;
  assign n5630 = n5230 & n5232;
  assign n5631 = n5255 & ~n5289;
  assign n5632 = ~n5630 & ~n5631;
  assign n5633 = ~n5266 & ~n5285;
  assign n5634 = n5240 & ~n5633;
  assign n5648 = n5286 ^ n5250;
  assign n5649 = n5250 ^ n5232;
  assign n5650 = n5649 ^ n5232;
  assign n5651 = ~n5240 & ~n5249;
  assign n5652 = n5651 ^ n5232;
  assign n5653 = ~n5650 & n5652;
  assign n5654 = n5653 ^ n5232;
  assign n5655 = ~n5648 & ~n5654;
  assign n5656 = n5655 ^ n5286;
  assign n5657 = ~n5293 & ~n5656;
  assign n5658 = ~n5257 & n5657;
  assign n5637 = ~n5281 & ~n5287;
  assign n5638 = ~n5257 & n5637;
  assign n5635 = ~n5242 & n5633;
  assign n5636 = ~n5244 & n5635;
  assign n5639 = n5638 ^ n5636;
  assign n5640 = ~n5255 & ~n5285;
  assign n5641 = n5640 ^ n5636;
  assign n5642 = n5641 ^ n5640;
  assign n5643 = n5640 ^ n5148;
  assign n5644 = n5642 & n5643;
  assign n5645 = n5644 ^ n5640;
  assign n5646 = n5639 & ~n5645;
  assign n5647 = n5646 ^ n5638;
  assign n5659 = n5658 ^ n5647;
  assign n5660 = n5265 & n5659;
  assign n5661 = n5660 ^ n5647;
  assign n5662 = ~n5634 & n5661;
  assign n5663 = n5244 ^ n5242;
  assign n5664 = n5663 ^ n5242;
  assign n5665 = n5255 ^ n5242;
  assign n5666 = n5665 ^ n5242;
  assign n5667 = n5664 & ~n5666;
  assign n5668 = n5667 ^ n5242;
  assign n5669 = ~n5148 & n5668;
  assign n5670 = n5669 ^ n5242;
  assign n5671 = n5662 & ~n5670;
  assign n5672 = n5632 & n5671;
  assign n5673 = n5239 & n5672;
  assign n5674 = ~n5231 & n5673;
  assign n5675 = n5629 & n5674;
  assign n5676 = n5675 ^ n3638;
  assign n5677 = n5676 ^ x258;
  assign n5678 = n5622 & n5677;
  assign n5679 = n5594 & n5678;
  assign n5680 = n5511 & n5679;
  assign n5681 = ~n5409 & n5510;
  assign n5682 = n5557 & n5593;
  assign n5683 = n5678 & n5682;
  assign n5684 = n5681 & n5683;
  assign n5685 = ~n5680 & ~n5684;
  assign n5686 = n5409 & ~n5510;
  assign n5687 = ~n5557 & ~n5593;
  assign n5688 = n5678 & n5687;
  assign n5689 = n5557 & ~n5593;
  assign n5690 = n5678 & n5689;
  assign n5691 = n5622 & ~n5677;
  assign n5692 = n5682 & n5691;
  assign n5693 = ~n5690 & ~n5692;
  assign n5694 = ~n5688 & n5693;
  assign n5695 = n5686 & ~n5694;
  assign n5696 = n5689 & n5691;
  assign n5697 = n5511 & n5696;
  assign n5698 = ~n5622 & ~n5677;
  assign n5699 = n5594 & n5698;
  assign n5700 = ~n5688 & ~n5699;
  assign n5701 = n5681 & ~n5700;
  assign n5702 = ~n5697 & ~n5701;
  assign n5703 = ~n5695 & n5702;
  assign n5704 = ~n5409 & ~n5510;
  assign n5705 = n5687 & n5691;
  assign n5706 = n5704 & n5705;
  assign n5707 = ~n5622 & n5677;
  assign n5708 = n5682 & n5707;
  assign n5709 = n5686 & n5708;
  assign n5710 = n5689 & n5707;
  assign n5711 = n5511 & n5710;
  assign n5712 = ~n5709 & ~n5711;
  assign n5713 = ~n5706 & n5712;
  assign n5714 = n5679 & n5704;
  assign n5715 = n5681 & n5696;
  assign n5716 = ~n5714 & ~n5715;
  assign n5717 = n5682 & n5698;
  assign n5718 = ~n5708 & ~n5710;
  assign n5719 = ~n5717 & n5718;
  assign n5720 = ~n5679 & n5719;
  assign n5721 = n5681 & ~n5720;
  assign n5722 = n5594 & n5707;
  assign n5723 = n5687 & n5698;
  assign n5724 = ~n5722 & ~n5723;
  assign n5725 = ~n5683 & ~n5705;
  assign n5726 = n5724 & n5725;
  assign n5727 = n5686 & ~n5726;
  assign n5728 = n5687 & n5707;
  assign n5729 = n5719 & ~n5728;
  assign n5730 = ~n5690 & n5729;
  assign n5731 = n5704 & ~n5730;
  assign n5732 = ~n5727 & ~n5731;
  assign n5733 = ~n5721 & n5732;
  assign n5734 = n5594 & n5691;
  assign n5735 = n5734 ^ n5511;
  assign n5736 = n5734 ^ n5704;
  assign n5737 = n5736 ^ n5704;
  assign n5738 = n5689 & n5698;
  assign n5739 = ~n5722 & ~n5738;
  assign n5740 = ~n5688 & n5739;
  assign n5741 = ~n5717 & n5740;
  assign n5742 = n5741 ^ n5704;
  assign n5743 = ~n5737 & n5742;
  assign n5744 = n5743 ^ n5704;
  assign n5745 = n5735 & n5744;
  assign n5746 = n5745 ^ n5511;
  assign n5747 = n5733 & ~n5746;
  assign n5748 = n5716 & n5747;
  assign n5749 = n5713 & n5748;
  assign n5750 = n5703 & n5749;
  assign n5751 = n5685 & n5750;
  assign n5752 = n5751 ^ n4908;
  assign n5753 = n5752 ^ x327;
  assign n5754 = ~n5376 & n5753;
  assign n5755 = n5076 & n5084;
  assign n5756 = n5075 & n5755;
  assign n5757 = n5031 & n5611;
  assign n5758 = ~n4987 & n5757;
  assign n5759 = ~n5756 & ~n5758;
  assign n5760 = n5037 & n5095;
  assign n5761 = ~n5105 & n5611;
  assign n5762 = ~n5760 & ~n5761;
  assign n5763 = ~n5029 & n5101;
  assign n5764 = ~n5079 & ~n5763;
  assign n5765 = n5119 & n5764;
  assign n5766 = n5765 ^ n5113;
  assign n5767 = n5115 & ~n5766;
  assign n5768 = n5767 ^ n5113;
  assign n5769 = n5108 & n5768;
  assign n5770 = n5762 & ~n5769;
  assign n5771 = n5759 & n5770;
  assign n5772 = n5771 ^ n2169;
  assign n5773 = n5772 ^ x284;
  assign n5774 = ~n4460 & ~n4465;
  assign n5775 = ~n4446 & n5774;
  assign n5776 = n4464 & ~n5775;
  assign n5777 = n4462 & n4484;
  assign n5778 = ~n4475 & n5777;
  assign n5779 = n4448 & ~n5778;
  assign n5781 = ~n4452 & n5573;
  assign n5780 = ~n4451 & n4484;
  assign n5782 = n5781 ^ n5780;
  assign n5783 = n5781 ^ n4434;
  assign n5784 = n5783 ^ n5781;
  assign n5785 = n5782 & ~n5784;
  assign n5786 = n5785 ^ n5781;
  assign n5787 = ~n4050 & ~n5786;
  assign n5788 = ~n5779 & ~n5787;
  assign n5789 = ~n5776 & n5788;
  assign n5790 = ~n4468 & ~n4486;
  assign n5791 = n4470 & n5790;
  assign n5792 = ~n4475 & n5791;
  assign n5793 = n5792 ^ n4476;
  assign n5794 = n5793 ^ n4476;
  assign n5795 = n4476 ^ n4434;
  assign n5796 = n5795 ^ n4476;
  assign n5797 = ~n5794 & n5796;
  assign n5798 = n5797 ^ n4476;
  assign n5799 = n4050 & n5798;
  assign n5800 = n5799 ^ n4476;
  assign n5801 = n5789 & ~n5800;
  assign n5802 = n4440 ^ n4435;
  assign n5803 = n4443 ^ n4440;
  assign n5804 = n5803 ^ n4443;
  assign n5805 = n4474 ^ n4443;
  assign n5806 = n5804 & ~n5805;
  assign n5807 = n5806 ^ n4443;
  assign n5808 = ~n5802 & n5807;
  assign n5809 = n5808 ^ n4435;
  assign n5810 = n5801 & ~n5809;
  assign n5811 = n5560 & n5810;
  assign n5812 = n5811 ^ n2591;
  assign n5813 = n5812 ^ x283;
  assign n5814 = n5773 & n5813;
  assign n5815 = n5232 & n5237;
  assign n5816 = n5255 & n5257;
  assign n5817 = ~n5815 & ~n5816;
  assign n5818 = n5147 ^ n5129;
  assign n5819 = n5295 ^ n5147;
  assign n5820 = n5819 ^ n5295;
  assign n5821 = n5282 & n5289;
  assign n5822 = ~n5263 & n5821;
  assign n5823 = n5822 ^ n5295;
  assign n5824 = ~n5820 & n5823;
  assign n5825 = n5824 ^ n5295;
  assign n5826 = ~n5818 & ~n5825;
  assign n5827 = ~n5293 & n5635;
  assign n5828 = ~n5237 & n5827;
  assign n5829 = n5828 ^ n5147;
  assign n5830 = n5829 ^ n5828;
  assign n5831 = ~n5244 & n5296;
  assign n5832 = n5831 ^ n5828;
  assign n5833 = n5830 & n5832;
  assign n5834 = n5833 ^ n5828;
  assign n5835 = n5818 & ~n5834;
  assign n5836 = ~n5826 & ~n5835;
  assign n5837 = n5261 & n5836;
  assign n5838 = n5817 & n5837;
  assign n5839 = n5270 & n5838;
  assign n5840 = ~n5231 & n5839;
  assign n5841 = n5629 & n5840;
  assign n5842 = n5841 ^ n1974;
  assign n5843 = n5842 ^ x282;
  assign n5844 = n4587 ^ x208;
  assign n5845 = n5171 ^ x213;
  assign n5846 = n5844 & ~n5845;
  assign n5847 = n4521 ^ x209;
  assign n5848 = ~n1383 & n2643;
  assign n5849 = ~n2607 & n2650;
  assign n5850 = ~n5848 & ~n5849;
  assign n5851 = n2597 & n2609;
  assign n5852 = ~n2610 & n2645;
  assign n5853 = n2327 & ~n5852;
  assign n5854 = ~n5851 & ~n5853;
  assign n5855 = n5850 & n5854;
  assign n5856 = n1689 & n2617;
  assign n5857 = ~n2595 & ~n2615;
  assign n5858 = n2625 & ~n5857;
  assign n5859 = ~n2601 & n2630;
  assign n5860 = ~n2643 & n5859;
  assign n5861 = n2327 & ~n5860;
  assign n5862 = ~n2610 & n4009;
  assign n5863 = n2609 & ~n5862;
  assign n5866 = n2630 & ~n2636;
  assign n5864 = ~n4012 & n5040;
  assign n5865 = ~n2601 & n5864;
  assign n5867 = n5866 ^ n5865;
  assign n5868 = n5866 ^ n1688;
  assign n5869 = n5868 ^ n5866;
  assign n5870 = n5867 & ~n5869;
  assign n5871 = n5870 ^ n5866;
  assign n5872 = ~n1383 & ~n5871;
  assign n5873 = ~n5863 & ~n5872;
  assign n5874 = ~n5861 & n5873;
  assign n5875 = n5039 & n5874;
  assign n5876 = ~n5858 & n5875;
  assign n5877 = ~n5856 & n5876;
  assign n5878 = n5855 & n5877;
  assign n5879 = ~n4047 & n5878;
  assign n5880 = n5879 ^ n2242;
  assign n5881 = n5880 ^ x211;
  assign n5882 = n5847 & ~n5881;
  assign n5883 = n5146 ^ x212;
  assign n5884 = n3094 & n3102;
  assign n5885 = n3078 & n3087;
  assign n5886 = ~n5884 & ~n5885;
  assign n5887 = ~n3074 & ~n3094;
  assign n5888 = n3092 & ~n5887;
  assign n5889 = ~n3076 & ~n3130;
  assign n5890 = n2749 & ~n5889;
  assign n5891 = ~n5888 & ~n5890;
  assign n5892 = ~n3114 & ~n3124;
  assign n5893 = n3078 & n3096;
  assign n5894 = n2749 & ~n3118;
  assign n5895 = ~n5893 & ~n5894;
  assign n5896 = n3094 & n3116;
  assign n5897 = n3080 ^ n3074;
  assign n5898 = n3094 ^ n3080;
  assign n5899 = n5898 ^ n3094;
  assign n5900 = n5889 ^ n3094;
  assign n5901 = ~n5899 & n5900;
  assign n5902 = n5901 ^ n3094;
  assign n5903 = n5897 & n5902;
  assign n5904 = n5903 ^ n3074;
  assign n5905 = ~n5896 & ~n5904;
  assign n5906 = n5895 & n5905;
  assign n5907 = n4815 & n5906;
  assign n5908 = n3089 & n5907;
  assign n5909 = ~n3099 & n5908;
  assign n5910 = ~n4532 & n5909;
  assign n5911 = ~n5892 & n5910;
  assign n5912 = n5891 & n5911;
  assign n5913 = n5886 & n5912;
  assign n5914 = n3113 & n5913;
  assign n5915 = ~n3136 & n5914;
  assign n5916 = n4525 & n5915;
  assign n5917 = n5916 ^ n2207;
  assign n5918 = n5917 ^ x210;
  assign n5919 = ~n5883 & n5918;
  assign n5920 = n5882 & n5919;
  assign n5921 = n5846 & n5920;
  assign n5922 = ~n5844 & ~n5845;
  assign n5923 = ~n5883 & ~n5918;
  assign n5924 = n5882 & n5923;
  assign n5925 = n5922 & n5924;
  assign n5926 = ~n5921 & ~n5925;
  assign n5927 = n5844 & n5845;
  assign n5928 = ~n5847 & n5881;
  assign n5929 = n5919 & n5928;
  assign n5930 = n5927 & n5929;
  assign n5931 = n5883 & ~n5918;
  assign n5932 = n5928 & n5931;
  assign n5933 = n5846 & n5932;
  assign n5934 = ~n5844 & n5845;
  assign n5935 = ~n5922 & ~n5934;
  assign n5936 = n5883 & n5918;
  assign n5937 = n5928 & n5936;
  assign n5938 = ~n5935 & n5937;
  assign n5939 = ~n5847 & ~n5881;
  assign n5940 = n5936 & n5939;
  assign n5941 = n5923 & n5928;
  assign n5942 = ~n5940 & ~n5941;
  assign n5943 = n5927 & ~n5942;
  assign n5944 = ~n5938 & ~n5943;
  assign n5945 = ~n5933 & n5944;
  assign n5946 = ~n5922 & ~n5927;
  assign n5947 = n5932 & ~n5946;
  assign n5948 = n5931 & n5939;
  assign n5949 = ~n5929 & ~n5948;
  assign n5950 = n5846 & ~n5949;
  assign n5951 = ~n5947 & ~n5950;
  assign n5952 = n5922 & n5929;
  assign n5953 = n5846 & n5937;
  assign n5954 = ~n5952 & ~n5953;
  assign n5955 = n5847 & n5881;
  assign n5956 = n5919 & n5955;
  assign n5957 = n5931 & n5955;
  assign n5958 = ~n5956 & ~n5957;
  assign n5959 = ~n5920 & n5958;
  assign n5960 = n5934 & ~n5959;
  assign n5961 = n5919 & n5939;
  assign n5962 = n5922 & n5961;
  assign n5963 = n5882 & n5936;
  assign n5964 = n5936 & n5955;
  assign n5965 = n5923 & n5955;
  assign n5966 = ~n5964 & ~n5965;
  assign n5967 = ~n5963 & n5966;
  assign n5968 = n5846 & ~n5967;
  assign n5969 = ~n5962 & ~n5968;
  assign n5970 = n5923 & n5939;
  assign n5971 = ~n5940 & ~n5970;
  assign n5972 = ~n5924 & n5971;
  assign n5973 = ~n5964 & n5972;
  assign n5974 = n5934 & ~n5973;
  assign n5975 = n5882 & n5931;
  assign n5976 = ~n5956 & ~n5963;
  assign n5977 = ~n5927 & n5976;
  assign n5978 = ~n5920 & ~n5963;
  assign n5979 = n5922 & n5956;
  assign n5980 = ~n5965 & ~n5979;
  assign n5981 = n5978 & n5980;
  assign n5982 = ~n5977 & ~n5981;
  assign n5983 = ~n5975 & ~n5982;
  assign n5984 = ~n5946 & ~n5983;
  assign n5985 = ~n5974 & ~n5984;
  assign n5986 = n5969 & n5985;
  assign n5987 = ~n5960 & n5986;
  assign n5988 = n5954 & n5987;
  assign n5989 = n5951 & n5988;
  assign n5990 = n5945 & n5989;
  assign n5991 = ~n5930 & n5990;
  assign n5992 = n5926 & n5991;
  assign n5993 = n5992 ^ n2322;
  assign n5994 = n5993 ^ x281;
  assign n5995 = ~n5843 & n5994;
  assign n5996 = n5814 & n5995;
  assign n5997 = n5843 & ~n5994;
  assign n5998 = n5814 & n5997;
  assign n5999 = ~n5996 & ~n5998;
  assign n6000 = n4704 & n4748;
  assign n6001 = n4700 & n4720;
  assign n6002 = ~n6000 & ~n6001;
  assign n6003 = n4704 & ~n5384;
  assign n6004 = ~n4706 & n4716;
  assign n6005 = n6004 ^ n4563;
  assign n6006 = n6005 ^ n6004;
  assign n6007 = ~n4720 & ~n4724;
  assign n6008 = ~n4748 & n6007;
  assign n6009 = n6008 ^ n6004;
  assign n6010 = n6006 & n6009;
  assign n6011 = n6010 ^ n6004;
  assign n6012 = ~n5388 & ~n6011;
  assign n6013 = ~n6003 & ~n6012;
  assign n6014 = n4709 & n5389;
  assign n6015 = ~n4732 & n6014;
  assign n6016 = n6015 ^ n4728;
  assign n6017 = n6016 ^ n4728;
  assign n6018 = n4728 ^ n4563;
  assign n6019 = n6018 ^ n4728;
  assign n6020 = ~n6017 & ~n6019;
  assign n6021 = n6020 ^ n4728;
  assign n6022 = n5388 & n6021;
  assign n6023 = n6022 ^ n4728;
  assign n6024 = n6013 & ~n6023;
  assign n6025 = ~n4743 & n6024;
  assign n6026 = n6002 & n6025;
  assign n6027 = n5382 & n6026;
  assign n6028 = n4737 & n6027;
  assign n6029 = n5379 & n6028;
  assign n6030 = ~n4699 & n6029;
  assign n6031 = n6030 ^ n1687;
  assign n6032 = n6031 ^ x285;
  assign n6033 = n3933 & n3950;
  assign n6034 = n3148 & n3937;
  assign n6035 = n3933 & n3935;
  assign n6036 = ~n6034 & ~n6035;
  assign n6037 = n3937 & n3950;
  assign n6038 = n3953 & n3964;
  assign n6039 = ~n6037 & ~n6038;
  assign n6040 = n3148 & n3964;
  assign n6042 = ~n3944 & ~n3991;
  assign n6041 = ~n3947 & ~n3951;
  assign n6043 = n6042 ^ n6041;
  assign n6044 = n6041 ^ n3953;
  assign n6045 = n6044 ^ n3953;
  assign n6046 = n3953 ^ n3148;
  assign n6047 = ~n6045 & ~n6046;
  assign n6048 = n6047 ^ n3953;
  assign n6049 = n6043 & ~n6048;
  assign n6050 = n6049 ^ n6042;
  assign n6051 = ~n3968 & n6050;
  assign n6052 = ~n3938 & n6051;
  assign n6053 = ~n3929 & n6052;
  assign n6054 = n3976 & ~n6053;
  assign n6055 = ~n6040 & ~n6054;
  assign n6056 = ~n3938 & n3979;
  assign n6057 = ~n3963 & n6056;
  assign n6058 = n3935 & ~n6057;
  assign n6060 = ~n3963 & ~n3977;
  assign n6059 = n3960 & ~n3970;
  assign n6061 = n6060 ^ n6059;
  assign n6062 = n6060 ^ n3950;
  assign n6063 = n6060 & n6062;
  assign n6064 = n6063 ^ n6060;
  assign n6065 = n6061 & n6064;
  assign n6066 = n6065 ^ n6063;
  assign n6067 = n6066 ^ n6060;
  assign n6068 = n6067 ^ n3950;
  assign n6069 = ~n6058 & n6068;
  assign n6070 = n6069 ^ n6058;
  assign n6071 = n6055 & ~n6070;
  assign n6072 = ~n3954 & ~n3991;
  assign n6073 = n6072 ^ n3978;
  assign n6074 = n6073 ^ n3978;
  assign n6075 = n3978 ^ n2669;
  assign n6076 = n6075 ^ n3978;
  assign n6077 = ~n6074 & ~n6076;
  assign n6078 = n6077 ^ n3978;
  assign n6079 = n3147 & n6078;
  assign n6080 = n6079 ^ n3978;
  assign n6081 = n6071 & ~n6080;
  assign n6082 = n3973 & n6081;
  assign n6083 = n6039 & n6082;
  assign n6084 = n6036 & n6083;
  assign n6085 = ~n6033 & n6084;
  assign n6086 = ~n3959 & n6085;
  assign n6087 = n6086 ^ n1382;
  assign n6088 = n6087 ^ x280;
  assign n6089 = n6032 & ~n6088;
  assign n6090 = ~n5999 & n6089;
  assign n6091 = ~n5773 & ~n5813;
  assign n6092 = n5997 & n6091;
  assign n6093 = ~n6032 & n6088;
  assign n6094 = n6092 & n6093;
  assign n6095 = n5843 & n5994;
  assign n6096 = n5814 & n6095;
  assign n6097 = n6032 & n6088;
  assign n6098 = n6096 & n6097;
  assign n6099 = n5995 & n6091;
  assign n6100 = ~n6032 & ~n6088;
  assign n6101 = n6099 & n6100;
  assign n6102 = n6089 & n6092;
  assign n6103 = ~n6101 & ~n6102;
  assign n6104 = ~n6098 & n6103;
  assign n6105 = ~n5773 & n5813;
  assign n6106 = n5995 & n6105;
  assign n6107 = n6100 & n6106;
  assign n6108 = n5773 & ~n5813;
  assign n6109 = ~n5843 & ~n5994;
  assign n6110 = n6108 & n6109;
  assign n6111 = n6105 & n6109;
  assign n6112 = ~n6110 & ~n6111;
  assign n6113 = n6089 & ~n6112;
  assign n6114 = ~n6107 & ~n6113;
  assign n6115 = n5997 & n6105;
  assign n6116 = n5814 & n6109;
  assign n6117 = ~n6092 & ~n6116;
  assign n6118 = ~n6115 & n6117;
  assign n6119 = n6097 & ~n6118;
  assign n6120 = ~n6097 & ~n6100;
  assign n6121 = n6095 & n6105;
  assign n6122 = n5995 & n6108;
  assign n6123 = ~n6121 & ~n6122;
  assign n6124 = ~n5998 & ~n6110;
  assign n6125 = n6093 & ~n6124;
  assign n6126 = n6123 & ~n6125;
  assign n6127 = n6120 & ~n6126;
  assign n6128 = n6095 & n6108;
  assign n6129 = ~n6121 & ~n6128;
  assign n6130 = ~n6106 & n6129;
  assign n6131 = ~n5996 & n6130;
  assign n6132 = n6093 & ~n6131;
  assign n6133 = n6091 & n6109;
  assign n6134 = ~n6115 & ~n6128;
  assign n6135 = ~n6133 & n6134;
  assign n6136 = ~n6116 & n6135;
  assign n6137 = ~n6096 & n6136;
  assign n6138 = n6100 & ~n6137;
  assign n6139 = ~n6132 & ~n6138;
  assign n6140 = ~n6127 & n6139;
  assign n6145 = n5997 & n6108;
  assign n6141 = n6091 & n6095;
  assign n6142 = ~n6122 & ~n6141;
  assign n6143 = ~n6111 & n6142;
  assign n6144 = ~n6099 & n6143;
  assign n6146 = n6145 ^ n6144;
  assign n6147 = n6146 ^ n6145;
  assign n6148 = n6145 ^ n6032;
  assign n6149 = n6148 ^ n6145;
  assign n6150 = ~n6147 & n6149;
  assign n6151 = n6150 ^ n6145;
  assign n6152 = n6088 & n6151;
  assign n6153 = n6152 ^ n6145;
  assign n6154 = n6140 & ~n6153;
  assign n6155 = ~n6119 & n6154;
  assign n6156 = n6114 & n6155;
  assign n6157 = n6104 & n6156;
  assign n6158 = ~n6094 & n6157;
  assign n6159 = ~n6090 & n6158;
  assign n6160 = n6159 ^ n5070;
  assign n6161 = n6160 ^ x324;
  assign n6162 = ~n5265 & n5266;
  assign n6163 = ~n5285 & ~n5293;
  assign n6164 = n5148 & ~n6163;
  assign n6165 = ~n6162 & ~n6164;
  assign n6166 = ~n5234 & n5288;
  assign n6167 = n5255 & ~n6166;
  assign n6168 = ~n5250 & ~n5651;
  assign n6169 = n5637 & ~n6168;
  assign n6170 = ~n5263 & n6169;
  assign n6171 = n5265 & ~n6170;
  assign n6172 = ~n6167 & ~n6171;
  assign n6173 = n6165 & n6172;
  assign n6174 = n5817 & n6173;
  assign n6175 = n5262 & n6174;
  assign n6176 = n5254 & n6175;
  assign n6177 = n5629 & n6176;
  assign n6178 = n6177 ^ n3475;
  assign n6179 = n6178 ^ x273;
  assign n6180 = n4945 & ~n4966;
  assign n6181 = ~n4913 & ~n4946;
  assign n6182 = n4931 & ~n6181;
  assign n6183 = ~n6180 & ~n6182;
  assign n6184 = ~n4916 & n4957;
  assign n6185 = ~n4955 & n4966;
  assign n6186 = ~n4918 & n6185;
  assign n6187 = n4931 & ~n6186;
  assign n6188 = ~n6184 & ~n6187;
  assign n6189 = n4945 & n4960;
  assign n6190 = n4939 & n4970;
  assign n6191 = n5522 & n6190;
  assign n6192 = n4812 & ~n6191;
  assign n6193 = ~n4937 & ~n4955;
  assign n6194 = ~n4911 & n6193;
  assign n6195 = n4914 & ~n4918;
  assign n6196 = ~n4945 & n6195;
  assign n6197 = ~n4916 & ~n6196;
  assign n6198 = ~n6194 & n6197;
  assign n6199 = ~n4938 & ~n6197;
  assign n6200 = ~n4965 & n6199;
  assign n6201 = n4950 & ~n6200;
  assign n6202 = ~n6198 & ~n6201;
  assign n6203 = ~n6192 & n6202;
  assign n6204 = ~n6189 & n6203;
  assign n6205 = n6188 & n6204;
  assign n6206 = ~n4928 & n6205;
  assign n6207 = n6183 & n6206;
  assign n6208 = n5515 & n6207;
  assign n6209 = n6208 ^ n2873;
  assign n6210 = n6209 ^ x268;
  assign n6211 = ~n6179 & n6210;
  assign n6212 = n5456 & n5486;
  assign n6213 = ~n5484 & ~n5496;
  assign n6214 = n6212 & ~n6213;
  assign n6215 = n5432 & n5457;
  assign n6216 = n5448 & n5486;
  assign n6217 = ~n6215 & ~n6216;
  assign n6218 = ~n5454 & ~n5484;
  assign n6219 = ~n6217 & ~n6218;
  assign n6220 = ~n5460 & ~n5485;
  assign n6221 = n5454 & ~n6220;
  assign n6222 = ~n5491 & n5496;
  assign n6223 = ~n6221 & ~n6222;
  assign n6224 = ~n6219 & n6223;
  assign n6225 = n5479 ^ n5453;
  assign n6226 = n6225 ^ n5479;
  assign n6227 = n5494 ^ n5479;
  assign n6228 = n6226 & ~n6227;
  assign n6229 = n6228 ^ n5479;
  assign n6230 = ~n5452 & ~n6229;
  assign n6231 = n6224 & ~n6230;
  assign n6232 = n5471 & n6231;
  assign n6233 = ~n6214 & n6232;
  assign n6234 = n6233 ^ n3411;
  assign n6235 = n6234 ^ x272;
  assign n6236 = n5927 & n5937;
  assign n6237 = ~n5930 & ~n6236;
  assign n6238 = ~n5937 & ~n5963;
  assign n6239 = n5934 & ~n6238;
  assign n6240 = ~n5957 & ~n5964;
  assign n6241 = n5846 & ~n6240;
  assign n6242 = ~n5924 & ~n5965;
  assign n6243 = ~n5963 & n6242;
  assign n6244 = n5927 & ~n6243;
  assign n6245 = ~n6241 & ~n6244;
  assign n6246 = ~n5932 & ~n5941;
  assign n6247 = ~n5975 & n6246;
  assign n6248 = n5934 & ~n6247;
  assign n6249 = ~n5920 & n5966;
  assign n6250 = ~n5948 & n6249;
  assign n6251 = n5922 & ~n6250;
  assign n6252 = ~n6248 & ~n6251;
  assign n6253 = n6245 & n6252;
  assign n6254 = n5845 ^ n5844;
  assign n6255 = n5971 ^ n5961;
  assign n6256 = n6254 & ~n6255;
  assign n6257 = n6256 ^ n5961;
  assign n6258 = n6253 & ~n6257;
  assign n6259 = ~n6239 & n6258;
  assign n6260 = n6237 & n6259;
  assign n6261 = n5951 & n6260;
  assign n6262 = n5926 & n6261;
  assign n6263 = ~n5956 & n6262;
  assign n6264 = n6263 ^ n2701;
  assign n6265 = n6264 ^ x269;
  assign n6266 = ~n6235 & n6265;
  assign n6267 = n5037 & n5604;
  assign n6268 = n5033 & n5595;
  assign n6269 = ~n5073 & ~n5098;
  assign n6270 = ~n5078 & n6269;
  assign n6271 = n5084 & ~n6270;
  assign n6272 = ~n6268 & ~n6271;
  assign n6273 = ~n6267 & n6272;
  assign n6274 = ~n5609 & n5611;
  assign n6275 = n5034 & n5616;
  assign n6276 = ~n6274 & ~n6275;
  assign n6277 = n6273 & n6276;
  assign n6278 = n5759 & n6277;
  assign n6279 = n6278 ^ n4183;
  assign n6280 = n6279 ^ x270;
  assign n6281 = ~n4460 & ~n4475;
  assign n6282 = n4443 & ~n6281;
  assign n6283 = ~n4482 & n5790;
  assign n6284 = n4444 & ~n6283;
  assign n6285 = ~n6282 & ~n6284;
  assign n6286 = n4446 ^ n4434;
  assign n6287 = n6286 ^ n4446;
  assign n6288 = n4440 & n4477;
  assign n6289 = ~n4452 & n6288;
  assign n6290 = n6289 ^ n4446;
  assign n6291 = n6290 ^ n4446;
  assign n6292 = ~n6287 & ~n6291;
  assign n6293 = n6292 ^ n4446;
  assign n6294 = n4050 & n6293;
  assign n6295 = n6294 ^ n4446;
  assign n6296 = n6285 & ~n6295;
  assign n6297 = n4435 & n4476;
  assign n6298 = ~n4451 & n4462;
  assign n6299 = n4464 & ~n6298;
  assign n6300 = ~n4451 & n5581;
  assign n6301 = ~n4443 & n6300;
  assign n6302 = ~n4451 & n4483;
  assign n6303 = n4435 & ~n6302;
  assign n6304 = n5577 & ~n6303;
  assign n6305 = n5790 & n6304;
  assign n6306 = ~n6301 & ~n6305;
  assign n6307 = ~n4444 & n6306;
  assign n6308 = ~n6299 & ~n6307;
  assign n6309 = ~n6297 & n6308;
  assign n6310 = n6296 & n6309;
  assign n6311 = n5565 & n6310;
  assign n6312 = n6311 ^ n4222;
  assign n6313 = n6312 ^ x271;
  assign n6314 = ~n6280 & ~n6313;
  assign n6315 = n6266 & n6314;
  assign n6316 = n6211 & n6315;
  assign n6317 = ~n6280 & n6313;
  assign n6318 = n6235 & n6317;
  assign n6319 = n6265 & n6318;
  assign n6320 = n6211 & n6319;
  assign n6321 = n6235 & n6280;
  assign n6322 = ~n6313 & n6321;
  assign n6323 = ~n6265 & n6322;
  assign n6324 = n6179 & ~n6210;
  assign n6325 = n6323 & n6324;
  assign n6326 = ~n6320 & ~n6325;
  assign n6327 = ~n6316 & n6326;
  assign n6328 = n6179 & n6210;
  assign n6329 = ~n6179 & ~n6210;
  assign n6330 = ~n6328 & ~n6329;
  assign n6331 = n6235 & n6314;
  assign n6332 = n6265 & n6331;
  assign n6333 = n6266 & n6313;
  assign n6334 = n6280 & n6333;
  assign n6335 = n6265 & n6322;
  assign n6336 = ~n6334 & ~n6335;
  assign n6337 = ~n6332 & n6336;
  assign n6338 = ~n6330 & ~n6337;
  assign n6339 = ~n6280 & n6333;
  assign n6340 = n6313 & n6321;
  assign n6341 = n6265 & n6340;
  assign n6342 = ~n6339 & ~n6341;
  assign n6343 = n6280 & ~n6313;
  assign n6344 = n6266 & ~n6343;
  assign n6345 = n6342 & ~n6344;
  assign n6346 = n6324 & ~n6345;
  assign n6347 = ~n6338 & ~n6346;
  assign n6348 = ~n6235 & n6314;
  assign n6349 = ~n6265 & n6348;
  assign n6350 = n6266 & n6343;
  assign n6351 = ~n6265 & n6313;
  assign n6352 = ~n6280 & n6351;
  assign n6353 = n6235 & n6352;
  assign n6354 = n6280 & n6351;
  assign n6355 = ~n6235 & n6354;
  assign n6356 = ~n6353 & ~n6355;
  assign n6357 = ~n6350 & n6356;
  assign n6358 = ~n6349 & n6357;
  assign n6359 = n6328 & ~n6358;
  assign n6360 = ~n6235 & n6343;
  assign n6361 = ~n6265 & n6360;
  assign n6362 = ~n6265 & n6331;
  assign n6363 = ~n6355 & ~n6362;
  assign n6364 = ~n6323 & n6363;
  assign n6365 = ~n6361 & n6364;
  assign n6366 = n6211 & ~n6365;
  assign n6367 = ~n6359 & ~n6366;
  assign n6368 = n6347 & n6367;
  assign n6369 = ~n6235 & n6352;
  assign n6370 = ~n6361 & ~n6362;
  assign n6371 = ~n6369 & n6370;
  assign n6372 = n6371 ^ n6179;
  assign n6373 = n6372 ^ n6371;
  assign n6374 = n6321 & n6351;
  assign n6375 = ~n6341 & ~n6374;
  assign n6376 = ~n6349 & ~n6353;
  assign n6377 = n6375 & n6376;
  assign n6378 = ~n6369 & n6377;
  assign n6379 = n6378 ^ n6371;
  assign n6380 = ~n6373 & n6379;
  assign n6381 = n6380 ^ n6371;
  assign n6382 = ~n6210 & ~n6381;
  assign n6383 = n6368 & ~n6382;
  assign n6384 = n6319 ^ n6179;
  assign n6385 = n6384 ^ n6319;
  assign n6386 = n6342 ^ n6319;
  assign n6387 = ~n6385 & ~n6386;
  assign n6388 = n6387 ^ n6319;
  assign n6389 = n6210 & n6388;
  assign n6390 = n6383 & ~n6389;
  assign n6391 = n6327 & n6390;
  assign n6392 = n6391 ^ n4810;
  assign n6393 = n6392 ^ x326;
  assign n6394 = n5621 ^ x303;
  assign n6395 = n5306 ^ x298;
  assign n6396 = n6394 & ~n6395;
  assign n6397 = ~n5948 & ~n5961;
  assign n6398 = n5846 & ~n6397;
  assign n6399 = n5922 & ~n6246;
  assign n6400 = ~n6398 & ~n6399;
  assign n6401 = ~n5940 & n5978;
  assign n6402 = ~n5964 & n6401;
  assign n6403 = n5922 & ~n6402;
  assign n6404 = n5966 & ~n5975;
  assign n6405 = n5972 & n6404;
  assign n6406 = n5927 & ~n6405;
  assign n6407 = ~n6403 & ~n6406;
  assign n6408 = ~n5941 & n5949;
  assign n6409 = n6408 ^ n5845;
  assign n6410 = n6409 ^ n6408;
  assign n6411 = n5958 & n6242;
  assign n6412 = n6411 ^ n6408;
  assign n6413 = ~n6410 & n6412;
  assign n6414 = n6413 ^ n6408;
  assign n6415 = n6254 & ~n6414;
  assign n6416 = n6407 & ~n6415;
  assign n6417 = ~n6239 & n6416;
  assign n6418 = ~n5960 & n6417;
  assign n6419 = n5954 & n6418;
  assign n6420 = n6237 & n6419;
  assign n6421 = n6400 & n6420;
  assign n6422 = n5926 & n6421;
  assign n6423 = n6422 ^ n4074;
  assign n6424 = n6423 ^ x301;
  assign n6425 = n5509 ^ x302;
  assign n6426 = n6424 & ~n6425;
  assign n6427 = n4501 ^ x299;
  assign n6428 = n3929 & n3953;
  assign n6429 = n3148 & ~n3960;
  assign n6430 = ~n6428 & ~n6429;
  assign n6431 = n2669 & n3944;
  assign n6432 = n3947 & n3976;
  assign n6433 = ~n6431 & ~n6432;
  assign n6434 = n3950 & n3968;
  assign n6435 = n3953 & n3970;
  assign n6436 = ~n3929 & ~n3978;
  assign n6437 = n3950 & ~n6436;
  assign n6438 = ~n3944 & n3965;
  assign n6439 = n3935 & ~n6438;
  assign n6440 = ~n6437 & ~n6439;
  assign n6441 = n3147 ^ n2669;
  assign n6442 = n3939 & ~n3964;
  assign n6443 = n6442 ^ n3147;
  assign n6444 = n6443 ^ n6442;
  assign n6445 = ~n3958 & ~n3991;
  assign n6446 = n6445 ^ n6442;
  assign n6447 = n6444 & n6446;
  assign n6448 = n6447 ^ n6442;
  assign n6449 = ~n6441 & ~n6448;
  assign n6450 = n6440 & ~n6449;
  assign n6451 = n3967 & n6450;
  assign n6452 = ~n3959 & n6451;
  assign n6453 = ~n6435 & n6452;
  assign n6454 = ~n6434 & n6453;
  assign n6455 = n6433 & n6454;
  assign n6456 = n3941 & n6455;
  assign n6457 = n6036 & n6456;
  assign n6458 = n6430 & n6457;
  assign n6459 = ~n6033 & n6458;
  assign n6460 = ~n3951 & n6459;
  assign n6461 = n6460 ^ n4105;
  assign n6462 = n6461 ^ x300;
  assign n6463 = ~n6427 & n6462;
  assign n6464 = n6426 & n6463;
  assign n6465 = ~n6424 & n6425;
  assign n6466 = n6463 & n6465;
  assign n6467 = ~n6464 & ~n6466;
  assign n6468 = n6396 & ~n6467;
  assign n6469 = ~n6394 & ~n6395;
  assign n6470 = n6424 & n6425;
  assign n6471 = n6427 & n6462;
  assign n6472 = n6470 & n6471;
  assign n6473 = n6427 & ~n6462;
  assign n6474 = n6426 & n6473;
  assign n6475 = ~n6472 & ~n6474;
  assign n6476 = n6469 & ~n6475;
  assign n6477 = ~n6468 & ~n6476;
  assign n6478 = n6470 & n6473;
  assign n6479 = n6469 & n6478;
  assign n6480 = ~n6394 & n6395;
  assign n6481 = n6465 & n6473;
  assign n6482 = n6465 & n6471;
  assign n6483 = ~n6474 & ~n6482;
  assign n6484 = ~n6481 & n6483;
  assign n6485 = n6480 & ~n6484;
  assign n6486 = ~n6479 & ~n6485;
  assign n6487 = ~n6424 & ~n6425;
  assign n6492 = n6471 & n6487;
  assign n6488 = n6463 & n6487;
  assign n6489 = ~n6427 & ~n6462;
  assign n6490 = n6465 & n6489;
  assign n6491 = ~n6488 & ~n6490;
  assign n6493 = n6492 ^ n6491;
  assign n6494 = n6493 ^ n6492;
  assign n6495 = n6492 ^ n6394;
  assign n6496 = n6495 ^ n6492;
  assign n6497 = ~n6494 & n6496;
  assign n6498 = n6497 ^ n6492;
  assign n6499 = ~n6395 & n6498;
  assign n6500 = n6499 ^ n6492;
  assign n6501 = n6486 & ~n6500;
  assign n6502 = n6395 ^ n6394;
  assign n6503 = n6473 & n6487;
  assign n6504 = ~n6502 & n6503;
  assign n6505 = n6394 & n6395;
  assign n6506 = n6426 & n6471;
  assign n6507 = ~n6472 & ~n6506;
  assign n6508 = n6505 & ~n6507;
  assign n6509 = n6469 & ~n6491;
  assign n6510 = n6463 & n6470;
  assign n6511 = n6480 & n6510;
  assign n6512 = n6396 & n6472;
  assign n6513 = ~n6511 & ~n6512;
  assign n6514 = ~n6467 & n6469;
  assign n6515 = n6487 & n6489;
  assign n6516 = ~n6464 & ~n6490;
  assign n6517 = ~n6515 & n6516;
  assign n6518 = n6480 & ~n6517;
  assign n6519 = ~n6514 & ~n6518;
  assign n6520 = ~n6478 & n6483;
  assign n6521 = n6396 & ~n6520;
  assign n6522 = n6470 & n6489;
  assign n6523 = n6426 & n6489;
  assign n6524 = ~n6466 & ~n6515;
  assign n6525 = ~n6523 & n6524;
  assign n6526 = ~n6522 & n6525;
  assign n6527 = n6505 & ~n6526;
  assign n6528 = ~n6521 & ~n6527;
  assign n6529 = n6519 & n6528;
  assign n6530 = n6513 & n6529;
  assign n6531 = ~n6509 & n6530;
  assign n6532 = ~n6508 & n6531;
  assign n6533 = ~n6504 & n6532;
  assign n6534 = n6501 & n6533;
  assign n6535 = n6477 & n6534;
  assign n6536 = n6535 ^ n5028;
  assign n6537 = n6536 ^ x325;
  assign n6538 = n6393 & n6537;
  assign n6539 = ~n6161 & n6538;
  assign n6540 = n6264 ^ x267;
  assign n6541 = n5592 ^ x262;
  assign n6542 = n6540 & ~n6541;
  assign n6543 = n3944 & ~n3976;
  assign n6544 = n2669 & ~n3965;
  assign n6545 = ~n6543 & ~n6544;
  assign n6546 = n3976 & n3978;
  assign n6547 = ~n3951 & ~n3963;
  assign n6548 = n3953 & ~n6547;
  assign n6549 = ~n6546 & ~n6548;
  assign n6550 = ~n3958 & ~n3977;
  assign n6551 = n3935 & ~n6550;
  assign n6552 = ~n3947 & n6072;
  assign n6553 = ~n3147 & ~n6552;
  assign n6554 = ~n6551 & ~n6553;
  assign n6555 = n6549 & n6554;
  assign n6556 = n6545 & n6555;
  assign n6557 = ~n6035 & n6556;
  assign n6558 = n6039 & n6557;
  assign n6559 = n6430 & n6558;
  assign n6560 = n3942 & n6559;
  assign n6561 = n3974 & n6560;
  assign n6562 = ~n6033 & n6561;
  assign n6563 = n6562 ^ n3069;
  assign n6564 = n6563 ^ x264;
  assign n6565 = n6209 ^ x266;
  assign n6566 = n5408 ^ x263;
  assign n6567 = n5454 & n5458;
  assign n6568 = n5454 & n5487;
  assign n6569 = n5464 & ~n5484;
  assign n6570 = ~n6568 & ~n6569;
  assign n6571 = ~n5461 & n5474;
  assign n6572 = ~n5454 & ~n5474;
  assign n6573 = n5450 & ~n6572;
  assign n6574 = n5484 & n5488;
  assign n6575 = n5459 & ~n6213;
  assign n6576 = n5446 & n6575;
  assign n6577 = ~n6574 & ~n6576;
  assign n6578 = n5460 & n5496;
  assign n6579 = ~n5465 & ~n5478;
  assign n6580 = ~n5485 & n6579;
  assign n6581 = n6580 ^ n5484;
  assign n6582 = n6581 ^ n6580;
  assign n6583 = ~n5472 & ~n5476;
  assign n6584 = ~n5496 & n6583;
  assign n6585 = ~n5488 & n6572;
  assign n6586 = ~n5485 & n6585;
  assign n6587 = ~n6584 & ~n6586;
  assign n6588 = ~n6216 & ~n6587;
  assign n6589 = n6588 ^ n6580;
  assign n6590 = ~n6582 & n6589;
  assign n6591 = n6590 ^ n6580;
  assign n6592 = ~n6578 & n6591;
  assign n6593 = n6577 & n6592;
  assign n6594 = ~n6573 & n6593;
  assign n6595 = ~n6571 & n6594;
  assign n6596 = n6570 & n6595;
  assign n6597 = ~n6567 & n6596;
  assign n6598 = ~n6214 & n6597;
  assign n6599 = n6598 ^ n3033;
  assign n6600 = n6599 ^ x265;
  assign n6601 = ~n6566 & ~n6600;
  assign n6602 = n6565 & n6601;
  assign n6603 = n6564 & n6602;
  assign n6604 = ~n6564 & ~n6565;
  assign n6605 = ~n6566 & n6604;
  assign n6606 = ~n6600 & n6605;
  assign n6607 = ~n6603 & ~n6606;
  assign n6608 = n6542 & ~n6607;
  assign n6609 = n6541 ^ n6540;
  assign n6610 = n6566 & ~n6600;
  assign n6611 = n6564 & ~n6565;
  assign n6612 = n6610 & n6611;
  assign n6613 = n6612 ^ n6541;
  assign n6614 = n6613 ^ n6612;
  assign n6615 = n6566 & n6600;
  assign n6616 = n6604 & n6615;
  assign n6617 = n6565 & n6610;
  assign n6618 = n6564 & n6617;
  assign n6619 = ~n6616 & ~n6618;
  assign n6620 = n6619 ^ n6612;
  assign n6621 = ~n6614 & ~n6620;
  assign n6622 = n6621 ^ n6612;
  assign n6623 = ~n6609 & n6622;
  assign n6624 = ~n6608 & ~n6623;
  assign n6625 = n6541 & n6618;
  assign n6626 = n6540 & n6541;
  assign n6627 = ~n6564 & n6617;
  assign n6628 = ~n6616 & ~n6627;
  assign n6629 = n6626 & ~n6628;
  assign n6630 = ~n6625 & ~n6629;
  assign n6631 = ~n6540 & ~n6541;
  assign n6632 = n6611 & n6615;
  assign n6633 = ~n6627 & ~n6632;
  assign n6634 = n6631 & ~n6633;
  assign n6635 = ~n6566 & n6600;
  assign n6636 = n6565 & n6635;
  assign n6637 = ~n6564 & n6636;
  assign n6638 = n6600 & n6605;
  assign n6639 = ~n6637 & ~n6638;
  assign n6640 = n6542 & ~n6639;
  assign n6641 = n6611 & n6635;
  assign n6642 = n6626 & n6641;
  assign n6643 = ~n6540 & n6541;
  assign n6644 = ~n6607 & n6643;
  assign n6645 = ~n6642 & ~n6644;
  assign n6646 = n6564 & n6636;
  assign n6647 = n6626 & n6646;
  assign n6648 = n6643 & n6646;
  assign n6649 = n6542 & ~n6628;
  assign n6650 = ~n6648 & ~n6649;
  assign n6651 = ~n6564 & n6602;
  assign n6652 = ~n6641 & ~n6651;
  assign n6653 = n6631 & ~n6652;
  assign n6654 = n6601 & n6611;
  assign n6655 = ~n6637 & ~n6654;
  assign n6656 = n6626 & ~n6655;
  assign n6657 = ~n6646 & ~n6654;
  assign n6658 = n6631 & ~n6657;
  assign n6659 = n6565 & n6615;
  assign n6660 = n6564 & n6659;
  assign n6661 = ~n6612 & ~n6660;
  assign n6662 = n6542 & ~n6661;
  assign n6663 = ~n6564 & n6659;
  assign n6664 = ~n6632 & ~n6663;
  assign n6665 = ~n6565 & n6610;
  assign n6666 = ~n6564 & n6665;
  assign n6667 = ~n6638 & ~n6666;
  assign n6668 = n6664 & n6667;
  assign n6669 = n6643 & ~n6668;
  assign n6670 = ~n6662 & ~n6669;
  assign n6671 = ~n6658 & n6670;
  assign n6672 = ~n6656 & n6671;
  assign n6673 = ~n6653 & n6672;
  assign n6674 = n6650 & n6673;
  assign n6675 = ~n6647 & n6674;
  assign n6676 = n6645 & n6675;
  assign n6677 = ~n6640 & n6676;
  assign n6678 = ~n6634 & n6677;
  assign n6679 = n6630 & n6678;
  assign n6680 = n6624 & n6679;
  assign n6681 = n6680 ^ n3146;
  assign n6682 = n6681 ^ x323;
  assign n6683 = ~n6393 & ~n6537;
  assign n6684 = n6683 ^ n6537;
  assign n6685 = n6684 ^ n6683;
  assign n6686 = n6683 ^ n6161;
  assign n6687 = n6686 ^ n6683;
  assign n6688 = n6685 & n6687;
  assign n6689 = n6688 ^ n6683;
  assign n6690 = n6682 & n6689;
  assign n6691 = n6690 ^ n6683;
  assign n6692 = ~n6539 & ~n6691;
  assign n6693 = n6161 & ~n6537;
  assign n6694 = n6393 & n6693;
  assign n6695 = n6682 & n6694;
  assign n6696 = ~n6161 & ~n6537;
  assign n6697 = n6393 & ~n6682;
  assign n6698 = n6696 & n6697;
  assign n6699 = ~n6695 & ~n6698;
  assign n6700 = n6692 & n6699;
  assign n6701 = n5754 & n6700;
  assign n6702 = ~n5376 & ~n5753;
  assign n6703 = n6161 & n6537;
  assign n6704 = ~n6393 & n6703;
  assign n6705 = ~n6682 & n6704;
  assign n6706 = n6537 & n6682;
  assign n6707 = ~n6393 & n6706;
  assign n6708 = ~n6161 & n6707;
  assign n6709 = ~n6705 & ~n6708;
  assign n6710 = ~n6393 & n6696;
  assign n6711 = n6539 & n6682;
  assign n6712 = ~n6710 & ~n6711;
  assign n6713 = n6693 & n6697;
  assign n6714 = n6712 & ~n6713;
  assign n6715 = n6709 & n6714;
  assign n6716 = n6699 & n6715;
  assign n6717 = n6702 & ~n6716;
  assign n6718 = ~n6701 & ~n6717;
  assign n6719 = n5376 & n5753;
  assign n6720 = n6537 ^ n6161;
  assign n6721 = n6720 ^ n6161;
  assign n6722 = n6537 ^ n6393;
  assign n6723 = n6722 ^ n6161;
  assign n6724 = n6723 ^ n6161;
  assign n6725 = ~n6721 & n6724;
  assign n6726 = n6725 ^ n6161;
  assign n6727 = ~n6682 & n6726;
  assign n6728 = n6727 ^ n6722;
  assign n6729 = n6719 & ~n6728;
  assign n6730 = n5376 & ~n5753;
  assign n6731 = n6161 & n6538;
  assign n6732 = ~n6393 & n6693;
  assign n6733 = ~n6731 & ~n6732;
  assign n6734 = n6682 & ~n6733;
  assign n6736 = ~n6161 & ~n6682;
  assign n6735 = n6696 ^ n6682;
  assign n6737 = n6736 ^ n6735;
  assign n6738 = n6393 & ~n6737;
  assign n6739 = n6738 ^ n6736;
  assign n6740 = ~n6734 & ~n6739;
  assign n6741 = n6730 & ~n6740;
  assign n6742 = ~n6729 & ~n6741;
  assign n6743 = n6718 & n6742;
  assign n6744 = n6743 ^ n5127;
  assign n6745 = n6744 ^ x390;
  assign n6746 = n6392 ^ x328;
  assign n6747 = n6396 & n6492;
  assign n6748 = n6513 & ~n6747;
  assign n6749 = n6505 & ~n6524;
  assign n6750 = ~n6488 & ~n6522;
  assign n6751 = n6396 & ~n6750;
  assign n6752 = ~n6749 & ~n6751;
  assign n6753 = n6488 & n6505;
  assign n6754 = ~n6467 & n6480;
  assign n6755 = ~n6753 & ~n6754;
  assign n6756 = ~n6396 & n6523;
  assign n6757 = ~n6478 & ~n6506;
  assign n6758 = ~n6482 & ~n6522;
  assign n6759 = n6757 & n6758;
  assign n6760 = ~n6503 & n6759;
  assign n6761 = n6469 & ~n6760;
  assign n6762 = n6483 & ~n6510;
  assign n6763 = ~n6503 & n6762;
  assign n6764 = n6396 & ~n6763;
  assign n6765 = ~n6464 & n6757;
  assign n6766 = n6505 & ~n6765;
  assign n6767 = ~n6480 & ~n6481;
  assign n6768 = ~n6481 & ~n6503;
  assign n6769 = n6475 & n6768;
  assign n6770 = ~n6767 & ~n6769;
  assign n6771 = ~n6766 & ~n6770;
  assign n6772 = n6395 & ~n6771;
  assign n6773 = ~n6764 & ~n6772;
  assign n6774 = ~n6761 & n6773;
  assign n6775 = ~n6756 & n6774;
  assign n6776 = n6755 & n6775;
  assign n6777 = n6752 & n6776;
  assign n6778 = ~n6509 & n6777;
  assign n6779 = n6748 & n6778;
  assign n6780 = n6779 ^ n4171;
  assign n6781 = n6780 ^ x333;
  assign n6782 = ~n6746 & ~n6781;
  assign n6783 = n6234 ^ x274;
  assign n6784 = n5993 ^ x279;
  assign n6785 = n6783 & n6784;
  assign n6786 = n6178 ^ x275;
  assign n6787 = ~n4766 & n4957;
  assign n6788 = ~n4923 & n4970;
  assign n6789 = n4945 & ~n6788;
  assign n6790 = ~n6787 & ~n6789;
  assign n6791 = n4941 & n5513;
  assign n6792 = n4950 & ~n6791;
  assign n6793 = n5523 & n6193;
  assign n6794 = n4812 & ~n6793;
  assign n6795 = n5522 & n6194;
  assign n6796 = ~n4951 & n6795;
  assign n6797 = n4931 & ~n6796;
  assign n6798 = ~n6794 & ~n6797;
  assign n6799 = ~n6792 & n6798;
  assign n6800 = n6790 & n6799;
  assign n6801 = n6183 & n6800;
  assign n6802 = n4929 & n6801;
  assign n6803 = ~n4954 & n6802;
  assign n6804 = n6803 ^ n3441;
  assign n6805 = n6804 ^ x276;
  assign n6806 = n6087 ^ x278;
  assign n6807 = n6805 & n6806;
  assign n6808 = ~n6786 & n6807;
  assign n6809 = n4732 & ~n5388;
  assign n6810 = n4727 & ~n4745;
  assign n6811 = ~n6809 & ~n6810;
  assign n6812 = n4700 & ~n4725;
  assign n6813 = ~n4734 & n5389;
  assign n6814 = n4704 & ~n6813;
  assign n6815 = ~n6812 & ~n6814;
  assign n6816 = ~n4713 & ~n4715;
  assign n6817 = n4564 & ~n6816;
  assign n6818 = ~n4706 & ~n4728;
  assign n6819 = n4564 & ~n6818;
  assign n6820 = ~n4714 & ~n4741;
  assign n6821 = n4700 & ~n6820;
  assign n6822 = ~n6819 & ~n6821;
  assign n6823 = n4727 & ~n5383;
  assign n6824 = ~n4697 & n4729;
  assign n6825 = n4704 & ~n6824;
  assign n6826 = ~n6823 & ~n6825;
  assign n6827 = n6822 & n6826;
  assign n6828 = n5379 & n6827;
  assign n6829 = ~n4699 & n6828;
  assign n6830 = ~n6817 & n6829;
  assign n6831 = n6815 & n6830;
  assign n6832 = n6811 & n6831;
  assign n6833 = n6002 & n6832;
  assign n6834 = n4740 & n6833;
  assign n6835 = n6834 ^ n3503;
  assign n6836 = n6835 ^ x277;
  assign n6837 = n6786 & n6836;
  assign n6838 = ~n6806 & n6837;
  assign n6839 = n6805 & n6838;
  assign n6840 = ~n6808 & ~n6839;
  assign n6841 = ~n6786 & ~n6806;
  assign n6842 = ~n6805 & n6841;
  assign n6843 = n6805 & n6841;
  assign n6844 = ~n6836 & n6843;
  assign n6845 = n6836 ^ n6806;
  assign n6846 = n6786 & ~n6845;
  assign n6847 = ~n6805 & n6846;
  assign n6848 = ~n6844 & ~n6847;
  assign n6849 = ~n6842 & n6848;
  assign n6850 = n6840 & n6849;
  assign n6851 = n6785 & ~n6850;
  assign n6852 = ~n6783 & n6784;
  assign n6853 = ~n6805 & n6838;
  assign n6854 = n6786 & n6807;
  assign n6855 = n6836 & n6841;
  assign n6856 = n6805 & n6836;
  assign n6857 = ~n6805 & ~n6836;
  assign n6858 = n6806 & n6857;
  assign n6859 = ~n6856 & ~n6858;
  assign n6860 = ~n6786 & ~n6859;
  assign n6861 = n6806 ^ n6786;
  assign n6862 = n6806 ^ n6805;
  assign n6863 = ~n6806 & ~n6862;
  assign n6864 = n6863 ^ n6806;
  assign n6865 = n6861 & ~n6864;
  assign n6866 = n6865 ^ n6863;
  assign n6867 = n6866 ^ n6806;
  assign n6868 = n6867 ^ n6805;
  assign n6869 = ~n6845 & ~n6868;
  assign n6870 = ~n6860 & ~n6869;
  assign n6871 = ~n6855 & n6870;
  assign n6872 = ~n6854 & n6871;
  assign n6873 = ~n6853 & n6872;
  assign n6874 = n6852 & ~n6873;
  assign n6875 = ~n6851 & ~n6874;
  assign n6876 = n6848 & n6870;
  assign n6877 = n6876 ^ n6783;
  assign n6878 = n6877 ^ n6876;
  assign n6879 = n6806 & n6836;
  assign n6880 = n6879 ^ n6786;
  assign n6881 = n6880 ^ n6879;
  assign n6882 = ~n6807 & ~n6836;
  assign n6883 = n6882 ^ n6879;
  assign n6884 = n6881 & n6883;
  assign n6885 = n6884 ^ n6879;
  assign n6886 = ~n6843 & ~n6885;
  assign n6887 = ~n6853 & n6886;
  assign n6888 = n6887 ^ n6876;
  assign n6889 = ~n6878 & ~n6888;
  assign n6890 = n6889 ^ n6876;
  assign n6891 = ~n6784 & n6890;
  assign n6892 = n6875 & ~n6891;
  assign n6893 = n6892 ^ n4433;
  assign n6894 = n6893 ^ x332;
  assign n6895 = n5772 ^ x286;
  assign n6896 = n4984 ^ x291;
  assign n6897 = n6895 & n6896;
  assign n6898 = n6031 ^ x287;
  assign n6899 = ~n5484 & n5485;
  assign n6900 = n6212 & ~n6218;
  assign n6901 = ~n6899 & ~n6900;
  assign n6902 = ~n5472 & ~n6216;
  assign n6903 = n5454 & ~n6902;
  assign n6904 = ~n5450 & n6217;
  assign n6905 = n5474 & ~n6904;
  assign n6906 = n5432 & n5486;
  assign n6907 = n5451 & ~n6906;
  assign n6908 = ~n5465 & n6907;
  assign n6909 = n5496 & ~n6908;
  assign n6910 = ~n6905 & ~n6909;
  assign n6911 = n5461 & n6902;
  assign n6912 = n5484 & ~n6911;
  assign n6913 = ~n5457 & ~n5474;
  assign n6914 = ~n6212 & ~n6567;
  assign n6915 = ~n5478 & n6914;
  assign n6916 = ~n5464 & n6915;
  assign n6917 = ~n6913 & ~n6916;
  assign n6918 = ~n6572 & n6917;
  assign n6919 = ~n6912 & ~n6918;
  assign n6920 = n6910 & n6919;
  assign n6921 = ~n5470 & n6920;
  assign n6922 = n6577 & n6921;
  assign n6923 = ~n6903 & n6922;
  assign n6924 = n6901 & n6923;
  assign n6925 = n6924 ^ n3851;
  assign n6926 = n6925 ^ x288;
  assign n6927 = n6898 & ~n6926;
  assign n6928 = n3998 ^ x290;
  assign n6929 = n5927 & n5961;
  assign n6930 = n5966 & n5978;
  assign n6931 = ~n5929 & n6930;
  assign n6932 = ~n5932 & n6931;
  assign n6933 = n5934 & ~n6932;
  assign n6934 = ~n6929 & ~n6933;
  assign n6935 = n5970 & n6254;
  assign n6936 = ~n5956 & n6404;
  assign n6937 = n5846 & ~n6936;
  assign n6938 = ~n5924 & ~n5964;
  assign n6939 = ~n5963 & n6938;
  assign n6940 = ~n5922 & n6939;
  assign n6941 = n5958 & n5978;
  assign n6942 = ~n5927 & n6941;
  assign n6943 = ~n6940 & ~n6942;
  assign n6944 = ~n5948 & ~n6943;
  assign n6945 = ~n5946 & ~n6944;
  assign n6946 = ~n6937 & ~n6945;
  assign n6947 = ~n6935 & n6946;
  assign n6948 = n6934 & n6947;
  assign n6949 = n6400 & n6948;
  assign n6950 = n5945 & n6949;
  assign n6951 = ~n5930 & n6950;
  assign n6952 = n6951 ^ n3819;
  assign n6953 = n6952 ^ x289;
  assign n6954 = n6928 & ~n6953;
  assign n6955 = n6927 & n6954;
  assign n6956 = n6897 & n6955;
  assign n6957 = ~n6895 & ~n6896;
  assign n6958 = n6898 & n6926;
  assign n6959 = ~n6928 & ~n6953;
  assign n6960 = n6958 & n6959;
  assign n6961 = n6957 & n6960;
  assign n6962 = ~n6956 & ~n6961;
  assign n6963 = ~n6898 & n6926;
  assign n6964 = n6928 & n6953;
  assign n6965 = n6963 & n6964;
  assign n6966 = n6959 & n6963;
  assign n6967 = ~n6965 & ~n6966;
  assign n6968 = n6897 & ~n6967;
  assign n6969 = n6895 & ~n6896;
  assign n6970 = ~n6928 & n6953;
  assign n6971 = n6958 & n6970;
  assign n6972 = n6954 & n6958;
  assign n6973 = ~n6971 & ~n6972;
  assign n6974 = n6969 & ~n6973;
  assign n6975 = ~n6968 & ~n6974;
  assign n6976 = n6958 & n6964;
  assign n6977 = n6969 & n6976;
  assign n6978 = n6897 & ~n6973;
  assign n6979 = ~n6977 & ~n6978;
  assign n6980 = n6927 & n6970;
  assign n6981 = ~n6957 & n6980;
  assign n6982 = n6963 & n6970;
  assign n6983 = ~n6898 & ~n6926;
  assign n6984 = n6954 & n6983;
  assign n6985 = ~n6982 & ~n6984;
  assign n6986 = n6897 & ~n6985;
  assign n6987 = ~n6981 & ~n6986;
  assign n6988 = n6927 & n6959;
  assign n6989 = ~n6895 & n6988;
  assign n6990 = ~n6895 & n6896;
  assign n6991 = ~n6966 & ~n6984;
  assign n6992 = ~n6976 & ~n6982;
  assign n6993 = n6927 & n6964;
  assign n6994 = n6954 & n6963;
  assign n6995 = ~n6993 & ~n6994;
  assign n6996 = n6992 & n6995;
  assign n6997 = n6991 & n6996;
  assign n6998 = n6990 & ~n6997;
  assign n6999 = ~n6989 & ~n6998;
  assign n7000 = n6957 & ~n6973;
  assign n7001 = n6964 & n6983;
  assign n7002 = n7001 ^ n6896;
  assign n7004 = n6959 & n6983;
  assign n7005 = n6970 & n6983;
  assign n7006 = ~n6965 & ~n7005;
  assign n7007 = ~n7004 & n7006;
  assign n7003 = ~n6955 & n6991;
  assign n7008 = n7007 ^ n7003;
  assign n7009 = n7007 ^ n6895;
  assign n7010 = n7009 ^ n7007;
  assign n7011 = n7008 & n7010;
  assign n7012 = n7011 ^ n7007;
  assign n7013 = n7012 ^ n7001;
  assign n7014 = n7002 & ~n7013;
  assign n7015 = n7014 ^ n7011;
  assign n7016 = n7015 ^ n7007;
  assign n7017 = n7016 ^ n6896;
  assign n7018 = ~n7001 & ~n7017;
  assign n7019 = n7018 ^ n7001;
  assign n7020 = n7019 ^ n6896;
  assign n7021 = ~n7000 & ~n7020;
  assign n7022 = n6999 & n7021;
  assign n7023 = n6987 & n7022;
  assign n7024 = n6979 & n7023;
  assign n7025 = n6975 & n7024;
  assign n7026 = n6962 & n7025;
  assign n7027 = n7026 ^ n4871;
  assign n7028 = n7027 ^ x331;
  assign n7029 = ~n6894 & ~n7028;
  assign n7030 = n5752 ^ x329;
  assign n7031 = n6643 & n6654;
  assign n7032 = ~n6638 & ~n6651;
  assign n7033 = n6626 & ~n7032;
  assign n7034 = ~n7031 & ~n7033;
  assign n7035 = n6626 & n6627;
  assign n7036 = n6643 & n6651;
  assign n7037 = ~n7035 & ~n7036;
  assign n7038 = n6541 & ~n6664;
  assign n7039 = n6639 & n6661;
  assign n7040 = n6631 & ~n7039;
  assign n7041 = ~n6603 & ~n6638;
  assign n7042 = ~n6663 & n7041;
  assign n7043 = ~n6665 & n7042;
  assign n7044 = ~n6627 & n7043;
  assign n7045 = ~n6646 & n7044;
  assign n7046 = n6542 & ~n7045;
  assign n7047 = ~n7040 & ~n7046;
  assign n7048 = ~n7038 & n7047;
  assign n7049 = n7037 & n7048;
  assign n7050 = ~n6623 & n7049;
  assign n7051 = ~n6658 & n7050;
  assign n7052 = n6641 ^ n6541;
  assign n7053 = n7052 ^ n6641;
  assign n7054 = n6641 ^ n6628;
  assign n7055 = n7053 & ~n7054;
  assign n7056 = n7055 ^ n6641;
  assign n7057 = n6609 & n7056;
  assign n7058 = n7051 & ~n7057;
  assign n7059 = n7034 & n7058;
  assign n7060 = ~n6647 & n7059;
  assign n7061 = n6645 & n7060;
  assign n7062 = n7061 ^ n4844;
  assign n7063 = n7062 ^ x330;
  assign n7064 = n7030 & ~n7063;
  assign n7065 = n7029 & n7064;
  assign n7066 = n6782 & n7065;
  assign n7067 = ~n6746 & n6781;
  assign n7068 = ~n7030 & ~n7063;
  assign n7069 = n7029 & n7068;
  assign n7070 = n7067 & n7069;
  assign n7071 = ~n7066 & ~n7070;
  assign n7072 = n6746 & n6781;
  assign n7073 = n6894 & n7028;
  assign n7074 = n7030 & n7063;
  assign n7075 = n7073 & n7074;
  assign n7076 = ~n6894 & n7028;
  assign n7077 = n7064 & n7076;
  assign n7078 = ~n7075 & ~n7077;
  assign n7079 = n7072 & ~n7078;
  assign n7080 = n6746 & ~n6781;
  assign n7081 = n7068 & n7073;
  assign n7082 = ~n7077 & ~n7081;
  assign n7083 = n7080 & ~n7082;
  assign n7084 = ~n7030 & n7063;
  assign n7085 = n7029 & n7084;
  assign n7086 = n7072 & n7085;
  assign n7087 = n7064 & n7073;
  assign n7088 = n6782 & n7087;
  assign n7089 = n7074 & n7076;
  assign n7090 = n6894 & ~n7028;
  assign n7091 = n7074 & n7090;
  assign n7092 = ~n7089 & ~n7091;
  assign n7093 = n7080 & ~n7092;
  assign n7094 = ~n7088 & ~n7093;
  assign n7095 = ~n7086 & n7094;
  assign n7096 = n7068 & n7090;
  assign n7097 = ~n7075 & ~n7096;
  assign n7098 = ~n7069 & n7097;
  assign n7099 = ~n7087 & n7098;
  assign n7100 = n7080 & ~n7099;
  assign n7101 = n7029 & n7074;
  assign n7102 = n7064 & n7090;
  assign n7103 = ~n7101 & ~n7102;
  assign n7104 = n7073 & n7084;
  assign n7105 = n7084 & n7090;
  assign n7106 = n7068 & n7076;
  assign n7107 = ~n7105 & ~n7106;
  assign n7108 = ~n7104 & n7107;
  assign n7109 = n7103 & n7108;
  assign n7110 = ~n7069 & n7109;
  assign n7111 = n6782 & ~n7110;
  assign n7112 = ~n7100 & ~n7111;
  assign n7113 = n7076 & n7084;
  assign n7114 = ~n7105 & ~n7113;
  assign n7115 = ~n7096 & n7114;
  assign n7116 = ~n7087 & ~n7101;
  assign n7117 = n7115 & n7116;
  assign n7118 = n7072 & ~n7117;
  assign n7119 = ~n7075 & n7103;
  assign n7120 = ~n7081 & n7119;
  assign n7121 = ~n7065 & n7120;
  assign n7122 = n7114 & n7121;
  assign n7123 = n7067 & ~n7122;
  assign n7124 = ~n7118 & ~n7123;
  assign n7125 = n7112 & n7124;
  assign n7126 = n7095 & n7125;
  assign n7127 = ~n7083 & n7126;
  assign n7128 = ~n7079 & n7127;
  assign n7129 = n7071 & n7128;
  assign n7130 = n7129 ^ n4984;
  assign n7131 = n7130 ^ x389;
  assign n7132 = n6745 & ~n7131;
  assign n7133 = ~n6839 & ~n6844;
  assign n7134 = n6783 & ~n6784;
  assign n7135 = ~n6805 & n6879;
  assign n7136 = n6857 ^ n6786;
  assign n7137 = n7136 ^ n6857;
  assign n7138 = n6857 ^ n6807;
  assign n7139 = n7137 & n7138;
  assign n7140 = n7139 ^ n6857;
  assign n7141 = ~n7135 & ~n7140;
  assign n7142 = n7134 & ~n7141;
  assign n7143 = n6841 & n6857;
  assign n7144 = ~n6808 & ~n7143;
  assign n7145 = n6786 & n6858;
  assign n7146 = n6836 & n6842;
  assign n7147 = ~n7145 & ~n7146;
  assign n7148 = ~n6786 & n6879;
  assign n7149 = ~n6869 & ~n7148;
  assign n7150 = n7147 & n7149;
  assign n7151 = n7144 & n7150;
  assign n7152 = n6852 & n7151;
  assign n7153 = ~n7142 & ~n7152;
  assign n7154 = ~n6783 & ~n6784;
  assign n7155 = n6807 & ~n6837;
  assign n7156 = ~n6853 & n7147;
  assign n7157 = ~n7155 & n7156;
  assign n7158 = n7154 & ~n7157;
  assign n7159 = n6785 & ~n7150;
  assign n7160 = ~n7158 & ~n7159;
  assign n7161 = n7153 & n7160;
  assign n7162 = n7133 & n7161;
  assign n7163 = n7162 ^ n4521;
  assign n7164 = n7163 ^ x351;
  assign n7165 = n6631 & ~n7041;
  assign n7166 = ~n6612 & ~n6618;
  assign n7167 = n6633 & n7166;
  assign n7168 = ~n6606 & ~n6637;
  assign n7169 = ~n6646 & n7168;
  assign n7170 = n7167 & n7169;
  assign n7171 = n6643 & ~n7170;
  assign n7172 = ~n6626 & ~n6631;
  assign n7173 = ~n6660 & ~n6666;
  assign n7174 = ~n7172 & ~n7173;
  assign n7175 = n6600 ^ n6566;
  assign n7176 = n7175 ^ n6565;
  assign n7177 = n6565 ^ n6564;
  assign n7178 = n6600 ^ n6564;
  assign n7179 = n7178 ^ n6564;
  assign n7180 = ~n7177 & ~n7179;
  assign n7181 = n7180 ^ n6564;
  assign n7182 = n7176 & n7181;
  assign n7183 = n7182 ^ n6566;
  assign n7184 = n6542 & n7183;
  assign n7185 = ~n7174 & ~n7184;
  assign n7186 = ~n7171 & n7185;
  assign n7187 = ~n7165 & n7186;
  assign n7188 = ~n6656 & n7187;
  assign n7189 = ~n6653 & n7188;
  assign n7190 = n6624 & n7189;
  assign n7191 = n7034 & n7190;
  assign n7192 = ~n6647 & n7191;
  assign n7193 = n7192 ^ n4562;
  assign n7194 = n7193 ^ x346;
  assign n7195 = ~n7164 & ~n7194;
  assign n7196 = n6990 & ~n7006;
  assign n7197 = ~n6994 & ~n7005;
  assign n7198 = n6969 & ~n7197;
  assign n7199 = ~n7196 & ~n7198;
  assign n7200 = n6897 & n7004;
  assign n7201 = n6969 & n6980;
  assign n7202 = n6897 & n7001;
  assign n7203 = ~n7201 & ~n7202;
  assign n7204 = ~n7200 & n7203;
  assign n7205 = n6897 & n6960;
  assign n7206 = ~n6972 & ~n6980;
  assign n7207 = n6990 & ~n7206;
  assign n7208 = ~n6955 & n6967;
  assign n7209 = n6957 & ~n7208;
  assign n7210 = ~n7207 & ~n7209;
  assign n7211 = ~n7205 & n7210;
  assign n7212 = ~n6895 & n6971;
  assign n7213 = n6965 & n6969;
  assign n7214 = ~n7212 & ~n7213;
  assign n7215 = n6897 & ~n6992;
  assign n7216 = n6995 & ~n7004;
  assign n7217 = n6957 & ~n7216;
  assign n7218 = ~n6969 & ~n6990;
  assign n7219 = ~n6988 & n6991;
  assign n7220 = ~n7218 & ~n7219;
  assign n7221 = ~n7217 & ~n7220;
  assign n7222 = ~n7215 & n7221;
  assign n7223 = n7214 & n7222;
  assign n7224 = n6979 & n7223;
  assign n7225 = n6962 & n7224;
  assign n7226 = n7211 & n7225;
  assign n7227 = n7204 & n7226;
  assign n7228 = n7199 & n7227;
  assign n7229 = n7228 ^ n4625;
  assign n7230 = n7229 ^ x347;
  assign n7231 = ~n6319 & ~n6334;
  assign n7232 = n6324 & ~n7231;
  assign n7233 = n6323 & n6329;
  assign n7234 = ~n6361 & ~n6374;
  assign n7235 = n6328 & ~n7234;
  assign n7236 = ~n7233 & ~n7235;
  assign n7237 = ~n6330 & n6332;
  assign n7238 = n6324 & ~n6363;
  assign n7239 = ~n7237 & ~n7238;
  assign n7240 = n6319 & ~n6330;
  assign n7241 = ~n6315 & ~n6335;
  assign n7242 = n7234 & n7241;
  assign n7243 = n6324 & ~n7242;
  assign n7244 = n6336 & n6357;
  assign n7245 = n6329 & ~n7244;
  assign n7246 = ~n6350 & ~n6369;
  assign n7247 = n6363 & n7246;
  assign n7248 = n6328 & ~n7247;
  assign n7249 = ~n7245 & ~n7248;
  assign n7250 = ~n6341 & n7241;
  assign n7251 = ~n6355 & n7250;
  assign n7252 = n6376 & n7251;
  assign n7253 = n7234 & n7252;
  assign n7254 = n6211 & ~n7253;
  assign n7255 = n7249 & ~n7254;
  assign n7256 = ~n7243 & n7255;
  assign n7257 = ~n7240 & n7256;
  assign n7258 = n7239 & n7257;
  assign n7259 = n7236 & n7258;
  assign n7260 = ~n7232 & n7259;
  assign n7261 = n7260 ^ n4661;
  assign n7262 = n7261 ^ x348;
  assign n7263 = n7230 & ~n7262;
  assign n7264 = n4503 & n5342;
  assign n7265 = n5331 & n5348;
  assign n7267 = n5325 & n5334;
  assign n7268 = ~n5352 & ~n7267;
  assign n7266 = n5346 & n5365;
  assign n7269 = n7268 ^ n7266;
  assign n7270 = n7269 ^ n7268;
  assign n7271 = n7268 ^ n4502;
  assign n7272 = n7271 ^ n7268;
  assign n7273 = ~n7270 & n7272;
  assign n7274 = n7273 ^ n7268;
  assign n7275 = ~n3999 & ~n7274;
  assign n7276 = n7275 ^ n7268;
  assign n7277 = ~n7265 & n7276;
  assign n7278 = n5343 ^ n4502;
  assign n7279 = n7278 ^ n5343;
  assign n7280 = ~n5316 & n5365;
  assign n7281 = n5332 & n7280;
  assign n7282 = ~n5329 & n7281;
  assign n7283 = n7282 ^ n5343;
  assign n7284 = ~n7279 & n7283;
  assign n7285 = n7284 ^ n5343;
  assign n7286 = n3999 & ~n7285;
  assign n7287 = n7277 & ~n7286;
  assign n7288 = ~n7264 & n7287;
  assign n7289 = n5328 & n7288;
  assign n7290 = n5321 & n7289;
  assign n7291 = n7290 ^ n4587;
  assign n7292 = n7291 ^ x350;
  assign n7293 = n5681 & n5690;
  assign n7294 = n5716 & ~n7293;
  assign n7295 = n5681 & n5692;
  assign n7296 = n5686 & n5738;
  assign n7297 = ~n7295 & ~n7296;
  assign n7298 = n5511 & n5705;
  assign n7299 = n5713 & ~n7298;
  assign n7300 = n5679 & n5686;
  assign n7301 = n5511 & n5708;
  assign n7302 = ~n7300 & ~n7301;
  assign n7303 = n5724 & ~n5734;
  assign n7304 = n5511 & ~n7303;
  assign n7305 = n5704 & ~n5741;
  assign n7306 = ~n7304 & ~n7305;
  assign n7307 = ~n5511 & ~n5704;
  assign n7308 = n5683 & ~n7307;
  assign n7309 = n5686 & n5699;
  assign n7310 = ~n7308 & ~n7309;
  assign n7311 = ~n5705 & ~n5728;
  assign n7312 = ~n5708 & n7311;
  assign n7313 = n7312 ^ n5710;
  assign n7314 = n7313 ^ n5710;
  assign n7315 = n5710 ^ n5409;
  assign n7316 = n7315 ^ n5710;
  assign n7317 = ~n7314 & ~n7316;
  assign n7318 = n7317 ^ n5710;
  assign n7319 = n5510 & n7318;
  assign n7320 = n7319 ^ n5710;
  assign n7321 = n7310 & ~n7320;
  assign n7322 = n7306 & n7321;
  assign n7323 = n7302 & n7322;
  assign n7324 = n7299 & n7323;
  assign n7325 = n7297 & n7324;
  assign n7326 = n5703 & n7325;
  assign n7327 = n7294 & n7326;
  assign n7328 = n7327 ^ n4691;
  assign n7329 = n7328 ^ x349;
  assign n7330 = ~n7292 & ~n7329;
  assign n7331 = n7263 & n7330;
  assign n7332 = n7195 & n7331;
  assign n7333 = n7164 & ~n7194;
  assign n7334 = ~n7230 & ~n7262;
  assign n7335 = ~n7292 & n7329;
  assign n7336 = n7334 & n7335;
  assign n7337 = ~n7230 & n7262;
  assign n7338 = n7292 & n7329;
  assign n7339 = n7337 & n7338;
  assign n7340 = ~n7336 & ~n7339;
  assign n7341 = n7333 & ~n7340;
  assign n7342 = ~n7332 & ~n7341;
  assign n7343 = ~n7164 & n7194;
  assign n7344 = n7331 & n7343;
  assign n7345 = ~n7292 & n7337;
  assign n7346 = n7329 & n7345;
  assign n7347 = n7292 & ~n7329;
  assign n7348 = n7334 & n7347;
  assign n7349 = ~n7346 & ~n7348;
  assign n7350 = n7333 & ~n7349;
  assign n7351 = ~n7344 & ~n7350;
  assign n7352 = n7263 & n7335;
  assign n7353 = n7195 & n7352;
  assign n7354 = n7164 & n7194;
  assign n7355 = n7230 & n7262;
  assign n7356 = n7335 & n7355;
  assign n7357 = n7347 & n7355;
  assign n7358 = ~n7356 & ~n7357;
  assign n7359 = n7354 & ~n7358;
  assign n7360 = ~n7353 & ~n7359;
  assign n7361 = n7263 & n7347;
  assign n7362 = n7333 & n7361;
  assign n7363 = ~n7340 & n7354;
  assign n7364 = ~n7362 & ~n7363;
  assign n7365 = ~n7352 & ~n7357;
  assign n7366 = n7343 & ~n7365;
  assign n7367 = ~n7329 & n7345;
  assign n7368 = n7354 & n7367;
  assign n7369 = n7354 & n7361;
  assign n7370 = n7333 & ~n7358;
  assign n7371 = ~n7369 & ~n7370;
  assign n7372 = ~n7368 & n7371;
  assign n7373 = n7331 & n7354;
  assign n7374 = n7330 & n7334;
  assign n7375 = n7338 & n7355;
  assign n7376 = n7263 & n7338;
  assign n7377 = ~n7375 & ~n7376;
  assign n7378 = n7337 & n7347;
  assign n7379 = ~n7367 & ~n7378;
  assign n7380 = n7377 & n7379;
  assign n7381 = ~n7374 & n7380;
  assign n7382 = n7195 & ~n7381;
  assign n7383 = n7334 & n7338;
  assign n7384 = n7349 & ~n7383;
  assign n7385 = ~n7378 & n7384;
  assign n7386 = ~n7375 & n7385;
  assign n7387 = n7343 & ~n7386;
  assign n7388 = ~n7382 & ~n7387;
  assign n7389 = ~n7373 & n7388;
  assign n7390 = n7194 ^ n7164;
  assign n7391 = n7330 & n7355;
  assign n7392 = n7391 ^ n7383;
  assign n7393 = n7392 ^ n7383;
  assign n7394 = n7383 ^ n7194;
  assign n7395 = n7394 ^ n7383;
  assign n7396 = n7393 & ~n7395;
  assign n7397 = n7396 ^ n7383;
  assign n7398 = n7390 & n7397;
  assign n7399 = n7398 ^ n7383;
  assign n7400 = n7389 & ~n7399;
  assign n7401 = n7372 & n7400;
  assign n7402 = ~n7366 & n7401;
  assign n7403 = n7364 & n7402;
  assign n7404 = n7360 & n7403;
  assign n7405 = n7351 & n7404;
  assign n7406 = n7342 & n7405;
  assign n7407 = n7406 ^ n4764;
  assign n7408 = n7407 ^ x391;
  assign n7409 = n6480 & n6523;
  assign n7410 = n6395 & n6515;
  assign n7411 = ~n7409 & ~n7410;
  assign n7412 = n6469 & n6510;
  assign n7413 = ~n6491 & n6505;
  assign n7414 = ~n7412 & ~n7413;
  assign n7415 = n7411 & n7414;
  assign n7416 = ~n6482 & ~n6492;
  assign n7417 = ~n6502 & ~n7416;
  assign n7418 = ~n6510 & ~n6515;
  assign n7419 = n6396 & ~n7418;
  assign n7420 = ~n7417 & ~n7419;
  assign n7421 = n6505 & ~n6757;
  assign n7422 = ~n6506 & n6768;
  assign n7423 = ~n6482 & n7422;
  assign n7424 = n6480 & ~n7423;
  assign n7425 = ~n7421 & ~n7424;
  assign n7426 = n7420 & n7425;
  assign n7427 = n6477 & n7426;
  assign n7428 = n6522 ^ n6396;
  assign n7429 = n7428 ^ n6522;
  assign n7430 = ~n6474 & ~n6481;
  assign n7431 = n7430 ^ n6522;
  assign n7432 = n7429 & ~n7431;
  assign n7433 = n7432 ^ n6522;
  assign n7434 = n7427 & ~n7433;
  assign n7435 = n7415 & n7434;
  assign n7436 = ~n6509 & n7435;
  assign n7437 = n6748 & n7436;
  assign n7438 = n7437 ^ n5171;
  assign n7439 = n7438 ^ x311;
  assign n7440 = n6328 & n6361;
  assign n7441 = ~n6211 & ~n6329;
  assign n7442 = n6369 & ~n7441;
  assign n7443 = ~n7440 & ~n7442;
  assign n7444 = ~n6332 & ~n6339;
  assign n7445 = n6324 & ~n7444;
  assign n7446 = ~n6362 & n7234;
  assign n7447 = n6211 & ~n7446;
  assign n7448 = ~n7445 & ~n7447;
  assign n7449 = ~n6353 & n6363;
  assign n7450 = ~n6330 & ~n7449;
  assign n7451 = ~n6349 & n7234;
  assign n7452 = n6324 & ~n7451;
  assign n7453 = ~n6332 & n7250;
  assign n7454 = n6211 & ~n7241;
  assign n7455 = ~n6328 & ~n7454;
  assign n7456 = ~n7453 & ~n7455;
  assign n7457 = ~n7452 & ~n7456;
  assign n7458 = n6350 ^ n6329;
  assign n7459 = n6329 ^ n6211;
  assign n7460 = n7459 ^ n6211;
  assign n7461 = n7250 ^ n6211;
  assign n7462 = n7460 & n7461;
  assign n7463 = n7462 ^ n6211;
  assign n7464 = n7458 & ~n7463;
  assign n7465 = n7464 ^ n6350;
  assign n7466 = n7457 & ~n7465;
  assign n7467 = n6326 & n7466;
  assign n7468 = ~n7450 & n7467;
  assign n7469 = n7448 & n7468;
  assign n7470 = n7443 & n7469;
  assign n7471 = ~n7232 & n7470;
  assign n7472 = n7471 ^ n5190;
  assign n7473 = n7472 ^ x312;
  assign n7474 = ~n7439 & ~n7473;
  assign n7475 = n5998 & n6100;
  assign n7476 = ~n6094 & ~n7475;
  assign n7477 = ~n6120 & n6133;
  assign n7478 = n6096 ^ n6032;
  assign n7479 = n7478 ^ n6096;
  assign n7480 = n6122 ^ n6096;
  assign n7481 = ~n7479 & n7480;
  assign n7482 = n7481 ^ n6096;
  assign n7483 = ~n6088 & n7482;
  assign n7484 = ~n7477 & ~n7483;
  assign n7485 = n6089 & n6133;
  assign n7486 = n6093 & n6111;
  assign n7487 = n6097 & n6110;
  assign n7488 = ~n7486 & ~n7487;
  assign n7489 = ~n7485 & n7488;
  assign n7490 = n6092 & n6100;
  assign n7491 = ~n6115 & ~n6145;
  assign n7492 = ~n6099 & n7491;
  assign n7493 = n6123 & n7492;
  assign n7494 = ~n5996 & n7493;
  assign n7495 = n6093 & ~n7494;
  assign n7496 = ~n7490 & ~n7495;
  assign n7497 = ~n6106 & ~n6141;
  assign n7498 = n6089 & ~n7497;
  assign n7499 = ~n6099 & ~n6106;
  assign n7500 = ~n6128 & n7499;
  assign n7501 = ~n6100 & n7500;
  assign n7502 = n6097 & ~n7499;
  assign n7503 = n6129 & ~n7502;
  assign n7504 = ~n6096 & n7503;
  assign n7505 = ~n7501 & ~n7504;
  assign n7506 = ~n6120 & n7505;
  assign n7507 = ~n7498 & ~n7506;
  assign n7508 = n7496 & n7507;
  assign n7509 = ~n6119 & n7508;
  assign n7510 = n7489 & n7509;
  assign n7511 = n6114 & n7510;
  assign n7512 = n7484 & n7511;
  assign n7513 = n7476 & n7512;
  assign n7514 = ~n6090 & n7513;
  assign n7515 = n7514 ^ n2668;
  assign n7516 = n7515 ^ x314;
  assign n7517 = n5307 ^ n5128;
  assign n7518 = n7517 ^ n4985;
  assign n7519 = n5307 ^ n4765;
  assign n7520 = n7519 ^ n4765;
  assign n7521 = n4985 ^ n4765;
  assign n7522 = n7520 & n7521;
  assign n7523 = n7522 ^ n4765;
  assign n7524 = ~n7518 & n7523;
  assign n7525 = n4503 & n7524;
  assign n7526 = n4986 & n5317;
  assign n7527 = ~n5316 & ~n7526;
  assign n7528 = n5345 & n7527;
  assign n7529 = ~n5342 & n7528;
  assign n7530 = n5331 & ~n7529;
  assign n7531 = ~n7525 & ~n7530;
  assign n7532 = ~n4503 & ~n5331;
  assign n7533 = ~n5312 & n5343;
  assign n7534 = ~n5341 & n7533;
  assign n7535 = ~n5308 & ~n5315;
  assign n7536 = n4986 & ~n7535;
  assign n7537 = n5332 & ~n7536;
  assign n7538 = ~n5318 & n7537;
  assign n7539 = ~n7534 & ~n7538;
  assign n7540 = ~n7267 & ~n7539;
  assign n7541 = n5354 & n7540;
  assign n7542 = ~n5336 & n7541;
  assign n7543 = n7532 & ~n7542;
  assign n7544 = n7531 & ~n7543;
  assign n7545 = ~n5370 & n7544;
  assign n7546 = ~n5330 & n7545;
  assign n7547 = ~n7264 & n7546;
  assign n7548 = n5328 & n7547;
  assign n7549 = n7548 ^ n5227;
  assign n7550 = n7549 ^ x313;
  assign n7551 = ~n7516 & n7550;
  assign n7552 = n7474 & n7551;
  assign n7553 = ~n5710 & n5724;
  assign n7554 = n5681 & ~n7553;
  assign n7555 = ~n5717 & n7303;
  assign n7556 = n5686 & ~n7555;
  assign n7557 = ~n7554 & ~n7556;
  assign n7558 = ~n5717 & ~n5728;
  assign n7559 = ~n7307 & ~n7558;
  assign n7560 = ~n5683 & ~n5696;
  assign n7561 = ~n5688 & n7560;
  assign n7562 = ~n5699 & n7561;
  assign n7563 = n5704 & ~n7562;
  assign n7564 = ~n7559 & ~n7563;
  assign n7565 = n7557 & n7564;
  assign n7566 = n5702 & n7565;
  assign n7567 = n7302 & n7566;
  assign n7568 = n7299 & n7567;
  assign n7569 = n7297 & n7568;
  assign n7570 = n5685 & n7569;
  assign n7571 = ~n5690 & n7570;
  assign n7572 = n7571 ^ n3784;
  assign n7573 = n7572 ^ x315;
  assign n7574 = ~n6895 & n6960;
  assign n7575 = ~n6976 & ~n6980;
  assign n7576 = ~n7001 & n7575;
  assign n7577 = ~n6988 & n7576;
  assign n7578 = n6957 & ~n7577;
  assign n7579 = ~n7574 & ~n7578;
  assign n7580 = n6926 ^ n6898;
  assign n7581 = n7580 ^ n6953;
  assign n7582 = n6928 ^ n6926;
  assign n7583 = n6953 ^ n6928;
  assign n7584 = n7583 ^ n6928;
  assign n7585 = n7582 & ~n7584;
  assign n7586 = n7585 ^ n6928;
  assign n7587 = n7581 & ~n7586;
  assign n7588 = n6897 & n7587;
  assign n7589 = n6985 & ~n6988;
  assign n7590 = ~n6994 & n7589;
  assign n7591 = ~n6990 & n7590;
  assign n7592 = ~n6969 & ~n6984;
  assign n7593 = ~n7589 & ~n7592;
  assign n7594 = n7197 & ~n7593;
  assign n7595 = ~n7004 & n7594;
  assign n7596 = ~n7591 & ~n7595;
  assign n7597 = ~n6993 & ~n7596;
  assign n7598 = ~n7218 & ~n7597;
  assign n7599 = ~n7588 & ~n7598;
  assign n7600 = n7579 & n7599;
  assign n7601 = n7203 & n7600;
  assign n7602 = n6975 & n7601;
  assign n7603 = n7211 & n7602;
  assign n7604 = n7603 ^ n5146;
  assign n7605 = n7604 ^ x310;
  assign n7606 = n7573 & ~n7605;
  assign n7607 = n7552 & n7606;
  assign n7608 = n7573 & n7605;
  assign n7609 = ~n7516 & ~n7550;
  assign n7610 = n7474 & n7609;
  assign n7611 = n7608 & n7610;
  assign n7612 = ~n7607 & ~n7611;
  assign n7613 = n7516 & ~n7550;
  assign n7614 = n7474 & n7613;
  assign n7615 = n7606 & n7614;
  assign n7616 = ~n7439 & n7473;
  assign n7617 = n7609 & n7616;
  assign n7618 = n7608 & n7617;
  assign n7619 = n7439 & ~n7473;
  assign n7620 = n7551 & n7619;
  assign n7621 = n7606 & n7620;
  assign n7622 = n7551 & n7616;
  assign n7623 = ~n7573 & ~n7605;
  assign n7624 = ~n7608 & ~n7623;
  assign n7625 = n7622 & ~n7624;
  assign n7626 = ~n7621 & ~n7625;
  assign n7627 = n7516 & n7550;
  assign n7628 = n7616 & n7627;
  assign n7629 = ~n7573 & n7605;
  assign n7630 = n7628 & n7629;
  assign n7631 = n7613 & n7616;
  assign n7632 = ~n7624 & n7631;
  assign n7633 = ~n7630 & ~n7632;
  assign n7634 = n7609 & n7619;
  assign n7635 = n7439 & n7473;
  assign n7636 = n7613 & n7635;
  assign n7637 = ~n7634 & ~n7636;
  assign n7638 = n7623 & ~n7637;
  assign n7639 = n7609 & n7635;
  assign n7640 = n7613 & n7619;
  assign n7641 = ~n7639 & ~n7640;
  assign n7642 = ~n7636 & n7641;
  assign n7643 = n7606 & ~n7642;
  assign n7644 = n7474 & n7627;
  assign n7645 = ~n7617 & ~n7644;
  assign n7646 = ~n7610 & n7645;
  assign n7647 = n7629 & ~n7646;
  assign n7648 = ~n7643 & ~n7647;
  assign n7649 = n7608 & n7644;
  assign n7650 = ~n7552 & ~n7614;
  assign n7651 = n7623 & ~n7650;
  assign n7660 = n7627 & n7635;
  assign n7661 = ~n7608 & ~n7620;
  assign n7654 = n7619 & n7627;
  assign n7662 = n7620 & n7623;
  assign n7663 = ~n7634 & ~n7662;
  assign n7664 = ~n7654 & n7663;
  assign n7665 = ~n7661 & ~n7664;
  assign n7666 = ~n7660 & ~n7665;
  assign n7652 = n7551 & n7635;
  assign n7653 = n7606 & n7628;
  assign n7655 = ~n7640 & ~n7654;
  assign n7656 = ~n7620 & n7655;
  assign n7657 = n7629 & ~n7656;
  assign n7658 = ~n7653 & ~n7657;
  assign n7659 = ~n7652 & n7658;
  assign n7667 = n7666 ^ n7659;
  assign n7668 = n7624 & n7667;
  assign n7669 = n7668 ^ n7666;
  assign n7670 = ~n7651 & n7669;
  assign n7671 = ~n7649 & n7670;
  assign n7672 = n7648 & n7671;
  assign n7673 = ~n7638 & n7672;
  assign n7674 = n7633 & n7673;
  assign n7675 = n7626 & n7674;
  assign n7676 = ~n7618 & n7675;
  assign n7677 = ~n7615 & n7676;
  assign n7678 = n7612 & n7677;
  assign n7679 = n7678 ^ n5306;
  assign n7680 = n7679 ^ x392;
  assign n7681 = ~n7408 & n7680;
  assign n7682 = n7132 & n7681;
  assign n7683 = n7515 ^ x316;
  assign n7684 = n6681 ^ x321;
  assign n7685 = ~n7683 & n7684;
  assign n7686 = n5375 ^ x320;
  assign n7687 = ~n6896 & n6976;
  assign n7688 = n6960 & ~n7218;
  assign n7689 = ~n7687 & ~n7688;
  assign n7690 = n6957 & n6971;
  assign n7691 = n6897 & ~n6991;
  assign n7692 = ~n7690 & ~n7691;
  assign n7693 = n7689 & n7692;
  assign n7694 = n6955 & n6990;
  assign n7695 = n6969 & n6972;
  assign n7696 = ~n7694 & ~n7695;
  assign n7697 = ~n6988 & ~n6993;
  assign n7698 = ~n6895 & ~n7697;
  assign n7699 = ~n6985 & n6990;
  assign n7700 = n6991 & n7006;
  assign n7701 = n6957 & ~n7700;
  assign n7702 = ~n7699 & ~n7701;
  assign n7703 = ~n6982 & ~n7001;
  assign n7704 = n6969 & ~n7703;
  assign n7705 = n6973 & n7697;
  assign n7706 = n6897 & ~n7705;
  assign n7707 = ~n7704 & ~n7706;
  assign n7708 = n7702 & n7707;
  assign n7709 = n7199 & n7708;
  assign n7710 = ~n7698 & n7709;
  assign n7711 = n7696 & n7710;
  assign n7712 = n7693 & n7711;
  assign n7713 = n7204 & n7712;
  assign n7714 = n7713 ^ n3926;
  assign n7715 = n7714 ^ x319;
  assign n7716 = n7686 & ~n7715;
  assign n7717 = n7133 & n7150;
  assign n7718 = n7134 & n7717;
  assign n7719 = ~n7151 & n7154;
  assign n7720 = ~n7718 & ~n7719;
  assign n7721 = n7133 & n7141;
  assign n7722 = n6785 & ~n7721;
  assign n7723 = ~n6836 & n6854;
  assign n7724 = n7156 & ~n7723;
  assign n7725 = n6840 & n7724;
  assign n7726 = ~n6844 & n7725;
  assign n7727 = n6852 & ~n7726;
  assign n7728 = ~n7722 & ~n7727;
  assign n7729 = n7720 & n7728;
  assign n7730 = n7729 ^ n3565;
  assign n7731 = n7730 ^ x318;
  assign n7732 = n7572 ^ x317;
  assign n7733 = ~n7731 & ~n7732;
  assign n7734 = n7716 & n7733;
  assign n7735 = n7685 & n7734;
  assign n7736 = n7683 & n7684;
  assign n7737 = ~n7686 & ~n7715;
  assign n7738 = n7731 & n7732;
  assign n7739 = n7737 & n7738;
  assign n7740 = ~n7731 & n7732;
  assign n7741 = n7716 & n7740;
  assign n7742 = ~n7739 & ~n7741;
  assign n7743 = n7736 & ~n7742;
  assign n7744 = ~n7686 & n7715;
  assign n7745 = n7731 & ~n7732;
  assign n7746 = n7744 & n7745;
  assign n7747 = n7716 & n7745;
  assign n7748 = ~n7746 & ~n7747;
  assign n7749 = n7685 & ~n7748;
  assign n7750 = ~n7743 & ~n7749;
  assign n7751 = n7684 ^ n7683;
  assign n7752 = n7733 & n7744;
  assign n7753 = n7751 & n7752;
  assign n7754 = n7686 & n7715;
  assign n7755 = n7745 & n7754;
  assign n7756 = ~n7684 & n7755;
  assign n7757 = ~n7753 & ~n7756;
  assign n7758 = n7738 & n7744;
  assign n7759 = n7733 & n7737;
  assign n7760 = ~n7758 & ~n7759;
  assign n7761 = n7736 & ~n7760;
  assign n7762 = ~n7683 & ~n7684;
  assign n7763 = n7737 & n7745;
  assign n7764 = ~n7734 & ~n7759;
  assign n7765 = ~n7763 & n7764;
  assign n7766 = n7762 & ~n7765;
  assign n7767 = n7741 & n7762;
  assign n7768 = n7740 & n7754;
  assign n7769 = n7685 & n7768;
  assign n7770 = n7683 & ~n7684;
  assign n7771 = n7768 & n7770;
  assign n7772 = n7733 & n7754;
  assign n7773 = ~n7734 & ~n7772;
  assign n7774 = n7770 & ~n7773;
  assign n7775 = n7738 & n7754;
  assign n7776 = n7740 & n7744;
  assign n7777 = ~n7775 & ~n7776;
  assign n7778 = ~n7739 & n7777;
  assign n7779 = n7762 & ~n7778;
  assign n7780 = ~n7774 & ~n7779;
  assign n7784 = n7716 & n7738;
  assign n7785 = n7737 & n7740;
  assign n7786 = ~n7784 & ~n7785;
  assign n7787 = ~n7758 & n7786;
  assign n7781 = ~n7763 & ~n7772;
  assign n7782 = ~n7755 & n7781;
  assign n7783 = ~n7752 & n7782;
  assign n7788 = n7787 ^ n7783;
  assign n7789 = n7788 ^ n7787;
  assign n7790 = n7787 ^ n7684;
  assign n7791 = n7790 ^ n7787;
  assign n7792 = ~n7789 & n7791;
  assign n7793 = n7792 ^ n7787;
  assign n7794 = ~n7751 & ~n7793;
  assign n7795 = n7794 ^ n7787;
  assign n7796 = n7780 & n7795;
  assign n7797 = ~n7771 & n7796;
  assign n7798 = ~n7769 & n7797;
  assign n7799 = ~n7767 & n7798;
  assign n7800 = ~n7766 & n7799;
  assign n7801 = ~n7761 & n7800;
  assign n7802 = n7757 & n7801;
  assign n7803 = n7750 & n7802;
  assign n7804 = ~n7735 & n7803;
  assign n7805 = n7804 ^ n3998;
  assign n7806 = n7805 ^ x388;
  assign n7807 = n6093 & n6116;
  assign n7808 = n6097 & n6115;
  assign n7809 = ~n7807 & ~n7808;
  assign n7810 = ~n6088 & n6111;
  assign n7811 = n6116 & ~n6120;
  assign n7812 = ~n7810 & ~n7811;
  assign n7813 = ~n6110 & ~n6115;
  assign n7814 = n6093 & ~n7813;
  assign n7815 = ~n5996 & ~n6096;
  assign n7816 = n7497 & n7815;
  assign n7817 = ~n6145 & n7816;
  assign n7818 = n6097 & ~n7817;
  assign n7819 = ~n7814 & ~n7818;
  assign n7820 = ~n5998 & n6142;
  assign n7821 = n7492 & n7820;
  assign n7822 = n6089 & ~n7821;
  assign n7823 = n7499 & n7815;
  assign n7824 = n6093 & ~n7823;
  assign n7825 = n6129 & ~n6141;
  assign n7826 = ~n6099 & n7825;
  assign n7827 = n6100 & ~n7826;
  assign n7828 = ~n7824 & ~n7827;
  assign n7829 = ~n7822 & n7828;
  assign n7830 = n7819 & n7829;
  assign n7831 = n7812 & n7830;
  assign n7832 = n7809 & n7831;
  assign n7833 = n7484 & n7832;
  assign n7834 = ~n6094 & n7833;
  assign n7835 = n7834 ^ n4049;
  assign n7836 = n7835 ^ x339;
  assign n7837 = n6893 ^ x334;
  assign n7838 = n7836 & ~n7837;
  assign n7839 = n5312 & n5315;
  assign n7840 = n5344 & ~n5360;
  assign n7841 = n5354 & n7840;
  assign n7842 = n5341 & ~n7841;
  assign n7843 = ~n7839 & ~n7842;
  assign n7844 = ~n7267 & n7527;
  assign n7845 = n4503 & ~n7844;
  assign n7846 = n5346 & ~n5353;
  assign n7847 = n5331 & ~n7846;
  assign n7848 = ~n7845 & ~n7847;
  assign n7849 = n7843 & n7848;
  assign n7850 = n5364 & n7532;
  assign n7851 = n5323 ^ n3999;
  assign n7852 = n7851 ^ n5323;
  assign n7853 = n5313 & ~n7526;
  assign n7854 = ~n5315 & n7853;
  assign n7855 = ~n5336 & ~n5353;
  assign n7856 = ~n5342 & n7855;
  assign n7857 = ~n5331 & n7856;
  assign n7858 = ~n7854 & ~n7857;
  assign n7859 = ~n5360 & ~n7858;
  assign n7860 = n7859 ^ n5323;
  assign n7861 = ~n7852 & ~n7860;
  assign n7862 = n7861 ^ n5323;
  assign n7863 = ~n7850 & ~n7862;
  assign n7864 = n7849 & n7863;
  assign n7865 = ~n5330 & n7864;
  assign n7866 = ~n7264 & n7865;
  assign n7867 = n5321 & n7866;
  assign n7868 = n7867 ^ n4339;
  assign n7869 = n7868 ^ x336;
  assign n7870 = n6780 ^ x335;
  assign n7871 = n7869 & n7870;
  assign n7872 = n6324 & n6349;
  assign n7873 = n6329 & n6362;
  assign n7874 = n6324 & ~n7246;
  assign n7875 = n6313 ^ n6235;
  assign n7876 = n7875 ^ n6313;
  assign n7877 = n7876 ^ n7875;
  assign n7878 = n7875 ^ n6265;
  assign n7879 = n7878 ^ n7875;
  assign n7880 = n7877 & ~n7879;
  assign n7881 = n7880 ^ n7875;
  assign n7882 = ~n6280 & n7881;
  assign n7883 = n7882 ^ n7875;
  assign n7884 = n6211 & n7883;
  assign n7885 = n6342 & n6376;
  assign n7886 = ~n6350 & n7885;
  assign n7887 = ~n6330 & ~n7886;
  assign n7888 = ~n7884 & ~n7887;
  assign n7889 = ~n7874 & n7888;
  assign n7890 = ~n7873 & n7889;
  assign n7891 = ~n7872 & n7890;
  assign n7892 = n7239 & n7891;
  assign n7893 = n6327 & n7892;
  assign n7894 = n7236 & n7893;
  assign n7895 = ~n7232 & n7894;
  assign n7896 = n7895 ^ n4305;
  assign n7897 = n7896 ^ x338;
  assign n7898 = n5681 & n5734;
  assign n7899 = n5720 & n7561;
  assign n7900 = ~n5723 & n7899;
  assign n7901 = n5686 & ~n7900;
  assign n7902 = ~n7898 & ~n7901;
  assign n7903 = ~n5694 & n5704;
  assign n7904 = ~n5710 & n5725;
  assign n7905 = n5511 & ~n7904;
  assign n7906 = ~n5510 & ~n5704;
  assign n7907 = ~n5708 & ~n5738;
  assign n7908 = ~n5717 & n7907;
  assign n7909 = ~n5510 & n7908;
  assign n7910 = ~n5723 & n7307;
  assign n7911 = ~n5717 & n7910;
  assign n7912 = ~n5704 & n5739;
  assign n7913 = ~n5681 & n7912;
  assign n7914 = ~n7911 & ~n7913;
  assign n7915 = ~n5728 & ~n7914;
  assign n7916 = ~n7909 & ~n7915;
  assign n7917 = ~n5699 & ~n7916;
  assign n7918 = ~n7906 & ~n7917;
  assign n7919 = ~n7905 & ~n7918;
  assign n7920 = ~n7903 & n7919;
  assign n7921 = n7902 & n7920;
  assign n7922 = n7294 & n7921;
  assign n7923 = n5685 & n7922;
  assign n7924 = n7923 ^ n4390;
  assign n7925 = n7924 ^ x337;
  assign n7926 = n7897 & ~n7925;
  assign n7927 = n7871 & n7926;
  assign n7928 = n7838 & n7927;
  assign n7929 = n7869 & ~n7870;
  assign n7930 = n7897 & n7925;
  assign n7931 = n7929 & n7930;
  assign n7932 = n7838 & n7931;
  assign n7933 = ~n7836 & n7837;
  assign n7934 = ~n7869 & ~n7870;
  assign n7935 = n7930 & n7934;
  assign n7936 = ~n7897 & ~n7925;
  assign n7937 = n7934 & n7936;
  assign n7938 = ~n7935 & ~n7937;
  assign n7939 = n7933 & ~n7938;
  assign n7940 = ~n7932 & ~n7939;
  assign n7941 = ~n7869 & n7870;
  assign n7942 = n7936 & n7941;
  assign n7943 = ~n7927 & ~n7942;
  assign n7944 = n7933 & ~n7943;
  assign n7945 = ~n7836 & ~n7837;
  assign n7946 = n7930 & n7941;
  assign n7947 = n7945 & n7946;
  assign n7948 = ~n7897 & n7925;
  assign n7949 = n7934 & n7948;
  assign n7950 = n7838 & n7949;
  assign n7951 = ~n7947 & ~n7950;
  assign n7952 = n7836 & n7837;
  assign n7953 = n7941 & n7948;
  assign n7954 = n7926 & n7941;
  assign n7955 = ~n7953 & ~n7954;
  assign n7956 = n7952 & ~n7955;
  assign n7957 = ~n7945 & ~n7952;
  assign n7958 = n7929 & n7936;
  assign n7959 = n7957 & n7958;
  assign n7960 = n7933 & n7953;
  assign n7961 = n7838 & ~n7955;
  assign n7962 = ~n7960 & ~n7961;
  assign n7963 = n7871 & n7936;
  assign n7964 = n7871 & n7948;
  assign n7965 = n7926 & n7934;
  assign n7966 = n7945 & n7965;
  assign n7967 = n7929 & n7948;
  assign n7968 = n7926 & n7929;
  assign n7969 = ~n7967 & ~n7968;
  assign n7970 = ~n7966 & n7969;
  assign n7971 = n7938 & n7970;
  assign n7972 = ~n7964 & n7971;
  assign n7973 = ~n7963 & n7972;
  assign n7974 = ~n7957 & ~n7973;
  assign n7975 = n7837 ^ n7836;
  assign n7976 = n7871 & n7930;
  assign n7977 = ~n7965 & ~n7976;
  assign n7978 = n7977 ^ n7837;
  assign n7979 = n7978 ^ n7977;
  assign n7980 = ~n7942 & ~n7946;
  assign n7981 = n7980 ^ n7977;
  assign n7982 = ~n7979 & n7981;
  assign n7983 = n7982 ^ n7977;
  assign n7984 = n7975 & ~n7983;
  assign n7985 = ~n7974 & ~n7984;
  assign n7986 = n7962 & n7985;
  assign n7987 = ~n7959 & n7986;
  assign n7988 = ~n7956 & n7987;
  assign n7989 = n7951 & n7988;
  assign n7990 = ~n7944 & n7989;
  assign n7991 = n7940 & n7990;
  assign n7992 = ~n7928 & n7991;
  assign n7993 = n7992 ^ n4501;
  assign n7994 = n7993 ^ x393;
  assign n7995 = ~n7806 & ~n7994;
  assign n7996 = n7682 & n7995;
  assign n7997 = ~n7806 & n7994;
  assign n7998 = n6745 & n7131;
  assign n7999 = n7681 & n7998;
  assign n8000 = ~n6745 & n7131;
  assign n8001 = ~n7408 & ~n7680;
  assign n8002 = n8000 & n8001;
  assign n8003 = ~n7999 & ~n8002;
  assign n8004 = n7997 & ~n8003;
  assign n8005 = ~n7996 & ~n8004;
  assign n8006 = ~n6745 & ~n7131;
  assign n8007 = n7681 & n8006;
  assign n8008 = n7997 & n8007;
  assign n8009 = n7408 & n7680;
  assign n8010 = n8000 & n8009;
  assign n8011 = n7408 & ~n7680;
  assign n8012 = n7998 & n8011;
  assign n8013 = ~n8010 & ~n8012;
  assign n8014 = n7995 & ~n8013;
  assign n8015 = ~n8008 & ~n8014;
  assign n8016 = n7806 & n7994;
  assign n8017 = n8000 & n8011;
  assign n8018 = n7681 & n8000;
  assign n8019 = ~n8012 & ~n8018;
  assign n8020 = ~n8017 & n8019;
  assign n8021 = n8016 & ~n8020;
  assign n8022 = n7682 & n8016;
  assign n8023 = n7132 & n8011;
  assign n8024 = n7997 & n8023;
  assign n8025 = ~n8022 & ~n8024;
  assign n8026 = n7998 & n8001;
  assign n8027 = n8006 & n8011;
  assign n8028 = ~n8026 & ~n8027;
  assign n8029 = n7806 & ~n7994;
  assign n8030 = ~n7997 & ~n8029;
  assign n8031 = ~n8028 & n8030;
  assign n8032 = n7132 & n8009;
  assign n8033 = n8001 & n8006;
  assign n8034 = ~n8032 & ~n8033;
  assign n8035 = n8016 & ~n8034;
  assign n8036 = ~n8031 & ~n8035;
  assign n8037 = n7131 ^ n6745;
  assign n8038 = n8037 ^ n7680;
  assign n8039 = n8038 ^ n7408;
  assign n8040 = n8039 ^ n7131;
  assign n8041 = n8040 ^ n7680;
  assign n8042 = n7680 ^ n7131;
  assign n8043 = n7408 ^ n7131;
  assign n8044 = n8043 ^ n7131;
  assign n8045 = n8042 & n8044;
  assign n8046 = n8045 ^ n7131;
  assign n8047 = n8041 & n8046;
  assign n8048 = n8047 ^ n8038;
  assign n8049 = n8029 & n8048;
  assign n8050 = ~n8007 & ~n8023;
  assign n8051 = ~n8018 & n8050;
  assign n8052 = n7995 & ~n8051;
  assign n8053 = n8006 & n8009;
  assign n8054 = ~n8027 & ~n8053;
  assign n8055 = ~n7682 & ~n8017;
  assign n8056 = n8054 & n8055;
  assign n8057 = n7997 & ~n8056;
  assign n8058 = ~n8052 & ~n8057;
  assign n8059 = ~n8049 & n8058;
  assign n8060 = n8036 & n8059;
  assign n8061 = n8025 & n8060;
  assign n8062 = ~n8021 & n8061;
  assign n8063 = n8015 & n8062;
  assign n8064 = n8005 & n8063;
  assign n8065 = n8064 ^ n5375;
  assign n8066 = n8065 ^ x418;
  assign n8067 = n7229 ^ x345;
  assign n8068 = n7896 ^ x340;
  assign n8069 = n8067 & n8068;
  assign n8070 = n7835 ^ x341;
  assign n8071 = ~n6850 & n7134;
  assign n8072 = ~n6873 & n7154;
  assign n8073 = ~n8071 & ~n8072;
  assign n8074 = n6784 & ~n6890;
  assign n8075 = n8073 & ~n8074;
  assign n8076 = n8075 ^ n5443;
  assign n8077 = n8076 ^ x342;
  assign n8078 = n8070 & ~n8077;
  assign n8079 = ~n6396 & n6490;
  assign n8080 = n6480 & ~n6750;
  assign n8081 = ~n8079 & ~n8080;
  assign n8082 = n6464 & ~n6502;
  assign n8083 = n6762 & n6768;
  assign n8084 = ~n6523 & n8083;
  assign n8085 = n6469 & ~n8084;
  assign n8086 = ~n8082 & ~n8085;
  assign n8087 = n6524 & n6757;
  assign n8088 = n6396 & ~n8087;
  assign n8091 = ~n6472 & n6483;
  assign n8092 = ~n6503 & n8091;
  assign n8089 = n6475 & ~n6492;
  assign n8090 = ~n6478 & n8089;
  assign n8093 = n8092 ^ n8090;
  assign n8094 = n8092 ^ n6394;
  assign n8095 = n8094 ^ n8092;
  assign n8096 = n8093 & n8095;
  assign n8097 = n8096 ^ n8092;
  assign n8098 = n6395 & ~n8097;
  assign n8099 = ~n8088 & ~n8098;
  assign n8100 = n8086 & n8099;
  assign n8101 = n8081 & n8100;
  assign n8102 = n6752 & n8101;
  assign n8103 = n6748 & n8102;
  assign n8104 = n8103 ^ n5429;
  assign n8105 = n8104 ^ x343;
  assign n8106 = n7193 ^ x344;
  assign n8107 = ~n8105 & n8106;
  assign n8108 = n8078 & n8107;
  assign n8109 = n8069 & n8108;
  assign n8110 = n8105 & ~n8106;
  assign n8111 = n8078 & n8110;
  assign n8112 = n8069 & n8111;
  assign n8115 = ~n8067 & n8068;
  assign n8113 = n8105 & n8106;
  assign n8114 = n8078 & n8113;
  assign n8116 = n8115 ^ n8114;
  assign n8117 = n8067 & ~n8068;
  assign n8118 = n8117 ^ n8114;
  assign n8119 = n8118 ^ n8117;
  assign n8120 = n8070 & n8077;
  assign n8121 = n8110 & n8120;
  assign n8122 = n8121 ^ n8117;
  assign n8123 = ~n8119 & ~n8122;
  assign n8124 = n8123 ^ n8117;
  assign n8125 = n8116 & n8124;
  assign n8126 = n8125 ^ n8115;
  assign n8127 = ~n8112 & ~n8126;
  assign n8128 = ~n8070 & ~n8077;
  assign n8129 = n8113 & n8128;
  assign n8130 = ~n8105 & ~n8106;
  assign n8131 = n8128 & n8130;
  assign n8132 = ~n8129 & ~n8131;
  assign n8133 = n8069 & ~n8132;
  assign n8134 = ~n8070 & n8077;
  assign n8135 = n8113 & n8134;
  assign n8136 = ~n8131 & ~n8135;
  assign n8137 = n8117 & ~n8136;
  assign n8138 = ~n8133 & ~n8137;
  assign n8139 = n8078 & n8130;
  assign n8140 = n8107 & n8134;
  assign n8141 = n8110 & n8128;
  assign n8142 = ~n8140 & ~n8141;
  assign n8143 = ~n8139 & n8142;
  assign n8144 = n8143 ^ n8115;
  assign n8145 = n8143 ^ n8117;
  assign n8146 = n8145 ^ n8117;
  assign n8147 = n8117 ^ n8108;
  assign n8148 = n8146 & ~n8147;
  assign n8149 = n8148 ^ n8117;
  assign n8150 = ~n8144 & n8149;
  assign n8151 = n8150 ^ n8115;
  assign n8152 = n8138 & ~n8151;
  assign n8153 = n8107 & n8128;
  assign n8154 = n8130 & n8134;
  assign n8155 = ~n8153 & ~n8154;
  assign n8156 = n8068 & ~n8155;
  assign n8157 = n8107 & n8120;
  assign n8158 = ~n8121 & ~n8157;
  assign n8159 = n8067 & ~n8158;
  assign n8160 = ~n8156 & ~n8159;
  assign n8161 = ~n8067 & ~n8068;
  assign n8162 = ~n8108 & ~n8157;
  assign n8163 = ~n8121 & n8136;
  assign n8164 = n8162 & n8163;
  assign n8165 = n8142 & n8164;
  assign n8166 = ~n8129 & n8165;
  assign n8167 = n8161 & n8166;
  assign n8168 = n8160 & ~n8167;
  assign n8169 = n8152 & n8168;
  assign n8170 = n8127 & n8169;
  assign n8171 = ~n8109 & n8170;
  assign n8172 = n8171 ^ n5509;
  assign n8173 = n8172 ^ x352;
  assign n8174 = n7331 & n7333;
  assign n8175 = n7343 & n7374;
  assign n8176 = ~n8174 & ~n8175;
  assign n8177 = n7195 & n7375;
  assign n8178 = n7354 & n7391;
  assign n8179 = ~n8177 & ~n8178;
  assign n8180 = ~n7376 & n7379;
  assign n8181 = n7333 & ~n8180;
  assign n8182 = ~n7352 & ~n7391;
  assign n8183 = n7377 & n8182;
  assign n8184 = ~n7348 & n8183;
  assign n8185 = ~n7336 & n8184;
  assign n8186 = n7343 & ~n8185;
  assign n8187 = ~n8181 & ~n8186;
  assign n8188 = ~n7164 & n7378;
  assign n8189 = n7195 & ~n7358;
  assign n8190 = ~n7384 & ~n7390;
  assign n8191 = ~n8189 & ~n8190;
  assign n8192 = n7354 ^ n7336;
  assign n8193 = ~n7336 & ~n8192;
  assign n8194 = n8193 ^ n7336;
  assign n8195 = ~n7356 & ~n7375;
  assign n8196 = n8195 ^ n7336;
  assign n8197 = ~n8194 & ~n8196;
  assign n8198 = n8197 ^ n8193;
  assign n8199 = n8198 ^ n7336;
  assign n8200 = n8199 ^ n7354;
  assign n8201 = n8191 & ~n8200;
  assign n8202 = n8201 ^ n8191;
  assign n8203 = ~n8188 & n8202;
  assign n8204 = n8187 & n8203;
  assign n8205 = n8179 & n8204;
  assign n8206 = n7371 & n8205;
  assign n8207 = n8176 & n8206;
  assign n8208 = n7342 & n8207;
  assign n8209 = n8208 ^ n5408;
  assign n8210 = n8209 ^ x357;
  assign n8211 = n8173 & n8210;
  assign n8212 = n7606 & n7631;
  assign n8213 = n7605 ^ n7573;
  assign n8214 = n7610 ^ n7605;
  assign n8215 = n8214 ^ n7610;
  assign n8216 = ~n7614 & ~n7654;
  assign n8217 = n8216 ^ n7610;
  assign n8218 = n8215 & ~n8217;
  assign n8219 = n8218 ^ n7610;
  assign n8220 = ~n8213 & n8219;
  assign n8221 = ~n8212 & ~n8220;
  assign n8222 = n7623 & n7654;
  assign n8223 = ~n7662 & ~n8222;
  assign n8224 = n7606 & n7660;
  assign n8225 = ~n7636 & ~n7652;
  assign n8226 = n7629 & ~n8225;
  assign n8227 = ~n8224 & ~n8226;
  assign n8228 = n7606 & ~n8225;
  assign n8229 = ~n7552 & ~n7610;
  assign n8230 = ~n7628 & n8229;
  assign n8231 = n7629 & ~n8230;
  assign n8232 = ~n8228 & ~n8231;
  assign n8233 = n7629 & n7660;
  assign n8234 = n7608 & n7620;
  assign n8235 = n7606 & n7634;
  assign n8236 = ~n8234 & ~n8235;
  assign n8237 = ~n8233 & n8236;
  assign n8238 = n7606 & n7622;
  assign n8239 = n7629 & ~n8216;
  assign n8240 = ~n8238 & ~n8239;
  assign n8241 = ~n7634 & ~n7639;
  assign n8242 = ~n7628 & n8241;
  assign n8243 = n7608 & ~n8242;
  assign n8244 = n7641 & ~n7660;
  assign n8245 = ~n7631 & n8244;
  assign n8246 = n7623 & ~n8245;
  assign n8247 = ~n8243 & ~n8246;
  assign n8248 = n8240 & n8247;
  assign n8249 = n8237 & n8248;
  assign n8250 = n7626 & n8249;
  assign n8251 = n8232 & n8250;
  assign n8252 = n8227 & n8251;
  assign n8253 = n8223 & n8252;
  assign n8254 = ~n7618 & n8253;
  assign n8255 = ~n7615 & n8254;
  assign n8256 = n8221 & n8255;
  assign n8257 = n8256 ^ n5676;
  assign n8258 = n8257 ^ x354;
  assign n8259 = n7067 & n7102;
  assign n8260 = n6782 & n7077;
  assign n8261 = ~n8259 & ~n8260;
  assign n8262 = n6782 & ~n7098;
  assign n8263 = ~n6782 & ~n7072;
  assign n8264 = ~n7085 & ~n7104;
  assign n8265 = ~n8263 & ~n8264;
  assign n8266 = n7067 & n7091;
  assign n8267 = n7065 & n7080;
  assign n8268 = ~n8266 & ~n8267;
  assign n8269 = ~n7081 & ~n7089;
  assign n8270 = ~n7105 & n8269;
  assign n8271 = ~n7065 & n8270;
  assign n8272 = n7072 & ~n8271;
  assign n8273 = n7080 ^ n7067;
  assign n8280 = ~n7106 & n7115;
  assign n8274 = n7063 ^ n6894;
  assign n8275 = n7030 ^ n7028;
  assign n8276 = n7063 ^ n7030;
  assign n8277 = n8275 & ~n8276;
  assign n8278 = n8274 & n8277;
  assign n8279 = n8278 ^ n8274;
  assign n8281 = n8280 ^ n8279;
  assign n8282 = n8280 ^ n7080;
  assign n8283 = n8282 ^ n8280;
  assign n8284 = n8281 & n8283;
  assign n8285 = n8284 ^ n8280;
  assign n8286 = n8273 & n8285;
  assign n8287 = n8286 ^ n7067;
  assign n8288 = ~n8272 & ~n8287;
  assign n8289 = n8268 & n8288;
  assign n8290 = ~n8265 & n8289;
  assign n8291 = ~n8262 & n8290;
  assign n8292 = n7116 ^ n7102;
  assign n8293 = n8292 ^ n7102;
  assign n8294 = n7102 ^ n6746;
  assign n8295 = n8294 ^ n7102;
  assign n8296 = ~n8293 & ~n8295;
  assign n8297 = n8296 ^ n7102;
  assign n8298 = n6781 & n8297;
  assign n8299 = n8298 ^ n7102;
  assign n8300 = n8291 & ~n8299;
  assign n8301 = n7094 & n8300;
  assign n8302 = n8261 & n8301;
  assign n8303 = ~n7079 & n8302;
  assign n8304 = n8303 ^ n5556;
  assign n8305 = n8304 ^ x355;
  assign n8306 = ~n8258 & ~n8305;
  assign n8307 = n6682 & n6696;
  assign n8308 = n6393 & n8307;
  assign n8309 = n6538 & n6736;
  assign n8310 = ~n8308 & ~n8309;
  assign n8311 = ~n6393 & n6736;
  assign n8312 = ~n6694 & ~n8311;
  assign n8313 = ~n6707 & n8312;
  assign n8314 = n6702 & ~n8313;
  assign n8315 = n6538 & ~n6682;
  assign n8316 = n6683 & ~n6736;
  assign n8317 = ~n8315 & ~n8316;
  assign n8318 = n6709 & n8317;
  assign n8319 = n6730 & ~n8318;
  assign n8320 = ~n8314 & ~n8319;
  assign n8321 = n6704 ^ n6693;
  assign n8322 = ~n6682 & n8321;
  assign n8323 = n8322 ^ n6704;
  assign n8324 = n6712 & ~n8323;
  assign n8325 = n8310 & n8324;
  assign n8326 = n8325 ^ n5376;
  assign n8327 = n8326 ^ n8325;
  assign n8328 = n6699 & n6709;
  assign n8329 = ~n6734 & n8328;
  assign n8330 = n8329 ^ n8325;
  assign n8331 = ~n8327 & n8330;
  assign n8332 = n8331 ^ n8325;
  assign n8333 = n5753 & ~n8332;
  assign n8334 = n8320 & ~n8333;
  assign n8335 = n8310 & n8334;
  assign n8336 = n8335 ^ n5621;
  assign n8337 = n8336 ^ x353;
  assign n8338 = n7931 & n7933;
  assign n8339 = n7945 & n7968;
  assign n8340 = ~n8338 & ~n8339;
  assign n8341 = n7945 & n7949;
  assign n8342 = ~n7946 & ~n7964;
  assign n8343 = n7933 & ~n8342;
  assign n8344 = ~n8341 & ~n8343;
  assign n8345 = ~n7957 & n7965;
  assign n8346 = n7938 & ~n7953;
  assign n8347 = ~n7967 & n8346;
  assign n8348 = ~n7942 & n8347;
  assign n8349 = n7838 & ~n8348;
  assign n8350 = ~n8345 & ~n8349;
  assign n8351 = n8344 & n8350;
  assign n8352 = n7942 & n7952;
  assign n8353 = n7955 & ~n8352;
  assign n8354 = ~n7942 & ~n7954;
  assign n8355 = ~n7945 & n8354;
  assign n8356 = ~n8353 & ~n8355;
  assign n8357 = ~n7976 & ~n8356;
  assign n8358 = ~n7964 & n8357;
  assign n8359 = ~n7957 & ~n8358;
  assign n8360 = n7963 ^ n7952;
  assign n8361 = n8360 ^ n7963;
  assign n8362 = ~n7958 & n7969;
  assign n8363 = n8362 ^ n7963;
  assign n8364 = n8361 & ~n8363;
  assign n8365 = n8364 ^ n7963;
  assign n8366 = ~n8359 & ~n8365;
  assign n8367 = n8351 & n8366;
  assign n8368 = ~n7944 & n8367;
  assign n8369 = n8340 & n8368;
  assign n8370 = ~n7928 & n8369;
  assign n8371 = n7940 & n8370;
  assign n8372 = n8371 ^ n5592;
  assign n8373 = n8372 ^ x356;
  assign n8374 = n8337 & ~n8373;
  assign n8375 = n8306 & n8374;
  assign n8376 = n8211 & n8375;
  assign n8377 = ~n8258 & n8305;
  assign n8378 = n8337 & n8373;
  assign n8379 = n8377 & n8378;
  assign n8380 = n8211 & n8379;
  assign n8381 = ~n8173 & ~n8210;
  assign n8382 = n8374 & n8377;
  assign n8383 = n8381 & n8382;
  assign n8384 = ~n8380 & ~n8383;
  assign n8385 = n8173 & ~n8210;
  assign n8386 = n8258 & n8305;
  assign n8387 = n8374 & n8386;
  assign n8388 = n8385 & n8387;
  assign n8389 = ~n8173 & n8210;
  assign n8390 = n8306 & n8378;
  assign n8391 = n8258 & ~n8305;
  assign n8392 = n8374 & n8391;
  assign n8393 = ~n8390 & ~n8392;
  assign n8394 = n8389 & ~n8393;
  assign n8395 = ~n8388 & ~n8394;
  assign n8396 = n8384 & n8395;
  assign n8397 = ~n8337 & n8373;
  assign n8398 = n8391 & n8397;
  assign n8399 = n8389 & n8398;
  assign n8400 = n8378 & n8386;
  assign n8401 = n8381 & n8400;
  assign n8402 = ~n8399 & ~n8401;
  assign n8403 = n8386 & n8397;
  assign n8404 = ~n8337 & ~n8373;
  assign n8405 = n8306 & n8404;
  assign n8406 = ~n8403 & ~n8405;
  assign n8407 = n8211 & ~n8406;
  assign n8408 = n8378 & n8391;
  assign n8409 = ~n8375 & ~n8408;
  assign n8410 = n8385 & ~n8409;
  assign n8411 = ~n8407 & ~n8410;
  assign n8412 = n8402 & n8411;
  assign n8413 = n8211 & n8400;
  assign n8414 = n8385 & n8400;
  assign n8415 = n8306 & n8397;
  assign n8416 = ~n8387 & ~n8415;
  assign n8417 = n8211 & ~n8416;
  assign n8418 = ~n8414 & ~n8417;
  assign n8419 = ~n8379 & ~n8392;
  assign n8420 = n8381 & ~n8419;
  assign n8421 = n8391 & n8404;
  assign n8422 = n8386 & n8404;
  assign n8423 = ~n8421 & ~n8422;
  assign n8424 = ~n8385 & n8423;
  assign n8425 = n8377 & n8397;
  assign n8426 = ~n8421 & ~n8425;
  assign n8427 = ~n8381 & n8426;
  assign n8428 = ~n8415 & n8427;
  assign n8429 = ~n8424 & ~n8428;
  assign n8430 = ~n8398 & ~n8429;
  assign n8431 = n8430 ^ n8173;
  assign n8432 = n8431 ^ n8430;
  assign n8433 = n8377 & n8404;
  assign n8434 = ~n8403 & ~n8433;
  assign n8435 = ~n8408 & n8434;
  assign n8436 = ~n8387 & n8435;
  assign n8437 = ~n8382 & n8436;
  assign n8438 = n8437 ^ n8430;
  assign n8439 = n8438 ^ n8430;
  assign n8440 = ~n8432 & ~n8439;
  assign n8441 = n8440 ^ n8430;
  assign n8442 = n8210 & ~n8441;
  assign n8443 = n8442 ^ n8430;
  assign n8444 = ~n8420 & n8443;
  assign n8445 = n8418 & n8444;
  assign n8446 = ~n8413 & n8445;
  assign n8447 = n8412 & n8446;
  assign n8448 = n8396 & n8447;
  assign n8449 = ~n8376 & n8448;
  assign n8450 = n8210 ^ n8173;
  assign n8451 = n8415 ^ n8210;
  assign n8452 = n8451 ^ n8415;
  assign n8453 = n8421 ^ n8415;
  assign n8454 = n8452 & n8453;
  assign n8455 = n8454 ^ n8415;
  assign n8456 = ~n8450 & n8455;
  assign n8457 = n8449 & ~n8456;
  assign n8458 = n8457 ^ n5752;
  assign n8459 = n8458 ^ x423;
  assign n8460 = ~n8066 & ~n8459;
  assign n8461 = n8209 ^ x359;
  assign n8462 = n7762 & ~n7777;
  assign n8463 = n7736 & ~n7748;
  assign n8464 = ~n8462 & ~n8463;
  assign n8465 = n7685 & n7775;
  assign n8466 = ~n7769 & ~n8465;
  assign n8467 = n7736 & n7755;
  assign n8468 = n7770 & n7775;
  assign n8469 = ~n8467 & ~n8468;
  assign n8470 = ~n7776 & ~n7784;
  assign n8471 = n7751 & ~n8470;
  assign n8472 = ~n7746 & n7781;
  assign n8473 = n7685 & ~n8472;
  assign n8474 = n7736 & n7785;
  assign n8475 = ~n7764 & n7770;
  assign n8476 = ~n8474 & ~n8475;
  assign n8477 = ~n7684 & n7758;
  assign n8478 = n7770 & ~n7781;
  assign n8479 = ~n8477 & ~n8478;
  assign n8480 = ~n7752 & ~n7768;
  assign n8481 = n7736 & ~n8480;
  assign n8482 = ~n7759 & ~n7772;
  assign n8483 = n7748 & n8482;
  assign n8484 = n7762 & ~n8483;
  assign n8485 = ~n8481 & ~n8484;
  assign n8486 = n8479 & n8485;
  assign n8487 = n8476 & n8486;
  assign n8488 = ~n8473 & n8487;
  assign n8489 = ~n8471 & n8488;
  assign n8490 = n8469 & n8489;
  assign n8491 = ~n7743 & n8490;
  assign n8492 = n8466 & n8491;
  assign n8493 = n8464 & n8492;
  assign n8494 = ~n7767 & n8493;
  assign n8495 = ~n7735 & n8494;
  assign n8496 = n8495 ^ n6563;
  assign n8497 = n8496 ^ x360;
  assign n8498 = n8461 & n8497;
  assign n8499 = ~n8115 & ~n8117;
  assign n8500 = n8120 & n8130;
  assign n8501 = n8499 & n8500;
  assign n8502 = ~n8114 & ~n8121;
  assign n8503 = n8161 & ~n8502;
  assign n8504 = ~n8501 & ~n8503;
  assign n8505 = ~n8112 & n8504;
  assign n8506 = n8140 & n8161;
  assign n8507 = n8113 & n8120;
  assign n8508 = n8069 & n8507;
  assign n8509 = ~n8506 & ~n8508;
  assign n8510 = n8161 & n8507;
  assign n8511 = n8111 & n8115;
  assign n8512 = n8117 & n8121;
  assign n8513 = ~n8511 & ~n8512;
  assign n8514 = ~n8132 & n8499;
  assign n8515 = n8110 & n8134;
  assign n8516 = ~n8140 & ~n8515;
  assign n8517 = ~n8157 & n8516;
  assign n8518 = n8069 & ~n8517;
  assign n8519 = ~n8514 & ~n8518;
  assign n8520 = n8513 & n8519;
  assign n8521 = n8139 & n8161;
  assign n8522 = ~n8153 & ~n8515;
  assign n8523 = ~n8141 & n8522;
  assign n8524 = n8162 & n8523;
  assign n8525 = ~n8135 & n8524;
  assign n8526 = ~n8154 & n8525;
  assign n8527 = ~n8499 & ~n8526;
  assign n8528 = ~n8521 & ~n8527;
  assign n8529 = n8520 & n8528;
  assign n8530 = ~n8510 & n8529;
  assign n8531 = n8509 & n8530;
  assign n8532 = n8505 & n8531;
  assign n8533 = n8532 ^ n6599;
  assign n8534 = n8533 ^ x361;
  assign n8535 = n6782 & n7091;
  assign n8536 = ~n7096 & ~n7106;
  assign n8537 = n7072 & ~n8536;
  assign n8538 = ~n8535 & ~n8537;
  assign n8539 = ~n7104 & n7115;
  assign n8540 = n6782 & ~n8539;
  assign n8541 = n7103 & n8264;
  assign n8542 = n7080 & ~n8541;
  assign n8543 = ~n8540 & ~n8542;
  assign n8544 = n7072 & ~n7121;
  assign n8545 = n7108 & n8269;
  assign n8546 = ~n7087 & n8545;
  assign n8547 = n7067 & ~n8546;
  assign n8548 = ~n8544 & ~n8547;
  assign n8549 = n8543 & n8548;
  assign n8550 = n8261 & n8549;
  assign n8551 = n7095 & n8550;
  assign n8552 = n8538 & n8551;
  assign n8553 = ~n7083 & n8552;
  assign n8554 = n7071 & n8553;
  assign n8555 = n8554 ^ n6209;
  assign n8556 = n8555 ^ x362;
  assign n8557 = ~n8534 & n8556;
  assign n8558 = n8498 & n8557;
  assign n8559 = n8461 & ~n8497;
  assign n8560 = n8534 & ~n8556;
  assign n8561 = n8559 & n8560;
  assign n8562 = ~n8558 & ~n8561;
  assign n8563 = n7163 ^ x305;
  assign n8564 = n6097 & n6121;
  assign n8565 = n7499 & n7820;
  assign n8566 = n6093 & ~n8565;
  assign n8567 = ~n8564 & ~n8566;
  assign n8568 = n6100 & ~n6131;
  assign n8569 = n6134 & n6142;
  assign n8570 = n6089 & ~n8569;
  assign n8571 = ~n6111 & ~n6145;
  assign n8572 = ~n6120 & ~n8571;
  assign n8573 = ~n8570 & ~n8572;
  assign n8574 = ~n8568 & n8573;
  assign n8575 = n8567 & n8574;
  assign n8576 = n7809 & n8575;
  assign n8577 = n7489 & n8576;
  assign n8578 = n6104 & n8577;
  assign n8579 = n7476 & n8578;
  assign n8580 = ~n7502 & n8579;
  assign n8581 = ~n6090 & n8580;
  assign n8582 = n8581 ^ n5880;
  assign n8583 = n8582 ^ x307;
  assign n8584 = n8563 & ~n8583;
  assign n8585 = n6643 & n6665;
  assign n8586 = ~n6651 & n6667;
  assign n8587 = n6542 & ~n8586;
  assign n8588 = ~n8585 & ~n8587;
  assign n8589 = n6631 & ~n6664;
  assign n8590 = ~n7166 & ~n7172;
  assign n8591 = n6626 & n6659;
  assign n8592 = ~n6618 & ~n6660;
  assign n8593 = n6542 & ~n8592;
  assign n8594 = ~n8591 & ~n8593;
  assign n8595 = n6641 & n6643;
  assign n8596 = ~n6651 & n7168;
  assign n8597 = ~n6631 & n8596;
  assign n8598 = ~n6626 & ~n6646;
  assign n8599 = n8586 & n8598;
  assign n8600 = ~n8597 & ~n8599;
  assign n8601 = ~n7172 & n8600;
  assign n8602 = ~n8595 & ~n8601;
  assign n8603 = n8594 & n8602;
  assign n8604 = n6650 & n8603;
  assign n8605 = n6645 & n8604;
  assign n8606 = ~n8590 & n8605;
  assign n8607 = ~n8589 & n8606;
  assign n8608 = n8588 & n8607;
  assign n8609 = ~n7057 & n8608;
  assign n8610 = n8609 ^ n5917;
  assign n8611 = n8610 ^ x306;
  assign n8612 = n7604 ^ x308;
  assign n8613 = n8611 & ~n8612;
  assign n8614 = n8584 & n8613;
  assign n8615 = n7291 ^ x304;
  assign n8616 = n7438 ^ x309;
  assign n8617 = ~n8615 & n8616;
  assign n8618 = n8563 & n8583;
  assign n8619 = n8611 & n8612;
  assign n8620 = n8618 & n8619;
  assign n8621 = n8617 & n8620;
  assign n8622 = ~n8615 & ~n8616;
  assign n8623 = ~n8563 & ~n8583;
  assign n8624 = ~n8611 & n8612;
  assign n8625 = n8623 & n8624;
  assign n8626 = n8622 & n8625;
  assign n8627 = n8615 & ~n8616;
  assign n8628 = ~n8563 & n8583;
  assign n8629 = n8624 & n8628;
  assign n8630 = n8627 & n8629;
  assign n8631 = ~n8626 & ~n8630;
  assign n8632 = ~n8621 & n8631;
  assign n8633 = n8615 & n8616;
  assign n8634 = ~n8611 & ~n8612;
  assign n8635 = n8618 & n8634;
  assign n8636 = n8633 & n8635;
  assign n8637 = n8584 & n8634;
  assign n8638 = n8633 & n8637;
  assign n8639 = n8620 & n8633;
  assign n8640 = n8619 & n8623;
  assign n8641 = n8617 & n8640;
  assign n8642 = ~n8639 & ~n8641;
  assign n8643 = n8618 & n8624;
  assign n8644 = n8617 & n8643;
  assign n8645 = ~n8622 & ~n8633;
  assign n8646 = n8613 & n8628;
  assign n8647 = ~n8645 & n8646;
  assign n8648 = ~n8644 & ~n8647;
  assign n8649 = n8613 & n8623;
  assign n8650 = ~n8640 & ~n8649;
  assign n8651 = ~n8625 & n8650;
  assign n8652 = n8633 & ~n8651;
  assign n8653 = n8612 ^ n8583;
  assign n8654 = n8583 ^ n8563;
  assign n8655 = n8654 ^ n8612;
  assign n8656 = n8655 ^ n8583;
  assign n8657 = ~n8653 & ~n8656;
  assign n8658 = n8657 ^ n8583;
  assign n8659 = ~n8611 & n8658;
  assign n8660 = n8659 ^ n8655;
  assign n8661 = n8627 & ~n8660;
  assign n8662 = n8619 & n8628;
  assign n8663 = n8628 & n8634;
  assign n8664 = ~n8662 & ~n8663;
  assign n8665 = n8623 & n8634;
  assign n8666 = ~n8625 & ~n8665;
  assign n8667 = n8664 & n8666;
  assign n8668 = n8617 & ~n8667;
  assign n8669 = n8584 & n8619;
  assign n8670 = n8613 & n8618;
  assign n8671 = ~n8669 & ~n8670;
  assign n8672 = ~n8637 & n8671;
  assign n8673 = ~n8629 & n8672;
  assign n8674 = ~n8635 & n8673;
  assign n8675 = n8622 & ~n8674;
  assign n8676 = ~n8668 & ~n8675;
  assign n8677 = ~n8661 & n8676;
  assign n8678 = ~n8652 & n8677;
  assign n8679 = n8648 & n8678;
  assign n8680 = n8642 & n8679;
  assign n8681 = ~n8638 & n8680;
  assign n8682 = ~n8636 & n8681;
  assign n8683 = n8632 & n8682;
  assign n8684 = ~n8614 & n8683;
  assign n8685 = n8684 ^ n6264;
  assign n8686 = n8685 ^ x363;
  assign n8687 = n8372 ^ x358;
  assign n8688 = ~n8686 & ~n8687;
  assign n8689 = ~n8562 & n8688;
  assign n8690 = ~n8461 & n8497;
  assign n8691 = n8557 & n8690;
  assign n8692 = ~n8461 & ~n8497;
  assign n8693 = n8560 & n8692;
  assign n8694 = ~n8691 & ~n8693;
  assign n8695 = n8686 & ~n8687;
  assign n8696 = ~n8694 & n8695;
  assign n8697 = ~n8534 & ~n8556;
  assign n8698 = n8692 & n8697;
  assign n8699 = ~n8686 & n8687;
  assign n8700 = n8698 & n8699;
  assign n8701 = n8498 & n8560;
  assign n8702 = n8695 & n8701;
  assign n8703 = n8534 & n8556;
  assign n8704 = n8690 & n8703;
  assign n8705 = n8699 & n8704;
  assign n8706 = n8559 & n8703;
  assign n8707 = n8686 & n8687;
  assign n8708 = n8706 & n8707;
  assign n8709 = ~n8705 & ~n8708;
  assign n8710 = ~n8702 & n8709;
  assign n8711 = ~n8700 & n8710;
  assign n8712 = n8558 & n8686;
  assign n8713 = n8561 & n8687;
  assign n8714 = ~n8712 & ~n8713;
  assign n8715 = n8692 & n8703;
  assign n8716 = ~n8556 & n8690;
  assign n8717 = ~n8534 & n8716;
  assign n8718 = ~n8715 & ~n8717;
  assign n8719 = n8707 & ~n8718;
  assign n8720 = n8534 & n8716;
  assign n8721 = n8557 & n8559;
  assign n8722 = ~n8715 & ~n8721;
  assign n8723 = ~n8720 & n8722;
  assign n8724 = n8688 & ~n8723;
  assign n8725 = ~n8719 & ~n8724;
  assign n8726 = n8557 & n8692;
  assign n8727 = ~n8698 & ~n8726;
  assign n8728 = ~n8701 & n8727;
  assign n8729 = n8687 ^ n8686;
  assign n8730 = ~n8728 & ~n8729;
  assign n8731 = n8559 & n8697;
  assign n8732 = ~n8706 & ~n8731;
  assign n8733 = ~n8704 & ~n8717;
  assign n8734 = n8732 & n8733;
  assign n8735 = n8695 & ~n8734;
  assign n8736 = n8498 & n8703;
  assign n8737 = ~n8691 & ~n8736;
  assign n8738 = n8498 & n8697;
  assign n8739 = ~n8721 & ~n8738;
  assign n8740 = n8737 & n8739;
  assign n8741 = ~n8693 & n8740;
  assign n8742 = n8699 & ~n8741;
  assign n8743 = ~n8735 & ~n8742;
  assign n8744 = ~n8730 & n8743;
  assign n8745 = n8725 & n8744;
  assign n8746 = n8714 & n8745;
  assign n8747 = n8711 & n8746;
  assign n8748 = ~n8696 & n8747;
  assign n8749 = ~n8689 & n8748;
  assign n8750 = n8749 ^ n6681;
  assign n8751 = n8750 ^ x419;
  assign n8752 = ~n7617 & ~n7628;
  assign n8753 = n7606 & ~n8752;
  assign n8754 = ~n7622 & ~n7640;
  assign n8755 = n7623 & ~n8754;
  assign n8756 = ~n8753 & ~n8755;
  assign n8757 = ~n7620 & ~n7631;
  assign n8758 = n7629 & ~n8757;
  assign n8759 = ~n7618 & n8225;
  assign n8760 = ~n7614 & n8759;
  assign n8761 = ~n7644 & n8760;
  assign n8762 = ~n7624 & ~n8761;
  assign n8763 = ~n8758 & ~n8762;
  assign n8764 = n8756 & n8763;
  assign n8765 = n8237 & n8764;
  assign n8766 = n7654 ^ n7605;
  assign n8767 = n8766 ^ n7654;
  assign n8768 = n7654 ^ n7641;
  assign n8769 = n8767 & ~n8768;
  assign n8770 = n8769 ^ n7654;
  assign n8771 = n8213 & n8770;
  assign n8772 = n8765 & ~n8771;
  assign n8773 = n8232 & n8772;
  assign n8774 = ~n7662 & n8773;
  assign n8775 = n7612 & n8774;
  assign n8776 = n8221 & n8775;
  assign n8777 = n8776 ^ n6178;
  assign n8778 = n8777 ^ x369;
  assign n8779 = n8555 ^ x364;
  assign n8780 = n8778 & n8779;
  assign n8781 = n8069 & ~n8163;
  assign n8782 = n8115 & n8166;
  assign n8783 = ~n8781 & ~n8782;
  assign n8784 = n8108 & n8161;
  assign n8785 = ~n8068 & ~n8522;
  assign n8786 = ~n8784 & ~n8785;
  assign n8787 = ~n8067 & ~n8161;
  assign n8788 = ~n8142 & ~n8787;
  assign n8789 = n8077 ^ n8070;
  assign n8790 = n8789 ^ n8106;
  assign n8791 = n8106 ^ n8077;
  assign n8792 = n8791 ^ n8077;
  assign n8793 = n8105 ^ n8077;
  assign n8794 = n8793 ^ n8077;
  assign n8795 = n8792 & ~n8794;
  assign n8796 = n8795 ^ n8077;
  assign n8797 = n8790 & ~n8796;
  assign n8798 = n8117 & n8797;
  assign n8799 = ~n8788 & ~n8798;
  assign n8800 = n8786 & n8799;
  assign n8801 = n8783 & n8800;
  assign n8802 = n8505 & n8801;
  assign n8803 = ~n8109 & n8802;
  assign n8804 = n8803 ^ n6234;
  assign n8805 = n8804 ^ x368;
  assign n8806 = n8685 ^ x365;
  assign n8807 = n8805 & ~n8806;
  assign n8808 = n6730 & n8325;
  assign n8809 = n6702 & n8329;
  assign n8810 = n8310 & n8809;
  assign n8811 = ~n8808 & ~n8810;
  assign n8812 = n8310 & n8313;
  assign n8813 = n5754 & ~n8812;
  assign n8814 = ~n8308 & n8318;
  assign n8815 = n6719 & ~n8814;
  assign n8816 = ~n8813 & ~n8815;
  assign n8817 = n8811 & n8816;
  assign n8818 = n8817 ^ n6279;
  assign n8819 = n8818 ^ x366;
  assign n8820 = ~n7949 & ~n7967;
  assign n8821 = ~n7957 & ~n8820;
  assign n8822 = ~n7963 & ~n7976;
  assign n8823 = ~n7946 & n8822;
  assign n8824 = n7933 & ~n8823;
  assign n8825 = ~n8821 & ~n8824;
  assign n8826 = ~n7935 & n8822;
  assign n8827 = ~n7927 & n8826;
  assign n8828 = n7952 & ~n8827;
  assign n8829 = ~n7965 & n8342;
  assign n8830 = n8354 & n8829;
  assign n8831 = n7945 & ~n8830;
  assign n8832 = n7933 & ~n7969;
  assign n8833 = ~n7937 & n8822;
  assign n8834 = ~n7958 & n8833;
  assign n8835 = ~n7968 & n8834;
  assign n8836 = n7838 & ~n8835;
  assign n8837 = ~n8832 & ~n8836;
  assign n8838 = ~n8831 & n8837;
  assign n8839 = ~n8828 & n8838;
  assign n8840 = n8825 & n8839;
  assign n8841 = n7931 ^ n7837;
  assign n8842 = n8841 ^ n7931;
  assign n8843 = n7968 ^ n7931;
  assign n8844 = n8842 & n8843;
  assign n8845 = n8844 ^ n7931;
  assign n8846 = ~n7975 & n8845;
  assign n8847 = n8840 & ~n8846;
  assign n8848 = ~n8352 & n8847;
  assign n8849 = n7962 & n8848;
  assign n8850 = n7940 & n8849;
  assign n8851 = n8850 ^ n6312;
  assign n8852 = n8851 ^ x367;
  assign n8853 = ~n8819 & n8852;
  assign n8854 = n8807 & n8853;
  assign n8855 = n8780 & n8854;
  assign n8856 = ~n8778 & ~n8779;
  assign n8857 = n8805 & n8806;
  assign n8858 = n8819 & ~n8852;
  assign n8859 = n8857 & n8858;
  assign n8860 = n8856 & n8859;
  assign n8861 = ~n8855 & ~n8860;
  assign n8862 = ~n8805 & ~n8806;
  assign n8863 = n8853 & n8862;
  assign n8864 = n8780 & n8863;
  assign n8865 = ~n8819 & ~n8852;
  assign n8866 = n8857 & n8865;
  assign n8867 = n8856 & n8866;
  assign n8868 = ~n8864 & ~n8867;
  assign n8869 = ~n8805 & n8806;
  assign n8870 = n8819 & n8869;
  assign n8871 = n8856 & n8870;
  assign n8872 = n8778 & ~n8779;
  assign n8873 = n8859 & n8872;
  assign n8874 = ~n8871 & ~n8873;
  assign n8875 = ~n8778 & n8779;
  assign n8876 = n8866 & n8875;
  assign n8877 = n8819 & n8852;
  assign n8878 = n8807 & n8877;
  assign n8879 = n8858 & n8862;
  assign n8880 = ~n8878 & ~n8879;
  assign n8881 = n8780 & ~n8880;
  assign n8882 = ~n8876 & ~n8881;
  assign n8883 = n8779 ^ n8778;
  assign n8884 = n8857 & n8877;
  assign n8885 = n8853 & n8857;
  assign n8886 = n8865 & n8869;
  assign n8887 = ~n8885 & ~n8886;
  assign n8888 = ~n8884 & n8887;
  assign n8889 = n8883 & ~n8888;
  assign n8890 = ~n8866 & ~n8886;
  assign n8891 = ~n8870 & n8890;
  assign n8892 = n8780 & ~n8891;
  assign n8893 = ~n8854 & ~n8863;
  assign n8894 = n8862 & n8865;
  assign n8895 = ~n8878 & ~n8894;
  assign n8896 = n8893 & n8895;
  assign n8897 = n8856 & ~n8896;
  assign n8898 = ~n8892 & ~n8897;
  assign n8899 = n8862 & n8877;
  assign n8900 = n8807 & n8858;
  assign n8901 = ~n8899 & ~n8900;
  assign n8902 = n8853 & n8869;
  assign n8903 = ~n8894 & ~n8902;
  assign n8904 = n8901 & n8903;
  assign n8905 = n8872 & ~n8904;
  assign n8906 = n8807 & n8865;
  assign n8907 = n8901 & ~n8906;
  assign n8908 = ~n8879 & n8907;
  assign n8909 = n8875 & ~n8908;
  assign n8910 = ~n8905 & ~n8909;
  assign n8911 = n8898 & n8910;
  assign n8912 = ~n8889 & n8911;
  assign n8913 = n8882 & n8912;
  assign n8914 = n8874 & n8913;
  assign n8915 = n8868 & n8914;
  assign n8916 = n8861 & n8915;
  assign n8917 = n8916 ^ n6392;
  assign n8918 = n8917 ^ x422;
  assign n8919 = n8336 ^ x399;
  assign n8920 = n7679 ^ x394;
  assign n8921 = ~n8919 & ~n8920;
  assign n8922 = n8172 ^ x398;
  assign n8923 = n8633 & n8649;
  assign n8924 = n8584 & n8624;
  assign n8925 = ~n8670 & ~n8924;
  assign n8926 = ~n8614 & n8925;
  assign n8927 = n8617 & ~n8926;
  assign n8928 = ~n8923 & ~n8927;
  assign n8929 = n8615 & n8640;
  assign n8930 = n8633 & n8663;
  assign n8931 = ~n8929 & ~n8930;
  assign n8932 = ~n8645 & n8662;
  assign n8933 = ~n8637 & n8926;
  assign n8934 = ~n8646 & n8933;
  assign n8935 = ~n8635 & n8934;
  assign n8936 = n8627 & ~n8935;
  assign n8937 = ~n8932 & ~n8936;
  assign n8938 = ~n8649 & ~n8665;
  assign n8939 = n8622 & ~n8938;
  assign n8940 = ~n8629 & ~n8665;
  assign n8941 = n8650 & n8940;
  assign n8942 = n8617 & ~n8941;
  assign n8943 = ~n8643 & ~n8669;
  assign n8944 = ~n8622 & n8943;
  assign n8945 = ~n8620 & ~n8635;
  assign n8946 = ~n8633 & n8945;
  assign n8947 = n8671 & n8946;
  assign n8948 = ~n8944 & ~n8947;
  assign n8949 = ~n8645 & n8948;
  assign n8950 = ~n8942 & ~n8949;
  assign n8951 = ~n8939 & n8950;
  assign n8952 = n8937 & n8951;
  assign n8953 = n8931 & n8952;
  assign n8954 = n8928 & n8953;
  assign n8955 = ~n8638 & n8954;
  assign n8956 = ~n8636 & n8955;
  assign n8957 = n8632 & n8956;
  assign n8958 = n8957 ^ n6423;
  assign n8959 = n8958 ^ x397;
  assign n8960 = n8922 & n8959;
  assign n8961 = n7741 & n7751;
  assign n8962 = ~n7734 & ~n7784;
  assign n8963 = n7762 & ~n8962;
  assign n8964 = ~n8961 & ~n8963;
  assign n8965 = n7736 & ~n7777;
  assign n8966 = n7684 & ~n7781;
  assign n8967 = ~n8965 & ~n8966;
  assign n8968 = n8964 & n8967;
  assign n8969 = n7685 & ~n7760;
  assign n8970 = n7715 ^ n7686;
  assign n8971 = n8970 ^ n7731;
  assign n8972 = n8971 ^ n7732;
  assign n8973 = n7732 ^ n7731;
  assign n8974 = n7731 ^ n7715;
  assign n8975 = n8974 ^ n7731;
  assign n8976 = ~n8973 & ~n8975;
  assign n8977 = n8976 ^ n7731;
  assign n8978 = n8972 & n8977;
  assign n8979 = ~n7762 & ~n8978;
  assign n8980 = n8979 ^ n7770;
  assign n8981 = ~n7739 & ~n7775;
  assign n8982 = n8981 ^ n8979;
  assign n8983 = n8982 ^ n8981;
  assign n8984 = ~n7752 & ~n7763;
  assign n8985 = n7748 & n8984;
  assign n8986 = n8985 ^ n8981;
  assign n8987 = ~n8983 & ~n8986;
  assign n8988 = n8987 ^ n8981;
  assign n8989 = ~n8980 & n8988;
  assign n8990 = n8989 ^ n7770;
  assign n8991 = ~n8969 & ~n8990;
  assign n8992 = n8968 & n8991;
  assign n8993 = n7750 & n8992;
  assign n8994 = n8464 & n8993;
  assign n8995 = ~n7771 & n8994;
  assign n8996 = ~n7769 & n8995;
  assign n8997 = n8996 ^ n6461;
  assign n8998 = n8997 ^ x396;
  assign n8999 = n7993 ^ x395;
  assign n9000 = ~n8998 & ~n8999;
  assign n9001 = n8960 & n9000;
  assign n9002 = n8921 & n9001;
  assign n9003 = n8919 & n8920;
  assign n9004 = ~n8922 & n8959;
  assign n9005 = n9000 & n9004;
  assign n9006 = n8998 & ~n8999;
  assign n9007 = n8960 & n9006;
  assign n9008 = ~n9005 & ~n9007;
  assign n9009 = n9003 & ~n9008;
  assign n9010 = ~n9002 & ~n9009;
  assign n9011 = ~n8922 & ~n8959;
  assign n9012 = n8998 & n8999;
  assign n9013 = n9011 & n9012;
  assign n9014 = n9003 & n9013;
  assign n9015 = ~n8998 & n8999;
  assign n9016 = n9004 & n9015;
  assign n9017 = n8921 & n9016;
  assign n9018 = n9004 & n9006;
  assign n9019 = n8921 & n9018;
  assign n9020 = ~n8919 & n8920;
  assign n9021 = n8960 & n9015;
  assign n9022 = n8960 & n9012;
  assign n9023 = ~n9021 & ~n9022;
  assign n9024 = n9020 & ~n9023;
  assign n9025 = n8919 & ~n8920;
  assign n9026 = n9006 & n9011;
  assign n9027 = ~n9007 & ~n9026;
  assign n9028 = n9025 & ~n9027;
  assign n9029 = ~n9024 & ~n9028;
  assign n9030 = n9011 & n9015;
  assign n9031 = n9020 & n9030;
  assign n9032 = n9004 & n9012;
  assign n9033 = n8920 & n9032;
  assign n9034 = ~n9031 & ~n9033;
  assign n9035 = ~n9001 & ~n9018;
  assign n9036 = n9025 & ~n9035;
  assign n9037 = n8998 ^ n8959;
  assign n9038 = n9037 ^ n8999;
  assign n9039 = n8999 ^ n8959;
  assign n9040 = n9039 ^ n8959;
  assign n9041 = n8959 ^ n8922;
  assign n9042 = n9041 ^ n8959;
  assign n9043 = n9040 & ~n9042;
  assign n9044 = n9043 ^ n8959;
  assign n9045 = ~n9038 & ~n9044;
  assign n9046 = n9003 & n9045;
  assign n9047 = ~n9036 & ~n9046;
  assign n9048 = n8922 & ~n8959;
  assign n9049 = n9015 & n9048;
  assign n9050 = n9012 & n9048;
  assign n9051 = ~n9030 & ~n9050;
  assign n9052 = n9027 & n9051;
  assign n9053 = ~n9049 & n9052;
  assign n9054 = n8921 & ~n9053;
  assign n9055 = ~n9022 & n9051;
  assign n9056 = ~n9049 & n9055;
  assign n9057 = n9025 & ~n9056;
  assign n9058 = n9006 & n9048;
  assign n9059 = ~n9005 & ~n9058;
  assign n9060 = ~n9026 & n9059;
  assign n9061 = ~n9001 & n9060;
  assign n9062 = n9020 & ~n9061;
  assign n9063 = ~n9057 & ~n9062;
  assign n9064 = ~n9054 & n9063;
  assign n9065 = n9047 & n9064;
  assign n9066 = n9034 & n9065;
  assign n9067 = n9029 & n9066;
  assign n9068 = ~n9019 & n9067;
  assign n9069 = ~n9017 & n9068;
  assign n9070 = ~n9014 & n9069;
  assign n9071 = n9010 & n9070;
  assign n9072 = n9071 ^ n6536;
  assign n9073 = n9072 ^ x421;
  assign n9074 = n8918 & ~n9073;
  assign n9075 = n8751 & n9074;
  assign n9310 = ~n8918 & n9073;
  assign n9076 = n7333 & n7375;
  assign n9077 = n7343 & ~n7379;
  assign n9078 = ~n9076 & ~n9077;
  assign n9079 = n7374 & ~n7390;
  assign n9080 = n7345 & ~n7384;
  assign n9081 = n7354 & n9080;
  assign n9082 = ~n9079 & ~n9081;
  assign n9083 = n7339 & n7343;
  assign n9084 = ~n7352 & ~n7378;
  assign n9085 = n7333 & ~n9084;
  assign n9086 = ~n9083 & ~n9085;
  assign n9087 = n7384 & n8182;
  assign n9088 = ~n7361 & n9087;
  assign n9089 = n9088 ^ n7376;
  assign n9090 = n9089 ^ n7376;
  assign n9091 = n7376 ^ n7164;
  assign n9092 = n9091 ^ n7376;
  assign n9093 = ~n9090 & ~n9092;
  assign n9094 = n9093 ^ n7376;
  assign n9095 = ~n7194 & n9094;
  assign n9096 = n9095 ^ n7376;
  assign n9097 = n9086 & ~n9096;
  assign n9098 = n9082 & n9097;
  assign n9099 = ~n7363 & n9098;
  assign n9100 = n8179 & n9099;
  assign n9101 = n9078 & n9100;
  assign n9102 = n7372 & n9101;
  assign n9103 = n8176 & n9102;
  assign n9104 = ~n7366 & n9103;
  assign n9105 = n7351 & n9104;
  assign n9106 = n9105 ^ n6031;
  assign n9107 = n9106 ^ x381;
  assign n9108 = n7739 & n7751;
  assign n9109 = n7685 & n7741;
  assign n9110 = ~n7776 & ~n7785;
  assign n9111 = n7762 & ~n9110;
  assign n9112 = n8470 & n8482;
  assign n9113 = ~n7746 & n9112;
  assign n9114 = ~n7739 & n9113;
  assign n9115 = n7736 & ~n9114;
  assign n9116 = ~n9111 & ~n9115;
  assign n9117 = ~n7684 & n7784;
  assign n9118 = ~n7747 & ~n7752;
  assign n9119 = n7770 & ~n9118;
  assign n9120 = ~n7758 & n8984;
  assign n9121 = n9120 ^ n7684;
  assign n9122 = n9121 ^ n9120;
  assign n9123 = ~n7746 & n7782;
  assign n9124 = n9123 ^ n9120;
  assign n9125 = ~n9122 & n9124;
  assign n9126 = n9125 ^ n9120;
  assign n9127 = ~n7683 & ~n9126;
  assign n9128 = ~n9119 & ~n9127;
  assign n9129 = ~n9117 & n9128;
  assign n9130 = n9116 & n9129;
  assign n9131 = n8476 & n9130;
  assign n9132 = ~n7735 & n9131;
  assign n9133 = ~n9109 & n9132;
  assign n9134 = ~n9108 & n9133;
  assign n9135 = n8469 & n9134;
  assign n9136 = n8466 & n9135;
  assign n9137 = ~n7767 & n9136;
  assign n9138 = ~n7771 & n9137;
  assign n9139 = n9138 ^ n6087;
  assign n9140 = n9139 ^ x376;
  assign n9141 = n9107 & n9140;
  assign n9142 = n5754 & ~n6716;
  assign n9143 = n6719 & ~n6740;
  assign n9144 = ~n9142 & ~n9143;
  assign n9145 = n6700 ^ n5376;
  assign n9146 = n9145 ^ n6700;
  assign n9147 = n6728 ^ n6700;
  assign n9148 = n9146 & ~n9147;
  assign n9149 = n9148 ^ n6700;
  assign n9150 = ~n5753 & ~n9149;
  assign n9151 = n9144 & ~n9150;
  assign n9152 = n9151 ^ n5772;
  assign n9153 = n9152 ^ x380;
  assign n9154 = n7623 & ~n7645;
  assign n9155 = ~n7552 & ~n7644;
  assign n9156 = ~n7622 & n9155;
  assign n9157 = n7629 & ~n9156;
  assign n9158 = ~n9154 & ~n9157;
  assign n9159 = ~n7639 & ~n7652;
  assign n9160 = ~n7610 & n9159;
  assign n9161 = n7606 & ~n9160;
  assign n9162 = n7641 & ~n7652;
  assign n9163 = ~n7622 & n9162;
  assign n9164 = n7608 & ~n9163;
  assign n9165 = ~n9161 & ~n9164;
  assign n9166 = n9158 & n9165;
  assign n9167 = ~n7638 & n9166;
  assign n9168 = n7633 & n9167;
  assign n9169 = ~n8771 & n9168;
  assign n9170 = n8227 & n9169;
  assign n9171 = n8223 & n9170;
  assign n9172 = ~n7615 & n9171;
  assign n9173 = n7612 & n9172;
  assign n9174 = n8221 & n9173;
  assign n9175 = n9174 ^ n5842;
  assign n9176 = n9175 ^ x378;
  assign n9177 = ~n9153 & ~n9176;
  assign n9178 = ~n8646 & n8650;
  assign n9179 = n8622 & ~n9178;
  assign n9180 = ~n8662 & n8666;
  assign n9181 = n8633 & ~n9180;
  assign n9182 = ~n8622 & ~n8670;
  assign n9183 = ~n8614 & n8946;
  assign n9184 = ~n9182 & ~n9183;
  assign n9185 = ~n8643 & ~n9184;
  assign n9186 = ~n8645 & ~n9185;
  assign n9187 = ~n9181 & ~n9186;
  assign n9188 = ~n9179 & n9187;
  assign n9189 = n8616 ^ n8615;
  assign n9190 = n8664 & ~n8669;
  assign n9191 = ~n8635 & n9190;
  assign n9192 = n9191 ^ n8616;
  assign n9193 = n9192 ^ n9191;
  assign n9194 = n8651 & n8672;
  assign n9195 = ~n8620 & n9194;
  assign n9196 = n9195 ^ n9191;
  assign n9197 = ~n9193 & n9196;
  assign n9198 = n9197 ^ n9191;
  assign n9199 = n9189 & ~n9198;
  assign n9200 = n9188 & ~n9199;
  assign n9201 = n8631 & n9200;
  assign n9202 = n8642 & n9201;
  assign n9203 = n8928 & n9202;
  assign n9204 = ~n8638 & n9203;
  assign n9205 = n9204 ^ n5993;
  assign n9206 = n9205 ^ x377;
  assign n9207 = n7927 & n7945;
  assign n9208 = n7838 & n7964;
  assign n9209 = n7937 & ~n7957;
  assign n9210 = ~n7935 & ~n7958;
  assign n9211 = ~n7967 & n9210;
  assign n9212 = n7933 & ~n9211;
  assign n9213 = ~n9209 & ~n9212;
  assign n9214 = n8822 & n8829;
  assign n9215 = ~n7949 & n9214;
  assign n9216 = n7952 & ~n9215;
  assign n9217 = n7938 & ~n7968;
  assign n9218 = ~n7949 & n9217;
  assign n9219 = n7838 & ~n9218;
  assign n9220 = ~n9216 & ~n9219;
  assign n9221 = n7945 & ~n8342;
  assign n9222 = ~n7942 & ~n7963;
  assign n9223 = n7933 & ~n9222;
  assign n9224 = ~n9221 & ~n9223;
  assign n9225 = n7955 & n9224;
  assign n9226 = ~n7836 & ~n9225;
  assign n9227 = n9220 & ~n9226;
  assign n9228 = n9213 & n9227;
  assign n9229 = ~n9208 & n9228;
  assign n9230 = ~n9207 & n9229;
  assign n9231 = ~n7961 & n9230;
  assign n9232 = n8340 & n9231;
  assign n9233 = ~n8846 & n9232;
  assign n9234 = ~n7928 & n9233;
  assign n9235 = n9234 ^ n5812;
  assign n9236 = n9235 ^ x379;
  assign n9237 = ~n9206 & ~n9236;
  assign n9238 = n9177 & n9237;
  assign n9239 = n9141 & n9238;
  assign n9240 = n9107 & ~n9140;
  assign n9241 = ~n9153 & n9176;
  assign n9242 = n9206 & n9236;
  assign n9243 = n9241 & n9242;
  assign n9244 = n9153 & n9176;
  assign n9245 = n9206 & ~n9236;
  assign n9246 = n9244 & n9245;
  assign n9247 = ~n9243 & ~n9246;
  assign n9248 = n9240 & ~n9247;
  assign n9249 = ~n9239 & ~n9248;
  assign n9250 = ~n9107 & n9140;
  assign n9251 = n9177 & n9245;
  assign n9252 = ~n9246 & ~n9251;
  assign n9253 = n9250 & ~n9252;
  assign n9254 = n9242 & n9244;
  assign n9255 = ~n9107 & n9254;
  assign n9256 = n9177 & n9242;
  assign n9257 = n9250 & n9256;
  assign n9258 = ~n9255 & ~n9257;
  assign n9259 = n9153 & ~n9176;
  assign n9260 = n9242 & n9259;
  assign n9261 = ~n9256 & ~n9260;
  assign n9262 = n9240 & ~n9261;
  assign n9263 = ~n9206 & n9236;
  assign n9264 = n9244 & n9263;
  assign n9265 = n9141 & n9264;
  assign n9266 = n9177 & n9263;
  assign n9267 = n9250 & n9266;
  assign n9268 = n9237 & n9259;
  assign n9269 = n9240 & n9268;
  assign n9270 = ~n9267 & ~n9269;
  assign n9271 = ~n9107 & ~n9140;
  assign n9272 = n9245 & n9259;
  assign n9273 = ~n9251 & ~n9272;
  assign n9274 = n9271 & ~n9273;
  assign n9275 = ~n9141 & ~n9271;
  assign n9276 = ~n9206 & n9241;
  assign n9277 = n9236 & n9276;
  assign n9278 = n9237 & n9244;
  assign n9279 = ~n9277 & ~n9278;
  assign n9280 = n9241 & n9245;
  assign n9281 = n9259 & n9263;
  assign n9282 = ~n9260 & ~n9272;
  assign n9283 = ~n9281 & n9282;
  assign n9284 = ~n9280 & n9283;
  assign n9285 = n9279 & n9284;
  assign n9286 = ~n9275 & ~n9285;
  assign n9287 = n9250 ^ n9240;
  assign n9289 = ~n9236 & n9276;
  assign n9290 = ~n9264 & ~n9289;
  assign n9291 = ~n9268 & n9290;
  assign n9288 = ~n9238 & ~n9276;
  assign n9292 = n9291 ^ n9288;
  assign n9293 = n9291 ^ n9240;
  assign n9294 = n9293 ^ n9291;
  assign n9295 = ~n9292 & n9294;
  assign n9296 = n9295 ^ n9291;
  assign n9297 = n9287 & n9296;
  assign n9298 = n9297 ^ n9250;
  assign n9299 = ~n9286 & ~n9298;
  assign n9300 = ~n9274 & n9299;
  assign n9301 = n9270 & n9300;
  assign n9302 = ~n9265 & n9301;
  assign n9303 = ~n9262 & n9302;
  assign n9304 = n9258 & n9303;
  assign n9305 = ~n9253 & n9304;
  assign n9306 = n9249 & n9305;
  assign n9307 = n9306 ^ n6160;
  assign n9308 = n9307 ^ x420;
  assign n9309 = ~n8751 & n9308;
  assign n9311 = n9310 ^ n9309;
  assign n9312 = ~n9075 & ~n9311;
  assign n9313 = n8460 & ~n9312;
  assign n9314 = n8066 & n8459;
  assign n9315 = ~n8751 & ~n9308;
  assign n9316 = n9073 & n9315;
  assign n9317 = n8918 & n9073;
  assign n9318 = ~n8918 & ~n9073;
  assign n9319 = ~n9317 & ~n9318;
  assign n9320 = n9308 & ~n9319;
  assign n9321 = ~n9316 & ~n9320;
  assign n9322 = n9074 ^ n9073;
  assign n9323 = ~n9308 & n9322;
  assign n9324 = n9323 ^ n9073;
  assign n9325 = n8751 & n9324;
  assign n9326 = n9321 & ~n9325;
  assign n9327 = n9314 & ~n9326;
  assign n9328 = ~n9313 & ~n9327;
  assign n9329 = ~n8066 & n8459;
  assign n9330 = n9308 ^ n8918;
  assign n9331 = n9330 ^ n8918;
  assign n9332 = n8918 ^ n8751;
  assign n9333 = n9332 ^ n9308;
  assign n9334 = n9333 ^ n8918;
  assign n9335 = n9334 ^ n8918;
  assign n9336 = n9331 & ~n9335;
  assign n9337 = n9336 ^ n8918;
  assign n9338 = n9073 & n9337;
  assign n9339 = n9338 ^ n9333;
  assign n9340 = n9329 & n9339;
  assign n9341 = n8751 & n9308;
  assign n9342 = n9310 & n9341;
  assign n9343 = n8066 & ~n8459;
  assign n9344 = ~n8751 & n9318;
  assign n9345 = n8751 & n9317;
  assign n9346 = ~n9315 & ~n9341;
  assign n9347 = n8918 & ~n9346;
  assign n9348 = ~n9345 & ~n9347;
  assign n9349 = ~n9344 & n9348;
  assign n9350 = n9343 & ~n9349;
  assign n9351 = ~n9342 & ~n9350;
  assign n9352 = ~n9340 & n9351;
  assign n9353 = n9328 & n9352;
  assign n9354 = n9353 ^ n8336;
  assign n9355 = n9354 ^ x449;
  assign n9356 = n9152 ^ x382;
  assign n9357 = n7130 ^ x387;
  assign n9358 = ~n9356 & ~n9357;
  assign n9359 = n9106 ^ x383;
  assign n9360 = n8622 & n8640;
  assign n9361 = n8615 & n8646;
  assign n9362 = ~n9360 & ~n9361;
  assign n9363 = n8617 & ~n8672;
  assign n9364 = n8633 & n8662;
  assign n9365 = ~n8620 & n8940;
  assign n9366 = n9365 ^ n8663;
  assign n9367 = ~n9189 & ~n9366;
  assign n9368 = n9367 ^ n8663;
  assign n9369 = n8625 ^ n8617;
  assign n9370 = n8627 ^ n8625;
  assign n9371 = n9370 ^ n8627;
  assign n9372 = n8650 ^ n8627;
  assign n9373 = ~n9371 & n9372;
  assign n9374 = n9373 ^ n8627;
  assign n9375 = n9369 & n9374;
  assign n9376 = n9375 ^ n8617;
  assign n9377 = ~n9368 & ~n9376;
  assign n9378 = n8622 & ~n8926;
  assign n9379 = ~n8637 & ~n8643;
  assign n9380 = ~n8614 & n9379;
  assign n9381 = n8627 & ~n9380;
  assign n9382 = ~n8923 & ~n9381;
  assign n9383 = ~n8669 & n9382;
  assign n9384 = n8615 & ~n9383;
  assign n9385 = ~n9378 & ~n9384;
  assign n9386 = n9377 & n9385;
  assign n9387 = ~n8636 & n9386;
  assign n9388 = ~n9364 & n9387;
  assign n9389 = ~n9363 & n9388;
  assign n9390 = n9362 & n9389;
  assign n9391 = n8632 & n9390;
  assign n9392 = n9391 ^ n6952;
  assign n9393 = n9392 ^ x385;
  assign n9394 = ~n9359 & n9393;
  assign n9395 = n7805 ^ x386;
  assign n9396 = n8117 & ~n8162;
  assign n9397 = n8136 & ~n8515;
  assign n9398 = n8161 & ~n9397;
  assign n9399 = ~n9396 & ~n9398;
  assign n9400 = n8067 & n8139;
  assign n9401 = ~n8157 & ~n8500;
  assign n9402 = n8115 & ~n9401;
  assign n9415 = ~n8108 & ~n8111;
  assign n9413 = ~n8135 & ~n8515;
  assign n9414 = ~n8129 & n9413;
  assign n9416 = n9415 ^ n9414;
  assign n9405 = n8068 ^ n8067;
  assign n9406 = n9405 ^ n8067;
  assign n9417 = n9414 ^ n8067;
  assign n9418 = n9406 & n9417;
  assign n9419 = n9418 ^ n8067;
  assign n9420 = n9416 & n9419;
  assign n9421 = n9420 ^ n9415;
  assign n9422 = ~n8500 & n9421;
  assign n9403 = n8142 & ~n8154;
  assign n9404 = n9403 ^ n8523;
  assign n9407 = n9403 ^ n8067;
  assign n9408 = ~n9406 & n9407;
  assign n9409 = n9408 ^ n8067;
  assign n9410 = n9404 & n9409;
  assign n9411 = n9410 ^ n8523;
  assign n9412 = ~n8129 & n9411;
  assign n9423 = n9422 ^ n9412;
  assign n9424 = n8068 & n9423;
  assign n9425 = n9424 ^ n9422;
  assign n9426 = ~n8510 & n9425;
  assign n9427 = ~n9402 & n9426;
  assign n9428 = ~n9400 & n9427;
  assign n9429 = n9399 & n9428;
  assign n9430 = n8509 & n9429;
  assign n9431 = n8127 & n9430;
  assign n9432 = ~n8109 & n9431;
  assign n9433 = n9432 ^ n6925;
  assign n9434 = n9433 ^ x384;
  assign n9435 = n9395 & ~n9434;
  assign n9436 = n9394 & n9435;
  assign n9437 = ~n9359 & ~n9393;
  assign n9438 = ~n9395 & ~n9434;
  assign n9439 = n9437 & n9438;
  assign n9440 = ~n9436 & ~n9439;
  assign n9441 = n9358 & ~n9440;
  assign n9442 = n9356 & n9357;
  assign n9443 = ~n9440 & n9442;
  assign n9444 = n9356 & ~n9357;
  assign n9445 = n9359 & n9393;
  assign n9446 = n9438 & n9445;
  assign n9447 = n9359 & ~n9393;
  assign n9448 = n9435 & n9447;
  assign n9449 = ~n9446 & ~n9448;
  assign n9450 = n9444 & ~n9449;
  assign n9451 = n9395 & n9434;
  assign n9452 = n9394 & n9451;
  assign n9453 = ~n9395 & n9434;
  assign n9454 = n9447 & n9453;
  assign n9455 = ~n9452 & ~n9454;
  assign n9456 = n9358 & ~n9455;
  assign n9457 = ~n9450 & ~n9456;
  assign n9458 = ~n9443 & n9457;
  assign n9459 = n9442 & n9452;
  assign n9460 = n9444 & n9454;
  assign n9461 = ~n9459 & ~n9460;
  assign n9462 = n9394 & n9438;
  assign n9463 = n9444 & n9462;
  assign n9464 = n9357 ^ n9356;
  assign n9465 = n9445 & n9453;
  assign n9466 = n9445 & n9451;
  assign n9467 = n9437 & n9451;
  assign n9468 = n9435 & n9437;
  assign n9469 = ~n9467 & ~n9468;
  assign n9470 = ~n9466 & n9469;
  assign n9471 = ~n9465 & n9470;
  assign n9472 = n9464 & ~n9471;
  assign n9473 = ~n9463 & ~n9472;
  assign n9474 = n9394 & n9453;
  assign n9475 = n9442 & n9474;
  assign n9476 = ~n9356 & n9357;
  assign n9477 = ~n9434 & n9447;
  assign n9478 = n9437 & n9453;
  assign n9479 = ~n9477 & ~n9478;
  assign n9480 = ~n9474 & n9479;
  assign n9481 = n9476 & ~n9480;
  assign n9482 = n9438 & n9447;
  assign n9483 = n9447 & n9451;
  assign n9484 = ~n9482 & ~n9483;
  assign n9485 = ~n9464 & ~n9484;
  assign n9486 = ~n9446 & ~n9454;
  assign n9487 = n9442 & ~n9486;
  assign n9488 = n9435 & n9445;
  assign n9489 = ~n9465 & ~n9488;
  assign n9490 = n9358 & ~n9489;
  assign n9491 = ~n9487 & ~n9490;
  assign n9492 = ~n9485 & n9491;
  assign n9493 = ~n9481 & n9492;
  assign n9494 = ~n9475 & n9493;
  assign n9495 = n9473 & n9494;
  assign n9496 = n9461 & n9495;
  assign n9497 = n9458 & n9496;
  assign n9498 = ~n9441 & n9497;
  assign n9499 = n9498 ^ n7604;
  assign n9500 = n9499 ^ x406;
  assign n9501 = n8211 & n8398;
  assign n9502 = ~n8456 & ~n9501;
  assign n9503 = ~n8379 & ~n8400;
  assign n9504 = ~n8398 & n9503;
  assign n9505 = n8389 & ~n9504;
  assign n9506 = ~n8422 & ~n8425;
  assign n9507 = ~n8382 & n9506;
  assign n9508 = n8381 & ~n9507;
  assign n9509 = ~n9505 & ~n9508;
  assign n9510 = ~n8415 & ~n8422;
  assign n9511 = n8211 & ~n9510;
  assign n9512 = ~n8415 & ~n8433;
  assign n9513 = n8389 & ~n9512;
  assign n9514 = ~n8413 & ~n9513;
  assign n9515 = n8211 & n8382;
  assign n9516 = n8389 & ~n8406;
  assign n9517 = ~n8387 & n8409;
  assign n9518 = n8381 & ~n9517;
  assign n9519 = ~n8390 & n8436;
  assign n9520 = n8426 & n9519;
  assign n9521 = n8385 & ~n9520;
  assign n9522 = ~n9518 & ~n9521;
  assign n9523 = ~n9516 & n9522;
  assign n9524 = ~n9515 & n9523;
  assign n9525 = n9514 & n9524;
  assign n9526 = ~n8376 & n9525;
  assign n9527 = ~n8392 & n9526;
  assign n9528 = ~n9511 & n9527;
  assign n9529 = n9509 & n9528;
  assign n9530 = n9502 & n9529;
  assign n9531 = n9530 ^ n7572;
  assign n9532 = n9531 ^ x411;
  assign n9533 = n9500 & n9532;
  assign n9534 = n8029 & ~n8050;
  assign n9535 = n8025 & ~n9534;
  assign n9536 = ~n8033 & ~n8053;
  assign n9537 = n8016 & ~n9536;
  assign n9538 = n8027 & ~n8030;
  assign n9539 = ~n9537 & ~n9538;
  assign n9540 = n7994 ^ n7806;
  assign n9541 = n8023 ^ n7994;
  assign n9542 = n9541 ^ n8023;
  assign n9543 = n7998 & n8009;
  assign n9544 = ~n8002 & ~n9543;
  assign n9545 = n9544 ^ n8023;
  assign n9546 = ~n9542 & ~n9545;
  assign n9547 = n9546 ^ n8023;
  assign n9548 = ~n9540 & n9547;
  assign n9560 = ~n8016 & ~n8026;
  assign n9561 = ~n7682 & n9560;
  assign n9562 = ~n8026 & ~n9543;
  assign n9563 = n8055 & n9562;
  assign n9564 = ~n7999 & n9563;
  assign n9565 = ~n9561 & ~n9564;
  assign n9566 = n9536 & ~n9565;
  assign n9549 = n7132 & n8001;
  assign n9550 = n8019 ^ n7994;
  assign n9551 = n9550 ^ n8019;
  assign n9552 = ~n8017 & ~n8018;
  assign n9553 = n9552 ^ n8019;
  assign n9554 = ~n9551 & n9553;
  assign n9555 = n9554 ^ n8019;
  assign n9556 = n9540 & ~n9555;
  assign n9557 = ~n8032 & ~n9556;
  assign n9558 = ~n9549 & n9557;
  assign n9559 = ~n7999 & n9558;
  assign n9567 = n9566 ^ n9559;
  assign n9568 = ~n8030 & n9567;
  assign n9569 = n9568 ^ n9566;
  assign n9570 = ~n9548 & n9569;
  assign n9571 = n9539 & n9570;
  assign n9572 = n8015 & n9571;
  assign n9573 = n9535 & n9572;
  assign n9574 = n9573 ^ n7549;
  assign n9575 = n9574 ^ x409;
  assign n9576 = n8921 & n9058;
  assign n9577 = n9020 & n9058;
  assign n9578 = ~n9032 & ~n9050;
  assign n9579 = n9025 & ~n9578;
  assign n9580 = ~n9577 & ~n9579;
  assign n9581 = ~n9576 & n9580;
  assign n9582 = n9025 & n9030;
  assign n9583 = n9003 & n9018;
  assign n9584 = ~n9582 & ~n9583;
  assign n9585 = n9000 & n9011;
  assign n9586 = n9020 & n9585;
  assign n9587 = n9021 & n9025;
  assign n9588 = n9016 & n9020;
  assign n9589 = n9003 & n9049;
  assign n9590 = ~n9588 & ~n9589;
  assign n9591 = n9013 & n9020;
  assign n9592 = n8920 & n9005;
  assign n9593 = ~n9591 & ~n9592;
  assign n9594 = n9022 ^ n8921;
  assign n9595 = n9022 ^ n9003;
  assign n9596 = n9595 ^ n9003;
  assign n9597 = n9051 ^ n9003;
  assign n9598 = ~n9596 & n9597;
  assign n9599 = n9598 ^ n9003;
  assign n9600 = n9594 & n9599;
  assign n9601 = n9600 ^ n8921;
  assign n9602 = n9593 & ~n9601;
  assign n9603 = n8920 ^ n8919;
  assign n9604 = ~n9001 & ~n9032;
  assign n9605 = ~n9603 & ~n9604;
  assign n9606 = n9000 & n9048;
  assign n9607 = n9606 ^ n9025;
  assign n9608 = n9607 ^ n9606;
  assign n9609 = n9606 ^ n9059;
  assign n9610 = n9608 & ~n9609;
  assign n9611 = n9610 ^ n9606;
  assign n9612 = ~n9605 & ~n9611;
  assign n9613 = n9602 & n9612;
  assign n9614 = n9590 & n9613;
  assign n9615 = n9029 & n9614;
  assign n9616 = ~n9014 & n9615;
  assign n9617 = ~n9587 & n9616;
  assign n9618 = ~n9586 & n9617;
  assign n9619 = n9584 & n9618;
  assign n9620 = n9581 & n9619;
  assign n9621 = ~n9019 & n9620;
  assign n9622 = n9621 ^ n7438;
  assign n9623 = n9622 ^ x407;
  assign n9624 = n9575 & ~n9623;
  assign n9625 = n8863 & n8872;
  assign n9626 = n8852 & n8870;
  assign n9627 = ~n8885 & ~n9626;
  assign n9628 = n8856 & ~n9627;
  assign n9629 = ~n8859 & ~n8886;
  assign n9630 = n8780 & ~n9629;
  assign n9631 = ~n9628 & ~n9630;
  assign n9632 = n8780 & n8899;
  assign n9633 = n8861 & ~n9632;
  assign n9634 = n8875 & n8879;
  assign n9635 = ~n8852 & n8870;
  assign n9636 = ~n8863 & ~n8906;
  assign n9637 = ~n9635 & n9636;
  assign n9638 = ~n8884 & n9637;
  assign n9639 = n8780 & ~n9638;
  assign n9640 = n8872 & n8884;
  assign n9641 = n8875 & n8902;
  assign n9642 = ~n9640 & ~n9641;
  assign n9643 = n8819 ^ n8805;
  assign n9644 = n9643 ^ n8806;
  assign n9645 = n8852 ^ n8806;
  assign n9646 = n8819 ^ n8806;
  assign n9647 = n9645 & ~n9646;
  assign n9648 = ~n9644 & n9647;
  assign n9649 = n9648 ^ n9644;
  assign n9650 = n8883 & ~n9649;
  assign n9651 = ~n8879 & ~n8902;
  assign n9652 = n9636 & n9651;
  assign n9653 = ~n8878 & n9652;
  assign n9654 = n8856 & ~n9653;
  assign n9655 = ~n9650 & ~n9654;
  assign n9656 = n9642 & n9655;
  assign n9657 = ~n9639 & n9656;
  assign n9658 = ~n9634 & n9657;
  assign n9659 = n9633 & n9658;
  assign n9660 = n9631 & n9659;
  assign n9661 = ~n9625 & n9660;
  assign n9662 = n9661 ^ n7472;
  assign n9663 = n9662 ^ x408;
  assign n9664 = n9240 & n9266;
  assign n9665 = n9141 & ~n9247;
  assign n9666 = ~n9664 & ~n9665;
  assign n9667 = ~n9238 & n9290;
  assign n9668 = n9271 & ~n9667;
  assign n9669 = n9141 & ~n9273;
  assign n9670 = ~n9668 & ~n9669;
  assign n9671 = n9240 & n9281;
  assign n9672 = ~n9140 & n9277;
  assign n9673 = n9141 & n9266;
  assign n9674 = ~n9254 & ~n9280;
  assign n9675 = n9250 & ~n9674;
  assign n9676 = ~n9673 & ~n9675;
  assign n9677 = ~n9260 & n9279;
  assign n9678 = n9250 & ~n9677;
  assign n9679 = ~n9238 & ~n9278;
  assign n9680 = ~n9281 & n9679;
  assign n9681 = n9141 & ~n9680;
  assign n9682 = ~n9678 & ~n9681;
  assign n9683 = n9261 & ~n9272;
  assign n9684 = ~n9280 & n9683;
  assign n9685 = n9271 & ~n9684;
  assign n9686 = ~n9251 & ~n9256;
  assign n9687 = ~n9289 & n9686;
  assign n9688 = ~n9254 & n9687;
  assign n9689 = n9240 & ~n9688;
  assign n9690 = ~n9685 & ~n9689;
  assign n9691 = n9682 & n9690;
  assign n9692 = n9676 & n9691;
  assign n9693 = ~n9253 & n9692;
  assign n9694 = ~n9672 & n9693;
  assign n9695 = ~n9671 & n9694;
  assign n9696 = n9670 & n9695;
  assign n9697 = n9666 & n9696;
  assign n9698 = n9270 & n9697;
  assign n9699 = n9698 ^ n7515;
  assign n9700 = n9699 ^ x410;
  assign n9701 = n9663 & ~n9700;
  assign n9702 = n9624 & n9701;
  assign n9703 = n9533 & n9702;
  assign n9704 = n9500 & ~n9532;
  assign n9705 = ~n9575 & ~n9623;
  assign n9706 = n9663 & n9700;
  assign n9707 = n9705 & n9706;
  assign n9708 = ~n9663 & ~n9700;
  assign n9709 = n9705 & n9708;
  assign n9710 = ~n9707 & ~n9709;
  assign n9711 = n9704 & ~n9710;
  assign n9712 = ~n9703 & ~n9711;
  assign n9713 = ~n9575 & n9623;
  assign n9714 = n9701 & n9713;
  assign n9715 = n9704 & n9714;
  assign n9716 = ~n9500 & n9532;
  assign n9717 = n9706 & n9713;
  assign n9718 = n9575 & n9623;
  assign n9719 = n9708 & n9718;
  assign n9720 = ~n9717 & ~n9719;
  assign n9721 = ~n9702 & n9720;
  assign n9722 = n9716 & ~n9721;
  assign n9723 = ~n9715 & ~n9722;
  assign n9724 = ~n9663 & n9700;
  assign n9725 = n9713 & n9724;
  assign n9726 = ~n9719 & ~n9725;
  assign n9727 = n9704 & ~n9726;
  assign n9728 = ~n9500 & ~n9532;
  assign n9729 = n9717 & n9728;
  assign n9730 = n9701 & n9718;
  assign n9731 = n9728 & n9730;
  assign n9732 = ~n9729 & ~n9731;
  assign n9733 = n9624 & n9706;
  assign n9734 = ~n9714 & ~n9733;
  assign n9735 = n9728 & ~n9734;
  assign n9736 = n9705 & n9724;
  assign n9737 = n9708 & n9713;
  assign n9738 = n9624 & n9708;
  assign n9739 = ~n9737 & ~n9738;
  assign n9740 = ~n9736 & n9739;
  assign n9741 = ~n9500 & ~n9740;
  assign n9742 = ~n9735 & ~n9741;
  assign n9743 = ~n9702 & ~n9737;
  assign n9744 = ~n9733 & n9743;
  assign n9745 = n9704 & ~n9744;
  assign n9746 = n9706 & n9718;
  assign n9747 = ~n9725 & ~n9746;
  assign n9748 = n9716 & ~n9747;
  assign n9749 = n9718 & n9724;
  assign n9750 = n9532 ^ n9500;
  assign n9751 = n9749 & ~n9750;
  assign n9752 = n9663 ^ n9623;
  assign n9753 = n9575 & ~n9700;
  assign n9754 = ~n9752 & n9753;
  assign n9755 = n9754 ^ n9752;
  assign n9756 = n9533 & ~n9755;
  assign n9757 = ~n9751 & ~n9756;
  assign n9758 = ~n9748 & n9757;
  assign n9759 = ~n9745 & n9758;
  assign n9760 = n9742 & n9759;
  assign n9761 = n9732 & n9760;
  assign n9762 = ~n9727 & n9761;
  assign n9763 = n9723 & n9762;
  assign n9764 = n9712 & n9763;
  assign n9765 = n9764 ^ n8257;
  assign n9766 = n9765 ^ x450;
  assign n9767 = n9355 & n9766;
  assign n9768 = n8917 ^ x424;
  assign n9769 = n8921 & n9022;
  assign n9770 = ~n9018 & ~n9606;
  assign n9771 = n9025 & ~n9770;
  assign n9772 = ~n9769 & ~n9771;
  assign n9773 = n9003 & n9026;
  assign n9774 = ~n9016 & ~n9058;
  assign n9775 = n9025 & ~n9774;
  assign n9776 = ~n9773 & ~n9775;
  assign n9777 = n8920 & n9021;
  assign n9778 = ~n9013 & ~n9606;
  assign n9779 = n8921 & ~n9778;
  assign n9780 = n9022 & n9025;
  assign n9781 = n9020 & ~n9052;
  assign n9782 = ~n9780 & ~n9781;
  assign n9783 = n9603 ^ n9585;
  assign n9784 = n9585 ^ n8920;
  assign n9785 = n9784 ^ n8920;
  assign n9786 = n9049 ^ n8920;
  assign n9787 = ~n9785 & ~n9786;
  assign n9788 = n9787 ^ n8920;
  assign n9789 = ~n9783 & ~n9788;
  assign n9790 = n9789 ^ n9585;
  assign n9791 = n9782 & ~n9790;
  assign n9792 = ~n9779 & n9791;
  assign n9793 = ~n9777 & n9792;
  assign n9794 = n9776 & n9793;
  assign n9795 = ~n9588 & n9794;
  assign n9796 = n9580 & n9795;
  assign n9797 = n9584 & n9796;
  assign n9798 = n9772 & n9797;
  assign n9799 = ~n9019 & n9798;
  assign n9800 = ~n9017 & n9799;
  assign n9801 = ~n9014 & n9800;
  assign n9802 = n9010 & n9801;
  assign n9803 = n9802 ^ n6780;
  assign n9804 = n9803 ^ x429;
  assign n9805 = n9768 & n9804;
  assign n9806 = n8804 ^ x370;
  assign n9807 = n9205 ^ x375;
  assign n9808 = n9806 & ~n9807;
  assign n9809 = n8777 ^ x371;
  assign n9810 = n7067 & ~n7078;
  assign n9811 = n7080 & ~n7116;
  assign n9812 = ~n9810 & ~n9811;
  assign n9813 = ~n7104 & ~n7113;
  assign n9814 = n7072 & ~n9813;
  assign n9817 = ~n7030 & n7090;
  assign n9818 = ~n7104 & ~n9817;
  assign n9815 = ~n7069 & n7114;
  assign n9816 = ~n7081 & n9815;
  assign n9819 = n9818 ^ n9816;
  assign n9820 = n9818 ^ n7080;
  assign n9821 = n9820 ^ n9818;
  assign n9822 = ~n9819 & n9821;
  assign n9823 = n9822 ^ n9818;
  assign n9824 = n8273 & n9823;
  assign n9825 = n9824 ^ n7067;
  assign n9826 = ~n9814 & ~n9825;
  assign n9827 = ~n6781 & n7089;
  assign n9830 = ~n7106 & n8264;
  assign n9828 = ~n7085 & ~n7091;
  assign n9829 = ~n7065 & n9828;
  assign n9831 = n9830 ^ n9829;
  assign n9832 = n6781 ^ n6746;
  assign n9833 = n9829 ^ n6781;
  assign n9834 = n9832 & n9833;
  assign n9835 = n9834 ^ n6781;
  assign n9836 = n9831 & n9835;
  assign n9837 = n9836 ^ n9830;
  assign n9838 = ~n7077 & n9837;
  assign n9839 = ~n8263 & ~n9838;
  assign n9840 = ~n9827 & ~n9839;
  assign n9841 = n9826 & n9840;
  assign n9842 = n9812 & n9841;
  assign n9843 = ~n8299 & n9842;
  assign n9844 = n8538 & n9843;
  assign n9845 = n7071 & n9844;
  assign n9846 = n9845 ^ n6804;
  assign n9847 = n9846 ^ x372;
  assign n9848 = ~n9809 & n9847;
  assign n9849 = ~n7164 & n7383;
  assign n9850 = n7329 ^ n7230;
  assign n9851 = n9850 ^ n7230;
  assign n9852 = n7292 ^ n7230;
  assign n9853 = n9852 ^ n7230;
  assign n9854 = ~n9851 & n9853;
  assign n9855 = n9854 ^ n7230;
  assign n9856 = n7262 & ~n9855;
  assign n9857 = ~n7383 & ~n9856;
  assign n9858 = ~n7331 & n9857;
  assign n9859 = n7333 & ~n9858;
  assign n9860 = ~n9849 & ~n9859;
  assign n9861 = n7336 & n7343;
  assign n9862 = ~n7348 & ~n7374;
  assign n9863 = n7354 & ~n9862;
  assign n9864 = n7354 & ~n8182;
  assign n9865 = ~n7356 & n7377;
  assign n9866 = ~n7331 & n9865;
  assign n9867 = n7343 & ~n9866;
  assign n9868 = ~n7361 & ~n9856;
  assign n9869 = n7195 & ~n9868;
  assign n9870 = ~n9867 & ~n9869;
  assign n9871 = ~n9864 & n9870;
  assign n9872 = n7360 & n9871;
  assign n9873 = ~n9863 & n9872;
  assign n9874 = ~n9861 & n9873;
  assign n9875 = n9860 & n9874;
  assign n9876 = ~n7332 & n9875;
  assign n9877 = n9078 & n9876;
  assign n9878 = n7364 & n9877;
  assign n9879 = n9878 ^ n6835;
  assign n9880 = n9879 ^ x373;
  assign n9881 = n9139 ^ x374;
  assign n9882 = n9880 & ~n9881;
  assign n9883 = n9848 & n9882;
  assign n9884 = n9881 ^ n9880;
  assign n9885 = n9809 & ~n9884;
  assign n9886 = ~n9809 & ~n9847;
  assign n9887 = ~n9882 & n9886;
  assign n9888 = ~n9885 & ~n9887;
  assign n9889 = ~n9883 & n9888;
  assign n9890 = n9808 & n9889;
  assign n9891 = ~n9806 & ~n9807;
  assign n9892 = n9880 & n9881;
  assign n9893 = n9809 & n9892;
  assign n9894 = n9809 & n9847;
  assign n9895 = ~n9886 & ~n9894;
  assign n9896 = n9881 & ~n9895;
  assign n9897 = ~n9893 & ~n9896;
  assign n9898 = n9894 ^ n9809;
  assign n9899 = n9898 ^ n9894;
  assign n9900 = n9894 ^ n9881;
  assign n9901 = n9900 ^ n9894;
  assign n9902 = ~n9899 & ~n9901;
  assign n9903 = n9902 ^ n9894;
  assign n9904 = ~n9880 & n9903;
  assign n9905 = n9904 ^ n9894;
  assign n9906 = n9897 & ~n9905;
  assign n9907 = n9891 & ~n9906;
  assign n9908 = ~n9890 & ~n9907;
  assign n9909 = ~n9880 & n9881;
  assign n9910 = ~n9847 & n9909;
  assign n9911 = n9809 & n9910;
  assign n9912 = n9886 & ~n9909;
  assign n9913 = ~n9880 & ~n9881;
  assign n9914 = n9894 & n9913;
  assign n9915 = n9848 & n9881;
  assign n9916 = n9847 & n9892;
  assign n9917 = ~n9915 & ~n9916;
  assign n9918 = ~n9914 & n9917;
  assign n9919 = ~n9912 & n9918;
  assign n9920 = ~n9911 & n9919;
  assign n9921 = n9920 ^ n9806;
  assign n9922 = n9921 ^ n9920;
  assign n9923 = n9881 ^ n9809;
  assign n9924 = n9881 ^ n9847;
  assign n9925 = n9924 ^ n9847;
  assign n9926 = n9880 ^ n9809;
  assign n9927 = n9926 ^ n9847;
  assign n9928 = n9927 ^ n9847;
  assign n9929 = n9928 ^ n9847;
  assign n9930 = ~n9925 & n9929;
  assign n9931 = n9930 ^ n9847;
  assign n9932 = n9923 & n9931;
  assign n9933 = n9932 ^ n9927;
  assign n9934 = n9933 ^ n9920;
  assign n9935 = ~n9922 & n9934;
  assign n9936 = n9935 ^ n9920;
  assign n9937 = n9807 & ~n9936;
  assign n9938 = n9908 & ~n9937;
  assign n9939 = n9938 ^ n6893;
  assign n9940 = n9939 ^ x428;
  assign n9941 = n8699 & n8715;
  assign n9942 = n8691 & ~n8729;
  assign n9943 = ~n9941 & ~n9942;
  assign n9944 = n8718 & n8732;
  assign n9945 = n8688 & ~n9944;
  assign n9946 = ~n8706 & ~n8736;
  assign n9947 = ~n8738 & n9946;
  assign n9948 = n8695 & ~n9947;
  assign n9949 = ~n9945 & ~n9948;
  assign n9950 = n8686 & ~n8727;
  assign n9951 = n8558 & n8699;
  assign n9952 = n8739 & ~n9951;
  assign n9953 = ~n8720 & n9952;
  assign n9954 = ~n8701 & n9953;
  assign n9955 = n8687 & ~n9954;
  assign n9956 = ~n9950 & ~n9955;
  assign n9957 = n9949 & n9956;
  assign n9958 = n9943 & n9957;
  assign n9959 = n8710 & n9958;
  assign n9960 = n8698 ^ n8687;
  assign n9961 = n9960 ^ n8698;
  assign n9962 = n8698 ^ n8693;
  assign n9963 = n9961 & n9962;
  assign n9964 = n9963 ^ n8698;
  assign n9965 = ~n8686 & n9964;
  assign n9966 = n9959 & ~n9965;
  assign n9967 = ~n8696 & n9966;
  assign n9968 = ~n8689 & n9967;
  assign n9969 = n9968 ^ n7062;
  assign n9970 = n9969 ^ x426;
  assign n9971 = n9940 & n9970;
  assign n9972 = ~n9454 & ~n9466;
  assign n9973 = n9476 & ~n9972;
  assign n9974 = n9444 & ~n9489;
  assign n9975 = ~n9973 & ~n9974;
  assign n9976 = n9442 & n9462;
  assign n9977 = n9439 & n9464;
  assign n9978 = ~n9478 & ~n9482;
  assign n9979 = n9358 & ~n9978;
  assign n9980 = ~n9977 & ~n9979;
  assign n9981 = ~n9976 & n9980;
  assign n9982 = n9442 & n9465;
  assign n9983 = n9358 & n9436;
  assign n9984 = ~n9982 & ~n9983;
  assign n9985 = ~n9449 & ~n9464;
  assign n9988 = ~n9467 & ~n9483;
  assign n9986 = n9469 & n9489;
  assign n9987 = ~n9462 & n9986;
  assign n9989 = n9988 ^ n9987;
  assign n9990 = n9989 ^ n9988;
  assign n9991 = n9988 ^ n9357;
  assign n9992 = n9991 ^ n9988;
  assign n9993 = ~n9990 & n9992;
  assign n9994 = n9993 ^ n9988;
  assign n9995 = ~n9356 & ~n9994;
  assign n9996 = n9995 ^ n9988;
  assign n9997 = ~n9985 & n9996;
  assign n9998 = n9984 & n9997;
  assign n9999 = n9981 & n9998;
  assign n10000 = n9452 ^ n9356;
  assign n10001 = n10000 ^ n9452;
  assign n10002 = n9474 ^ n9452;
  assign n10003 = ~n10001 & n10002;
  assign n10004 = n10003 ^ n9452;
  assign n10005 = ~n9357 & n10004;
  assign n10006 = n9999 & ~n10005;
  assign n10007 = n9458 & n10006;
  assign n10008 = n9975 & n10007;
  assign n10009 = n10008 ^ n7027;
  assign n10010 = n10009 ^ x427;
  assign n10011 = n8458 ^ x425;
  assign n10012 = n10010 & ~n10011;
  assign n10013 = n9971 & n10012;
  assign n10014 = n9805 & n10013;
  assign n10015 = ~n9768 & n9804;
  assign n10016 = ~n9940 & ~n9970;
  assign n10017 = ~n10010 & n10011;
  assign n10018 = n10016 & n10017;
  assign n10019 = n9971 & n10017;
  assign n10020 = ~n10018 & ~n10019;
  assign n10021 = n10015 & ~n10020;
  assign n10022 = n9768 & ~n9804;
  assign n10023 = n10012 & n10016;
  assign n10024 = ~n10010 & ~n10011;
  assign n10025 = n9971 & n10024;
  assign n10026 = ~n10023 & ~n10025;
  assign n10027 = n10022 & ~n10026;
  assign n10028 = ~n10021 & ~n10027;
  assign n10029 = ~n9768 & ~n9804;
  assign n10030 = n9940 & ~n9970;
  assign n10031 = n10017 & n10030;
  assign n10032 = n10029 & n10031;
  assign n10033 = n10012 & n10030;
  assign n10034 = n10022 & n10033;
  assign n10035 = ~n10032 & ~n10034;
  assign n10036 = ~n9805 & ~n10029;
  assign n10037 = ~n9940 & n9970;
  assign n10038 = n10024 & n10037;
  assign n10039 = ~n10033 & ~n10038;
  assign n10040 = ~n10036 & ~n10039;
  assign n10041 = n10016 & n10024;
  assign n10042 = n9805 & n10041;
  assign n10043 = n10012 & n10037;
  assign n10044 = ~n9804 & n10043;
  assign n10045 = ~n10020 & n10022;
  assign n10046 = ~n10044 & ~n10045;
  assign n10047 = ~n9805 & ~n10022;
  assign n10048 = n10010 & n10011;
  assign n10049 = n10030 & n10048;
  assign n10050 = ~n10031 & ~n10049;
  assign n10051 = ~n10047 & ~n10050;
  assign n10052 = n10017 & n10037;
  assign n10053 = ~n10049 & ~n10052;
  assign n10054 = n10016 & n10048;
  assign n10055 = n9971 & n10048;
  assign n10056 = ~n10054 & ~n10055;
  assign n10057 = n10053 & n10056;
  assign n10058 = n10029 & ~n10057;
  assign n10059 = ~n10051 & ~n10058;
  assign n10060 = n10046 & n10059;
  assign n10061 = n9805 & n10055;
  assign n10062 = n10024 & n10030;
  assign n10063 = n10037 & n10048;
  assign n10064 = n9805 & n10063;
  assign n10065 = ~n10043 & ~n10064;
  assign n10066 = ~n10013 & n10065;
  assign n10067 = ~n10025 & n10066;
  assign n10068 = ~n10062 & n10067;
  assign n10069 = n10068 ^ n10015;
  assign n10070 = n10068 ^ n10064;
  assign n10071 = n10070 ^ n10064;
  assign n10072 = ~n10052 & ~n10054;
  assign n10073 = n10072 ^ n10064;
  assign n10074 = n10071 & n10073;
  assign n10075 = n10074 ^ n10064;
  assign n10076 = ~n10069 & n10075;
  assign n10077 = n10076 ^ n10015;
  assign n10078 = ~n10061 & ~n10077;
  assign n10079 = n10060 & n10078;
  assign n10080 = ~n10042 & n10079;
  assign n10081 = ~n10040 & n10080;
  assign n10082 = n10035 & n10081;
  assign n10083 = n10028 & n10082;
  assign n10084 = ~n10014 & n10083;
  assign n10085 = n10084 ^ n8304;
  assign n10086 = n10085 ^ x451;
  assign n10087 = n9939 ^ x430;
  assign n10088 = n9246 ^ n9107;
  assign n10089 = n10088 ^ n9246;
  assign n10090 = n9290 ^ n9246;
  assign n10091 = n10089 & ~n10090;
  assign n10092 = n10091 ^ n9246;
  assign n10093 = ~n9140 & n10092;
  assign n10094 = ~n9250 & ~n9281;
  assign n10095 = ~n9276 & n10094;
  assign n10096 = ~n9238 & ~n9260;
  assign n10097 = ~n9271 & n10096;
  assign n10098 = ~n10095 & ~n10097;
  assign n10099 = ~n9268 & ~n10098;
  assign n10100 = ~n9256 & n10099;
  assign n10101 = n10100 ^ n9140;
  assign n10102 = n10101 ^ n10100;
  assign n10103 = n9261 & ~n9278;
  assign n10104 = n9290 & n10103;
  assign n10105 = n10104 ^ n10100;
  assign n10106 = n10105 ^ n10100;
  assign n10107 = n10102 & ~n10106;
  assign n10108 = n10107 ^ n10100;
  assign n10109 = n9107 & ~n10108;
  assign n10110 = n10109 ^ n10100;
  assign n10111 = ~n10093 & n10110;
  assign n10112 = n9273 ^ n9107;
  assign n10113 = n10112 ^ n9273;
  assign n10114 = n9273 ^ n9243;
  assign n10115 = n10114 ^ n9273;
  assign n10116 = ~n10113 & n10115;
  assign n10117 = n10116 ^ n9273;
  assign n10118 = n9140 & ~n10117;
  assign n10119 = n10118 ^ n9273;
  assign n10120 = n10111 & n10119;
  assign n10121 = ~n9675 & n10120;
  assign n10122 = n9249 & n10121;
  assign n10123 = n9666 & n10122;
  assign n10124 = n9270 & n10123;
  assign n10125 = n10124 ^ n7835;
  assign n10126 = n10125 ^ x435;
  assign n10127 = n10087 & n10126;
  assign n10128 = n8856 & n8900;
  assign n10129 = n8854 & n8875;
  assign n10130 = n8883 & n8884;
  assign n10131 = ~n10129 & ~n10130;
  assign n10132 = ~n10128 & n10131;
  assign n10133 = n8856 & n8894;
  assign n10134 = n9631 & ~n10133;
  assign n10135 = ~n8902 & ~n9635;
  assign n10136 = ~n8866 & n10135;
  assign n10137 = n8883 & ~n10136;
  assign n10138 = ~n8854 & ~n8886;
  assign n10139 = ~n8879 & n10138;
  assign n10140 = n8856 & ~n10139;
  assign n10141 = ~n10137 & ~n10140;
  assign n10142 = n8872 & ~n8907;
  assign n10143 = n8895 & n9651;
  assign n10144 = n8780 & ~n10143;
  assign n10145 = ~n8878 & n8901;
  assign n10146 = n8875 & ~n10145;
  assign n10147 = ~n10144 & ~n10146;
  assign n10148 = ~n10142 & n10147;
  assign n10149 = n10141 & n10148;
  assign n10150 = n9633 & n10149;
  assign n10151 = n10134 & n10150;
  assign n10152 = n10132 & n10151;
  assign n10153 = ~n9625 & n10152;
  assign n10154 = n10153 ^ n7896;
  assign n10155 = n10154 ^ x434;
  assign n10156 = ~n8023 & n8034;
  assign n10157 = n7995 & ~n10156;
  assign n10158 = n8013 & ~n8026;
  assign n10159 = ~n7999 & n10158;
  assign n10160 = n8029 & ~n10159;
  assign n10161 = ~n10157 & ~n10160;
  assign n10162 = n9544 & n9552;
  assign n10163 = n8016 & ~n10162;
  assign n10164 = n8016 & n9549;
  assign n10165 = ~n8016 & ~n8029;
  assign n10166 = ~n8054 & ~n10165;
  assign n10167 = ~n10164 & ~n10166;
  assign n10168 = n9552 & n9562;
  assign n10169 = n7995 & ~n10168;
  assign n10170 = ~n8010 & n9560;
  assign n10171 = ~n8053 & n10170;
  assign n10172 = ~n8032 & n10171;
  assign n10173 = ~n8018 & n10172;
  assign n10174 = n7997 & ~n10173;
  assign n10175 = ~n10169 & ~n10174;
  assign n10176 = n10167 & n10175;
  assign n10177 = n9535 & n10176;
  assign n10178 = ~n10163 & n10177;
  assign n10179 = n10161 & n10178;
  assign n10180 = n8005 & n10179;
  assign n10181 = n10180 ^ n7868;
  assign n10182 = n10181 ^ x432;
  assign n10183 = ~n10155 & ~n10182;
  assign n10184 = n8211 & n8408;
  assign n10185 = n8381 & n8387;
  assign n10186 = ~n10184 & ~n10185;
  assign n10187 = n8337 & n8386;
  assign n10188 = n8389 & n10187;
  assign n10189 = ~n9515 & ~n10188;
  assign n10190 = n8409 & ~n8421;
  assign n10191 = n8389 & ~n10190;
  assign n10192 = n8419 & n9512;
  assign n10193 = n9506 & n10192;
  assign n10194 = n8385 & ~n10193;
  assign n10195 = ~n10191 & ~n10194;
  assign n10196 = n8211 & ~n9506;
  assign n10197 = n8393 & ~n8398;
  assign n10198 = ~n8405 & n10197;
  assign n10199 = ~n8425 & n10198;
  assign n10200 = n8381 & ~n10199;
  assign n10201 = ~n10196 & ~n10200;
  assign n10202 = n10195 & n10201;
  assign n10203 = n8412 & n10202;
  assign n10204 = n10189 & n10203;
  assign n10205 = n9514 & n10204;
  assign n10206 = n10186 & n10205;
  assign n10207 = ~n8456 & n10206;
  assign n10208 = n10207 ^ n7924;
  assign n10209 = n10208 ^ x433;
  assign n10210 = n9803 ^ x431;
  assign n10211 = n10209 & ~n10210;
  assign n10212 = n10183 & n10211;
  assign n10213 = n10155 & ~n10182;
  assign n10214 = ~n10209 & ~n10210;
  assign n10215 = n10213 & n10214;
  assign n10216 = ~n10212 & ~n10215;
  assign n10217 = n10127 & ~n10216;
  assign n10218 = ~n10087 & ~n10126;
  assign n10219 = n10215 & n10218;
  assign n10220 = n10087 & ~n10126;
  assign n10221 = n10155 & n10182;
  assign n10222 = n10211 & n10221;
  assign n10223 = ~n10155 & n10182;
  assign n10224 = n10214 & n10223;
  assign n10225 = ~n10222 & ~n10224;
  assign n10226 = n10220 & ~n10225;
  assign n10227 = ~n10219 & ~n10226;
  assign n10228 = n10211 & n10213;
  assign n10229 = n10220 & n10228;
  assign n10230 = n10211 & n10223;
  assign n10231 = n10218 & n10230;
  assign n10232 = ~n10229 & ~n10231;
  assign n10233 = ~n10209 & n10210;
  assign n10234 = n10183 & n10233;
  assign n10235 = ~n10126 & n10234;
  assign n10236 = n10214 & n10221;
  assign n10237 = ~n10087 & n10126;
  assign n10238 = ~n10220 & ~n10237;
  assign n10239 = n10236 & n10238;
  assign n10240 = n10183 & n10214;
  assign n10241 = n10127 & n10240;
  assign n10242 = n10209 & n10210;
  assign n10243 = n10221 & n10242;
  assign n10244 = n10183 & n10242;
  assign n10245 = ~n10243 & ~n10244;
  assign n10246 = n10220 & ~n10245;
  assign n10247 = ~n10241 & ~n10246;
  assign n10248 = n10223 & n10242;
  assign n10249 = ~n10234 & ~n10248;
  assign n10250 = ~n10212 & ~n10228;
  assign n10251 = n10225 & n10250;
  assign n10252 = n10249 & n10251;
  assign n10253 = n10237 & ~n10252;
  assign n10254 = n10223 & n10233;
  assign n10255 = n10213 & n10233;
  assign n10256 = ~n10254 & ~n10255;
  assign n10257 = n10256 ^ n10238;
  assign n10258 = n10257 ^ n10256;
  assign n10259 = n10213 & n10242;
  assign n10260 = n10221 & n10233;
  assign n10261 = ~n10244 & ~n10260;
  assign n10262 = ~n10254 & n10261;
  assign n10263 = ~n10218 & n10262;
  assign n10264 = ~n10248 & n10261;
  assign n10265 = ~n10127 & n10264;
  assign n10266 = ~n10263 & ~n10265;
  assign n10267 = ~n10259 & ~n10266;
  assign n10268 = n10267 ^ n10256;
  assign n10269 = n10258 & n10268;
  assign n10270 = n10269 ^ n10256;
  assign n10271 = ~n10253 & n10270;
  assign n10272 = n10247 & n10271;
  assign n10273 = ~n10239 & n10272;
  assign n10274 = ~n10235 & n10273;
  assign n10275 = n10232 & n10274;
  assign n10276 = n10227 & n10275;
  assign n10277 = ~n10217 & n10276;
  assign n10278 = n10277 ^ n8372;
  assign n10279 = n10278 ^ x452;
  assign n10280 = n10086 & ~n10279;
  assign n10281 = n9767 & n10280;
  assign n10282 = n8699 & n8701;
  assign n10283 = n8711 & ~n10282;
  assign n10284 = ~n8561 & ~n8706;
  assign n10285 = ~n8721 & n10284;
  assign n10286 = n8699 & ~n10285;
  assign n10287 = ~n8704 & n8739;
  assign n10288 = n8695 & ~n10287;
  assign n10289 = ~n10286 & ~n10288;
  assign n10290 = n8687 & ~n8718;
  assign n10291 = ~n8731 & n8737;
  assign n10292 = ~n8729 & ~n10291;
  assign n10293 = ~n10290 & ~n10292;
  assign n10294 = n10289 & n10293;
  assign n10295 = ~n8693 & ~n8726;
  assign n10296 = n10295 ^ n8686;
  assign n10297 = n10296 ^ n10295;
  assign n10298 = n10295 ^ n8698;
  assign n10299 = n10298 ^ n10295;
  assign n10300 = n10297 & n10299;
  assign n10301 = n10300 ^ n10295;
  assign n10302 = n8687 & ~n10301;
  assign n10303 = n10302 ^ n10295;
  assign n10304 = n10294 & n10303;
  assign n10305 = n8720 ^ n8687;
  assign n10306 = n10305 ^ n8720;
  assign n10307 = n8720 ^ n8562;
  assign n10308 = n10307 ^ n8720;
  assign n10309 = ~n10306 & ~n10308;
  assign n10310 = n10309 ^ n8720;
  assign n10311 = n8729 & n10310;
  assign n10312 = n10311 ^ n8720;
  assign n10313 = n10304 & ~n10312;
  assign n10314 = n10283 & n10313;
  assign n10315 = ~n8689 & n10314;
  assign n10316 = n10315 ^ n7193;
  assign n10317 = n10316 ^ x440;
  assign n10318 = n8998 & ~n9603;
  assign n10319 = ~n8999 & n10318;
  assign n10320 = n9011 & n10319;
  assign n10321 = ~n9013 & ~n9049;
  assign n10322 = n9025 & ~n10321;
  assign n10323 = ~n9008 & n9025;
  assign n10324 = ~n9032 & n9051;
  assign n10325 = n10324 ^ n8919;
  assign n10326 = n10325 ^ n10324;
  assign n10327 = n9055 & n9770;
  assign n10328 = n10327 ^ n10324;
  assign n10329 = ~n10326 & n10328;
  assign n10330 = n10329 ^ n10324;
  assign n10331 = n8920 & ~n10330;
  assign n10332 = ~n10323 & ~n10331;
  assign n10333 = ~n9021 & ~n9030;
  assign n10334 = ~n9585 & n10333;
  assign n10335 = n10334 ^ n9001;
  assign n10336 = n10335 ^ n9001;
  assign n10337 = n9001 ^ n8919;
  assign n10338 = n10337 ^ n9001;
  assign n10339 = ~n10336 & ~n10338;
  assign n10340 = n10339 ^ n9001;
  assign n10341 = ~n8920 & n10340;
  assign n10342 = n10341 ^ n9001;
  assign n10343 = n10332 & ~n10342;
  assign n10344 = n9590 & n10343;
  assign n10345 = n9772 & n10344;
  assign n10346 = ~n9017 & n10345;
  assign n10347 = ~n10322 & n10346;
  assign n10348 = ~n10320 & n10347;
  assign n10349 = n9581 & n10348;
  assign n10350 = n9010 & n10349;
  assign n10351 = n10350 ^ n8104;
  assign n10352 = n10351 ^ x439;
  assign n10353 = n10317 & n10352;
  assign n10354 = n10154 ^ x436;
  assign n10355 = n9449 & ~n9478;
  assign n10356 = n9442 & ~n10355;
  assign n10357 = n9464 & n9474;
  assign n10358 = ~n9436 & ~n9467;
  assign n10359 = n9476 & ~n10358;
  assign n10360 = ~n10357 & ~n10359;
  assign n10361 = n9358 & n9468;
  assign n10362 = ~n9436 & n9986;
  assign n10363 = n9444 & ~n10362;
  assign n10364 = ~n9466 & ~n9483;
  assign n10365 = ~n9446 & n10364;
  assign n10366 = n9358 & ~n10365;
  assign n10367 = n9484 & ~n9488;
  assign n10368 = n9442 & ~n10367;
  assign n10369 = n9449 & ~n9465;
  assign n10370 = ~n9454 & n10369;
  assign n10371 = n9476 & ~n10370;
  assign n10372 = ~n10368 & ~n10371;
  assign n10373 = ~n10366 & n10372;
  assign n10374 = ~n10363 & n10373;
  assign n10375 = ~n10361 & n10374;
  assign n10376 = n9981 & n10375;
  assign n10377 = n9461 & n10376;
  assign n10378 = n10360 & n10377;
  assign n10379 = ~n10356 & n10378;
  assign n10380 = ~n9441 & n10379;
  assign n10381 = n10380 ^ n7229;
  assign n10382 = n10381 ^ x441;
  assign n10383 = n10354 & n10382;
  assign n10384 = n9806 & n9807;
  assign n10385 = ~n9889 & n10384;
  assign n10386 = n9891 & ~n9933;
  assign n10387 = ~n10385 & ~n10386;
  assign n10388 = n9808 & ~n9920;
  assign n10389 = ~n9806 & n9807;
  assign n10390 = n9906 & n10389;
  assign n10391 = ~n10388 & ~n10390;
  assign n10392 = n10387 & n10391;
  assign n10393 = n10392 ^ n8076;
  assign n10394 = n10393 ^ x438;
  assign n10395 = n10125 ^ x437;
  assign n10396 = n10394 & ~n10395;
  assign n10397 = n10383 & n10396;
  assign n10398 = n10353 & n10397;
  assign n10399 = ~n10354 & n10382;
  assign n10400 = ~n10394 & ~n10395;
  assign n10401 = n10353 & n10400;
  assign n10402 = n10399 & n10401;
  assign n10403 = ~n10317 & ~n10352;
  assign n10404 = n10400 & n10403;
  assign n10405 = n10383 & n10404;
  assign n10406 = ~n10402 & ~n10405;
  assign n10407 = ~n10398 & n10406;
  assign n10408 = ~n10317 & n10352;
  assign n10409 = n10394 & n10395;
  assign n10410 = n10408 & n10409;
  assign n10411 = n10383 & n10410;
  assign n10412 = n10397 & n10403;
  assign n10413 = ~n10411 & ~n10412;
  assign n10414 = n10403 & n10409;
  assign n10415 = n10317 & ~n10352;
  assign n10416 = ~n10394 & n10395;
  assign n10417 = n10415 & n10416;
  assign n10418 = ~n10414 & ~n10417;
  assign n10419 = n10399 & ~n10418;
  assign n10420 = n10413 & ~n10419;
  assign n10421 = n10383 & n10417;
  assign n10422 = n10396 & n10408;
  assign n10423 = n10399 & n10422;
  assign n10424 = ~n10421 & ~n10423;
  assign n10425 = n10354 & ~n10382;
  assign n10426 = ~n10399 & ~n10425;
  assign n10427 = n10408 & n10416;
  assign n10428 = n10353 & n10409;
  assign n10429 = ~n10427 & ~n10428;
  assign n10430 = ~n10426 & ~n10429;
  assign n10431 = n10409 & n10415;
  assign n10432 = ~n10427 & ~n10431;
  assign n10433 = n10383 & ~n10432;
  assign n10434 = ~n10430 & ~n10433;
  assign n10435 = n10397 & n10415;
  assign n10436 = n10400 & n10415;
  assign n10437 = ~n10422 & ~n10436;
  assign n10438 = ~n10414 & ~n10431;
  assign n10439 = n10396 & n10415;
  assign n10440 = ~n10404 & ~n10439;
  assign n10441 = n10438 & n10440;
  assign n10442 = n10437 & n10441;
  assign n10443 = n10425 & ~n10442;
  assign n10444 = ~n10435 & ~n10443;
  assign n10445 = n10396 & n10403;
  assign n10446 = ~n10436 & ~n10445;
  assign n10447 = n10399 & ~n10446;
  assign n10448 = ~n10354 & ~n10382;
  assign n10449 = n10353 & n10396;
  assign n10450 = n10446 & ~n10449;
  assign n10451 = n10395 ^ n10352;
  assign n10452 = n10395 ^ n10317;
  assign n10453 = n10452 ^ n10317;
  assign n10454 = n10394 ^ n10317;
  assign n10455 = n10454 ^ n10317;
  assign n10456 = ~n10453 & n10455;
  assign n10457 = n10456 ^ n10317;
  assign n10458 = n10451 & n10457;
  assign n10459 = n10450 & ~n10458;
  assign n10460 = ~n10427 & n10459;
  assign n10461 = n10448 & n10460;
  assign n10462 = ~n10447 & ~n10461;
  assign n10463 = n10444 & n10462;
  assign n10464 = n10434 & n10463;
  assign n10465 = n10424 & n10464;
  assign n10466 = n10420 & n10465;
  assign n10467 = n10407 & n10466;
  assign n10468 = n10467 ^ n8172;
  assign n10469 = n10468 ^ x448;
  assign n10470 = n10316 ^ x442;
  assign n10471 = n9848 & n9909;
  assign n10472 = n9809 & n9882;
  assign n10473 = n9909 ^ n9886;
  assign n10474 = n10473 ^ n9886;
  assign n10475 = n9894 ^ n9886;
  assign n10476 = n10474 & n10475;
  assign n10477 = n10476 ^ n9886;
  assign n10478 = ~n10472 & ~n10477;
  assign n10479 = ~n10471 & n10478;
  assign n10480 = n9891 & ~n10479;
  assign n10481 = ~n9809 & n9892;
  assign n10482 = n9847 & n9913;
  assign n10483 = ~n9881 & n9895;
  assign n10484 = ~n10482 & ~n10483;
  assign n10485 = ~n10481 & n10484;
  assign n10486 = n9808 & ~n10485;
  assign n10487 = ~n10480 & ~n10486;
  assign n10488 = n9882 & n9894;
  assign n10489 = ~n9847 & ~n9884;
  assign n10490 = ~n9880 & n9895;
  assign n10491 = ~n10489 & ~n10490;
  assign n10492 = ~n10488 & n10491;
  assign n10493 = n10384 & ~n10492;
  assign n10494 = ~n9880 & n9894;
  assign n10495 = n9882 & n9895;
  assign n10496 = ~n10494 & ~n10495;
  assign n10497 = ~n9910 & n10496;
  assign n10498 = ~n9896 & n10497;
  assign n10499 = n10389 & ~n10498;
  assign n10500 = ~n10493 & ~n10499;
  assign n10501 = n10487 & n10500;
  assign n10502 = ~n9911 & n10501;
  assign n10503 = n10502 ^ n7163;
  assign n10504 = n10503 ^ x447;
  assign n10505 = n10470 & n10504;
  assign n10506 = n7999 & n8016;
  assign n10507 = ~n8007 & ~n9549;
  assign n10508 = ~n10165 & ~n10507;
  assign n10509 = ~n10506 & ~n10508;
  assign n10510 = ~n7682 & n8013;
  assign n10511 = n10510 ^ n8029;
  assign n10512 = n10510 ^ n7997;
  assign n10513 = n10512 ^ n7997;
  assign n10514 = ~n8002 & ~n8018;
  assign n10515 = n10514 ^ n7997;
  assign n10516 = n10513 & n10515;
  assign n10517 = n10516 ^ n7997;
  assign n10518 = ~n10511 & n10517;
  assign n10519 = n10518 ^ n8029;
  assign n10520 = n10509 & ~n10519;
  assign n10521 = n7997 & ~n8034;
  assign n10522 = n7995 & n8048;
  assign n10523 = ~n10521 & ~n10522;
  assign n10524 = n10520 & n10523;
  assign n10525 = ~n8004 & n10524;
  assign n10526 = ~n8021 & n10525;
  assign n10527 = n9539 & n10526;
  assign n10528 = n10527 ^ n7291;
  assign n10529 = n10528 ^ x446;
  assign n10530 = n10381 ^ x443;
  assign n10531 = n8859 & n8883;
  assign n10532 = n8780 & ~n9627;
  assign n10533 = ~n10531 & ~n10532;
  assign n10534 = n8872 & ~n9651;
  assign n10535 = n8887 & n8903;
  assign n10536 = ~n8900 & n10535;
  assign n10537 = n8875 & ~n10536;
  assign n10538 = ~n10534 & ~n10537;
  assign n10540 = n8895 & ~n8906;
  assign n10539 = ~n8899 & n9636;
  assign n10541 = n10540 ^ n10539;
  assign n10542 = n10541 ^ n10540;
  assign n10543 = n10540 ^ n8779;
  assign n10544 = n10543 ^ n10540;
  assign n10545 = ~n10542 & ~n10544;
  assign n10546 = n10545 ^ n10540;
  assign n10547 = ~n8778 & ~n10546;
  assign n10548 = n10547 ^ n10540;
  assign n10549 = n10538 & n10548;
  assign n10550 = n10533 & n10549;
  assign n10551 = n8868 & n10550;
  assign n10552 = n10134 & n10551;
  assign n10553 = n10132 & n10552;
  assign n10554 = ~n9625 & n10553;
  assign n10555 = n10554 ^ n7261;
  assign n10556 = n10555 ^ x444;
  assign n10557 = n10530 & n10556;
  assign n10558 = n8211 & ~n8434;
  assign n10559 = n8406 & ~n8408;
  assign n10560 = ~n8421 & n10559;
  assign n10561 = n8381 & ~n10560;
  assign n10562 = ~n10558 & ~n10561;
  assign n10563 = ~n8405 & n8426;
  assign n10564 = n8389 & ~n10563;
  assign n10565 = n9507 & n10197;
  assign n10566 = ~n8375 & n10565;
  assign n10567 = n8385 & ~n10566;
  assign n10568 = ~n10564 & ~n10567;
  assign n10569 = n10562 & n10568;
  assign n10570 = n8402 & n10569;
  assign n10571 = n9502 & n10570;
  assign n10572 = n10189 & n10571;
  assign n10573 = n10186 & n10572;
  assign n10574 = n8396 & n10573;
  assign n10575 = ~n8376 & n10574;
  assign n10576 = n10575 ^ n7328;
  assign n10577 = n10576 ^ x445;
  assign n10578 = n10557 & ~n10577;
  assign n10579 = ~n10529 & n10578;
  assign n10580 = n10505 & n10579;
  assign n10581 = n10556 & n10577;
  assign n10582 = n10530 & n10581;
  assign n10583 = ~n10529 & n10582;
  assign n10584 = n10505 & n10583;
  assign n10585 = n10470 & ~n10504;
  assign n10586 = ~n10529 & ~n10556;
  assign n10587 = n10530 & n10586;
  assign n10588 = ~n10577 & n10587;
  assign n10589 = n10585 & n10588;
  assign n10590 = ~n10470 & n10504;
  assign n10591 = n10529 & n10530;
  assign n10592 = n10581 & n10591;
  assign n10593 = ~n10579 & ~n10592;
  assign n10594 = n10590 & ~n10593;
  assign n10595 = ~n10589 & ~n10594;
  assign n10596 = n10556 & n10591;
  assign n10597 = ~n10577 & n10596;
  assign n10598 = n10585 & n10597;
  assign n10599 = ~n10530 & n10581;
  assign n10600 = n10529 & n10599;
  assign n10601 = n10600 ^ n10470;
  assign n10602 = n10601 ^ n10600;
  assign n10603 = ~n10556 & n10591;
  assign n10604 = n10577 & n10603;
  assign n10605 = n10604 ^ n10600;
  assign n10606 = n10605 ^ n10600;
  assign n10607 = n10602 & n10606;
  assign n10608 = n10607 ^ n10600;
  assign n10609 = n10504 & n10608;
  assign n10610 = n10609 ^ n10600;
  assign n10611 = ~n10598 & ~n10610;
  assign n10612 = n10504 ^ n10470;
  assign n10613 = n10597 & ~n10612;
  assign n10614 = n10583 & n10585;
  assign n10615 = ~n10470 & ~n10504;
  assign n10616 = n10577 & n10587;
  assign n10617 = ~n10592 & ~n10616;
  assign n10618 = ~n10579 & n10617;
  assign n10619 = n10615 & ~n10618;
  assign n10620 = ~n10530 & ~n10577;
  assign n10621 = ~n10556 & n10620;
  assign n10622 = ~n10530 & ~n10556;
  assign n10623 = n10577 & n10622;
  assign n10624 = n10529 & n10623;
  assign n10625 = n10556 & n10620;
  assign n10626 = ~n10529 & n10625;
  assign n10627 = ~n10624 & ~n10626;
  assign n10628 = ~n10621 & n10627;
  assign n10629 = n10505 & ~n10628;
  assign n10630 = ~n10619 & ~n10629;
  assign n10631 = ~n10577 & n10603;
  assign n10632 = ~n10616 & ~n10631;
  assign n10633 = n10586 & n10620;
  assign n10634 = n10529 & n10625;
  assign n10635 = ~n10599 & n10634;
  assign n10636 = n10635 ^ n10599;
  assign n10637 = ~n10633 & ~n10636;
  assign n10638 = n10632 & n10637;
  assign n10639 = n10590 & ~n10638;
  assign n10640 = ~n10530 & n10586;
  assign n10641 = n10577 & n10640;
  assign n10642 = ~n10633 & ~n10641;
  assign n10643 = n10585 & ~n10642;
  assign n10644 = ~n10624 & ~n10643;
  assign n10645 = ~n10504 & ~n10644;
  assign n10646 = ~n10639 & ~n10645;
  assign n10647 = n10630 & n10646;
  assign n10648 = ~n10614 & n10647;
  assign n10649 = ~n10613 & n10648;
  assign n10650 = n10631 ^ n10470;
  assign n10651 = n10650 ^ n10631;
  assign n10652 = n10529 & n10621;
  assign n10653 = ~n10626 & ~n10652;
  assign n10654 = n10653 ^ n10631;
  assign n10655 = ~n10651 & ~n10654;
  assign n10656 = n10655 ^ n10631;
  assign n10657 = ~n10504 & n10656;
  assign n10658 = n10649 & ~n10657;
  assign n10659 = n10611 & n10658;
  assign n10660 = n10595 & n10659;
  assign n10661 = ~n10584 & n10660;
  assign n10662 = ~n10580 & n10661;
  assign n10663 = n10662 ^ n8209;
  assign n10664 = n10663 ^ x453;
  assign n10665 = n10469 & ~n10664;
  assign n10666 = ~n9355 & ~n9766;
  assign n10667 = ~n10086 & n10279;
  assign n10668 = n10666 & n10667;
  assign n10669 = n10665 & n10668;
  assign n10670 = ~n10469 & ~n10664;
  assign n10671 = n10086 & n10279;
  assign n10672 = n10666 & n10671;
  assign n10673 = n10670 & n10672;
  assign n10674 = ~n10669 & ~n10673;
  assign n10675 = ~n10469 & n10664;
  assign n10676 = ~n9355 & n9766;
  assign n10677 = n10671 & n10676;
  assign n10678 = n10675 & n10677;
  assign n10679 = n10280 & n10676;
  assign n10680 = n10469 & n10679;
  assign n10681 = n10667 & n10676;
  assign n10682 = ~n10086 & ~n10279;
  assign n10683 = n10666 & n10682;
  assign n10684 = ~n10681 & ~n10683;
  assign n10685 = n10665 & ~n10684;
  assign n10686 = ~n10680 & ~n10685;
  assign n10687 = n9767 & n10667;
  assign n10688 = n9355 & ~n9766;
  assign n10689 = n10667 & n10688;
  assign n10690 = ~n10687 & ~n10689;
  assign n10691 = n10675 & ~n10690;
  assign n10692 = n10469 & n10664;
  assign n10693 = ~n10670 & ~n10692;
  assign n10694 = n10676 & n10682;
  assign n10695 = n10682 & n10688;
  assign n10696 = ~n10694 & ~n10695;
  assign n10697 = ~n10693 & ~n10696;
  assign n10698 = n9767 & n10671;
  assign n10699 = n10280 & n10688;
  assign n10700 = ~n10698 & ~n10699;
  assign n10701 = n9767 & n10682;
  assign n10702 = ~n10668 & ~n10701;
  assign n10703 = n10700 & n10702;
  assign n10704 = n10670 & ~n10703;
  assign n10705 = n10280 & n10666;
  assign n10706 = ~n10681 & ~n10705;
  assign n10707 = ~n10672 & ~n10683;
  assign n10708 = n10706 & n10707;
  assign n10709 = n10675 & ~n10708;
  assign n10710 = ~n10704 & ~n10709;
  assign n10711 = n10671 & n10688;
  assign n10712 = ~n10698 & ~n10711;
  assign n10713 = ~n10701 & n10712;
  assign n10714 = n10713 ^ n10664;
  assign n10715 = n10714 ^ n10713;
  assign n10716 = n10086 ^ n9355;
  assign n10717 = n10716 ^ n10279;
  assign n10718 = n10279 ^ n10086;
  assign n10719 = n10086 ^ n9766;
  assign n10720 = n10719 ^ n10086;
  assign n10721 = n10718 & n10720;
  assign n10722 = n10721 ^ n10086;
  assign n10723 = ~n10717 & n10722;
  assign n10724 = n10723 ^ n10713;
  assign n10725 = n10715 & ~n10724;
  assign n10726 = n10725 ^ n10713;
  assign n10727 = n10469 & ~n10726;
  assign n10728 = n10710 & ~n10727;
  assign n10729 = ~n10697 & n10728;
  assign n10730 = ~n10691 & n10729;
  assign n10731 = n10686 & n10730;
  assign n10732 = ~n10678 & n10731;
  assign n10733 = n10674 & n10732;
  assign n10734 = ~n10281 & n10733;
  assign n10735 = n10734 ^ n9531;
  assign n10736 = n10735 ^ x507;
  assign n10737 = ~n9073 & n9309;
  assign n10738 = ~n9308 & n9318;
  assign n10739 = ~n10737 & ~n10738;
  assign n10740 = n9330 ^ n8751;
  assign n10741 = ~n9073 & n9330;
  assign n10742 = ~n10740 & n10741;
  assign n10743 = n10742 ^ n10740;
  assign n10744 = n10739 & n10743;
  assign n10745 = n10744 ^ n8459;
  assign n10746 = n10745 ^ n10744;
  assign n10747 = ~n8751 & n9324;
  assign n10748 = ~n9315 & n9318;
  assign n10749 = ~n9345 & ~n10748;
  assign n10750 = ~n10747 & n10749;
  assign n10751 = n10750 ^ n10744;
  assign n10752 = ~n10746 & ~n10751;
  assign n10753 = n10752 ^ n10744;
  assign n10754 = n8066 & ~n10753;
  assign n10755 = n9308 ^ n9073;
  assign n10756 = n9073 ^ n8751;
  assign n10757 = n10756 ^ n8918;
  assign n10758 = n10757 ^ n8918;
  assign n10759 = n9331 & n10758;
  assign n10760 = n10759 ^ n8918;
  assign n10761 = n10755 & ~n10760;
  assign n10762 = n10761 ^ n10756;
  assign n10763 = n10762 ^ n8459;
  assign n10764 = n10763 ^ n10762;
  assign n10765 = n9330 ^ n9073;
  assign n10766 = n10765 ^ n9330;
  assign n10767 = n9341 ^ n9330;
  assign n10768 = ~n10766 & ~n10767;
  assign n10769 = n10768 ^ n9330;
  assign n10770 = ~n10747 & n10769;
  assign n10771 = n10770 ^ n10762;
  assign n10772 = n10764 & ~n10771;
  assign n10773 = n10772 ^ n10762;
  assign n10774 = ~n8066 & n10773;
  assign n10775 = ~n10754 & ~n10774;
  assign n10776 = n10775 ^ n9152;
  assign n10777 = n10776 ^ x478;
  assign n10778 = n10022 & n10041;
  assign n10779 = ~n10014 & ~n10778;
  assign n10780 = n10013 & n10022;
  assign n10781 = n9805 & n10038;
  assign n10782 = ~n10780 & ~n10781;
  assign n10783 = ~n10031 & ~n10063;
  assign n10784 = n10015 & ~n10783;
  assign n10785 = ~n10049 & ~n10054;
  assign n10786 = ~n10063 & n10785;
  assign n10787 = ~n10031 & n10786;
  assign n10788 = n10022 & ~n10787;
  assign n10789 = ~n10015 & ~n10064;
  assign n10790 = n10039 & n10066;
  assign n10791 = ~n10789 & ~n10790;
  assign n10792 = ~n10788 & ~n10791;
  assign n10793 = ~n10784 & n10792;
  assign n10794 = ~n10023 & ~n10062;
  assign n10795 = ~n10052 & ~n10055;
  assign n10796 = ~n10031 & n10795;
  assign n10797 = n10796 ^ n10785;
  assign n10798 = n9804 ^ n9768;
  assign n10799 = n10796 ^ n9804;
  assign n10800 = n10798 & ~n10799;
  assign n10801 = n10800 ^ n9804;
  assign n10802 = n10797 & ~n10801;
  assign n10803 = n10802 ^ n10785;
  assign n10804 = n10794 & n10803;
  assign n10805 = ~n10019 & n10804;
  assign n10806 = n10805 ^ n10029;
  assign n10807 = n10805 ^ n9805;
  assign n10808 = n10807 ^ n9805;
  assign n10809 = ~n10018 & ~n10033;
  assign n10810 = n10809 ^ n9805;
  assign n10811 = n10808 & n10810;
  assign n10812 = n10811 ^ n9805;
  assign n10813 = ~n10806 & n10812;
  assign n10814 = n10813 ^ n10029;
  assign n10815 = n10793 & ~n10814;
  assign n10816 = n10782 & n10815;
  assign n10817 = n10028 & n10816;
  assign n10818 = n10779 & n10817;
  assign n10819 = n10818 ^ n7130;
  assign n10820 = n10819 ^ x483;
  assign n10821 = ~n10777 & n10820;
  assign n10822 = n10528 ^ x400;
  assign n10823 = n9622 ^ x405;
  assign n10824 = ~n10822 & n10823;
  assign n10825 = n8686 & n8731;
  assign n10826 = n8733 & ~n8738;
  assign n10827 = ~n8561 & n10826;
  assign n10828 = n8707 & ~n10827;
  assign n10829 = ~n8558 & n9946;
  assign n10830 = n8699 & ~n10829;
  assign n10831 = n8740 & n10284;
  assign n10832 = n8688 & ~n10831;
  assign n10833 = ~n10830 & ~n10832;
  assign n10834 = ~n10828 & n10833;
  assign n10835 = ~n10825 & n10834;
  assign n10836 = n8726 ^ n8695;
  assign n10837 = ~n8720 & n8737;
  assign n10838 = n10837 ^ n8695;
  assign n10839 = n10838 ^ n10837;
  assign n10840 = n10837 ^ n8687;
  assign n10841 = ~n10839 & n10840;
  assign n10842 = n10841 ^ n10837;
  assign n10843 = n10836 & ~n10842;
  assign n10844 = n10843 ^ n8726;
  assign n10845 = n10835 & ~n10844;
  assign n10846 = ~n9965 & n10845;
  assign n10847 = ~n10312 & n10846;
  assign n10848 = n10283 & n10847;
  assign n10849 = n10848 ^ n8610;
  assign n10850 = n10849 ^ x402;
  assign n10851 = n9499 ^ x404;
  assign n10852 = n10850 & n10851;
  assign n10853 = n10503 ^ x401;
  assign n10854 = ~n9140 & ~n9686;
  assign n10855 = n9250 & ~n9273;
  assign n10856 = ~n10854 & ~n10855;
  assign n10857 = ~n9246 & ~n9280;
  assign n10858 = n9240 & ~n10857;
  assign n10859 = n9279 & ~n9289;
  assign n10860 = n9141 & ~n10859;
  assign n10861 = ~n10858 & ~n10860;
  assign n10862 = ~n9243 & ~n9260;
  assign n10863 = n9271 & ~n10862;
  assign n10864 = ~n9264 & n9679;
  assign n10865 = ~n9256 & n10864;
  assign n10866 = n9250 & ~n10865;
  assign n10867 = n9667 & n10094;
  assign n10868 = n9240 & ~n10867;
  assign n10869 = ~n9268 & n9279;
  assign n10870 = ~n9238 & n10869;
  assign n10871 = n9271 & ~n10870;
  assign n10872 = ~n9254 & n9282;
  assign n10873 = ~n9243 & n10872;
  assign n10874 = n9141 & ~n10873;
  assign n10875 = ~n10871 & ~n10874;
  assign n10876 = ~n10868 & n10875;
  assign n10877 = ~n10866 & n10876;
  assign n10878 = ~n10863 & n10877;
  assign n10879 = n10861 & n10878;
  assign n10880 = n10856 & n10879;
  assign n10881 = n9676 & n10880;
  assign n10882 = n10881 ^ n8582;
  assign n10883 = n10882 ^ x403;
  assign n10884 = n10853 & ~n10883;
  assign n10885 = n10852 & n10884;
  assign n10886 = n10824 & n10885;
  assign n10887 = ~n10822 & ~n10823;
  assign n10888 = n10850 & ~n10851;
  assign n10889 = n10884 & n10888;
  assign n10890 = n10887 & n10889;
  assign n10891 = ~n10850 & n10851;
  assign n10892 = ~n10853 & n10883;
  assign n10893 = n10891 & n10892;
  assign n10894 = n10852 & n10892;
  assign n10895 = ~n10893 & ~n10894;
  assign n10896 = n10887 & ~n10895;
  assign n10897 = n10824 & n10889;
  assign n10898 = n10822 & n10823;
  assign n10899 = ~n10850 & ~n10851;
  assign n10900 = n10892 & n10899;
  assign n10901 = ~n10853 & ~n10883;
  assign n10902 = n10852 & n10901;
  assign n10903 = ~n10900 & ~n10902;
  assign n10904 = n10898 & ~n10903;
  assign n10905 = ~n10897 & ~n10904;
  assign n10906 = n10891 & n10901;
  assign n10907 = n10888 & n10901;
  assign n10908 = ~n10906 & ~n10907;
  assign n10909 = n10822 & ~n10908;
  assign n10910 = n10822 & ~n10823;
  assign n10911 = n10853 & n10883;
  assign n10912 = n10852 & n10911;
  assign n10913 = n10899 & n10911;
  assign n10914 = ~n10912 & ~n10913;
  assign n10915 = n10888 & n10911;
  assign n10916 = n10884 & n10891;
  assign n10917 = ~n10915 & ~n10916;
  assign n10918 = n10914 & n10917;
  assign n10919 = n10910 & ~n10918;
  assign n10920 = ~n10909 & ~n10919;
  assign n10921 = n10899 & n10901;
  assign n10922 = n10888 & n10892;
  assign n10923 = ~n10893 & ~n10922;
  assign n10924 = ~n10894 & n10923;
  assign n10925 = ~n10921 & n10924;
  assign n10926 = n10824 & ~n10925;
  assign n10927 = n10824 & ~n10914;
  assign n10928 = n10891 & n10911;
  assign n10929 = ~n10915 & ~n10928;
  assign n10930 = ~n10900 & ~n10906;
  assign n10931 = n10929 & n10930;
  assign n10932 = ~n10885 & n10931;
  assign n10933 = n10887 & ~n10932;
  assign n10934 = ~n10927 & ~n10933;
  assign n10935 = ~n10893 & ~n10921;
  assign n10936 = n10910 & ~n10935;
  assign n10937 = n10884 & n10899;
  assign n10938 = ~n10885 & ~n10937;
  assign n10939 = ~n10912 & n10938;
  assign n10940 = ~n10922 & n10939;
  assign n10941 = n10898 & ~n10940;
  assign n10942 = ~n10936 & ~n10941;
  assign n10943 = n10934 & n10942;
  assign n10944 = ~n10926 & n10943;
  assign n10945 = n10920 & n10944;
  assign n10946 = n10905 & n10945;
  assign n10947 = ~n10896 & n10946;
  assign n10948 = ~n10890 & n10947;
  assign n10949 = ~n10886 & n10948;
  assign n10950 = n10949 ^ n9392;
  assign n10951 = n10950 ^ x481;
  assign n10952 = n10585 & ~n10617;
  assign n10953 = ~n10633 & ~n10634;
  assign n10954 = n10505 & ~n10953;
  assign n10955 = ~n10952 & ~n10954;
  assign n10956 = ~n10588 & ~n10597;
  assign n10957 = n10615 & ~n10956;
  assign n10958 = n10590 & ~n10627;
  assign n10959 = ~n10957 & ~n10958;
  assign n10960 = n10595 & n10959;
  assign n10961 = n10505 & n10641;
  assign n10962 = n10590 & n10597;
  assign n10963 = ~n10961 & ~n10962;
  assign n10964 = ~n10504 & n10641;
  assign n10965 = ~n10600 & ~n10616;
  assign n10966 = ~n10588 & n10965;
  assign n10967 = n10590 & ~n10966;
  assign n10968 = ~n10583 & ~n10604;
  assign n10969 = ~n10624 & n10968;
  assign n10970 = n10615 & ~n10969;
  assign n10971 = ~n10967 & ~n10970;
  assign n10972 = ~n10964 & n10971;
  assign n10973 = n10585 & n10636;
  assign n10974 = ~n10529 & n10599;
  assign n10975 = ~n10626 & ~n10631;
  assign n10976 = ~n10604 & n10975;
  assign n10977 = ~n10974 & n10976;
  assign n10978 = n10505 & ~n10977;
  assign n10979 = ~n10973 & ~n10978;
  assign n10980 = n10972 & n10979;
  assign n10981 = n10963 & n10980;
  assign n10982 = n10960 & n10981;
  assign n10983 = n10955 & n10982;
  assign n10984 = ~n10657 & n10983;
  assign n10985 = ~n10584 & n10984;
  assign n10986 = n10985 ^ n9106;
  assign n10987 = n10986 ^ x479;
  assign n10988 = n10951 & n10987;
  assign n10989 = n8750 ^ x417;
  assign n10990 = n9699 ^ x412;
  assign n10991 = ~n10989 & ~n10990;
  assign n10992 = n9476 & ~n9484;
  assign n10993 = ~n9467 & n9972;
  assign n10994 = ~n9464 & ~n10993;
  assign n10995 = ~n10992 & ~n10994;
  assign n10996 = ~n9468 & ~n9477;
  assign n10997 = n9444 & ~n10996;
  assign n10998 = ~n9446 & ~n9488;
  assign n10999 = n9358 & ~n10998;
  assign n11000 = ~n10997 & ~n10999;
  assign n11001 = ~n9439 & ~n9452;
  assign n11002 = n11001 ^ n9462;
  assign n11003 = n11002 ^ n9462;
  assign n11004 = n9462 ^ n9357;
  assign n11005 = n11004 ^ n9462;
  assign n11006 = ~n11003 & n11005;
  assign n11007 = n11006 ^ n9462;
  assign n11008 = ~n9464 & n11007;
  assign n11009 = n11008 ^ n9462;
  assign n11010 = n11000 & ~n11009;
  assign n11011 = n10995 & n11010;
  assign n11012 = n10360 & n11011;
  assign n11013 = ~n10005 & n11012;
  assign n11014 = ~n10356 & n11013;
  assign n11015 = n9975 & n11014;
  assign n11016 = ~n9441 & n11015;
  assign n11017 = n11016 ^ n7714;
  assign n11018 = n11017 ^ x415;
  assign n11019 = n8065 ^ x416;
  assign n11020 = n11018 & n11019;
  assign n11021 = n9895 & n9909;
  assign n11022 = n10478 & ~n11021;
  assign n11023 = n10389 & ~n11022;
  assign n11024 = ~n9911 & n10485;
  assign n11025 = n10384 & ~n11024;
  assign n11026 = ~n11023 & ~n11025;
  assign n11027 = n10492 ^ n9806;
  assign n11028 = n11027 ^ n10492;
  assign n11029 = n10498 ^ n10492;
  assign n11030 = ~n11028 & n11029;
  assign n11031 = n11030 ^ n10492;
  assign n11032 = ~n9807 & n11031;
  assign n11033 = n11026 & ~n11032;
  assign n11034 = n11033 ^ n7730;
  assign n11035 = n11034 ^ x414;
  assign n11036 = n9531 ^ x413;
  assign n11037 = ~n11035 & n11036;
  assign n11038 = n11020 & n11037;
  assign n11039 = n10991 & n11038;
  assign n11040 = n10989 & ~n10990;
  assign n11041 = ~n11018 & ~n11019;
  assign n11042 = n11035 & ~n11036;
  assign n11043 = n11041 & n11042;
  assign n11044 = n11040 & n11043;
  assign n11045 = ~n11039 & ~n11044;
  assign n11046 = n11035 & n11036;
  assign n11047 = n11020 & n11046;
  assign n11048 = n11040 & n11047;
  assign n11049 = n11018 & ~n11019;
  assign n11050 = n11037 & n11049;
  assign n11051 = n11040 & n11050;
  assign n11052 = ~n11048 & ~n11051;
  assign n11053 = n10989 & n10990;
  assign n11054 = ~n11035 & ~n11036;
  assign n11055 = n11041 & n11054;
  assign n11056 = n11020 & n11054;
  assign n11057 = ~n11055 & ~n11056;
  assign n11058 = n11053 & ~n11057;
  assign n11059 = n11052 & ~n11058;
  assign n11060 = n11046 & n11049;
  assign n11061 = ~n11038 & ~n11060;
  assign n11062 = n11053 & ~n11061;
  assign n11063 = ~n10991 & ~n11053;
  assign n11064 = n11020 & n11042;
  assign n11065 = ~n11043 & ~n11064;
  assign n11066 = ~n11063 & ~n11065;
  assign n11067 = ~n11062 & ~n11066;
  assign n11068 = ~n10989 & n10990;
  assign n11069 = ~n11018 & n11019;
  assign n11070 = n11037 & n11069;
  assign n11071 = ~n11050 & ~n11070;
  assign n11072 = n11041 & n11046;
  assign n11073 = ~n11047 & ~n11072;
  assign n11074 = n11071 & n11073;
  assign n11075 = n11068 & ~n11074;
  assign n11076 = n11054 & n11069;
  assign n11077 = n11049 & n11054;
  assign n11078 = ~n11076 & ~n11077;
  assign n11079 = n11037 & n11041;
  assign n11080 = n11042 & n11069;
  assign n11081 = ~n11079 & ~n11080;
  assign n11082 = n11078 & n11081;
  assign n11083 = n11040 & ~n11082;
  assign n11084 = ~n11075 & ~n11083;
  assign n11085 = n11042 & n11049;
  assign n11086 = n11063 & n11085;
  assign n11087 = ~n11064 & n11078;
  assign n11088 = n11068 & ~n11087;
  assign n11089 = ~n11060 & n11081;
  assign n11090 = ~n11076 & n11089;
  assign n11091 = n10991 & ~n11090;
  assign n11092 = ~n11088 & ~n11091;
  assign n11093 = ~n11086 & n11092;
  assign n11094 = n11084 & n11093;
  assign n11095 = n11067 & n11094;
  assign n11096 = n11059 & n11095;
  assign n11097 = n11045 & n11096;
  assign n11098 = n11046 & n11069;
  assign n11099 = n11098 ^ n11053;
  assign n11100 = n11098 ^ n10991;
  assign n11101 = n11100 ^ n10991;
  assign n11102 = n11079 ^ n10991;
  assign n11103 = ~n11101 & ~n11102;
  assign n11104 = n11103 ^ n10991;
  assign n11105 = n11099 & n11104;
  assign n11106 = n11105 ^ n11053;
  assign n11107 = n11097 & ~n11106;
  assign n11108 = n11107 ^ n7805;
  assign n11109 = n11108 ^ x482;
  assign n11110 = n10431 & n10448;
  assign n11111 = n10400 & n10408;
  assign n11112 = n10399 & n11111;
  assign n11113 = n10383 & ~n10437;
  assign n11114 = ~n11112 & ~n11113;
  assign n11115 = ~n11110 & n11114;
  assign n11116 = n10403 & n10416;
  assign n11117 = ~n10354 & n11116;
  assign n11118 = ~n10401 & n10446;
  assign n11119 = ~n11111 & n11118;
  assign n11120 = n10448 & ~n11119;
  assign n11121 = ~n11117 & ~n11120;
  assign n11122 = ~n10439 & ~n11111;
  assign n11123 = ~n10422 & n11122;
  assign n11124 = n11123 ^ n10399;
  assign n11125 = n11124 ^ n11123;
  assign n11126 = n10353 & n10416;
  assign n11127 = ~n10410 & ~n11126;
  assign n11128 = n11127 ^ n11123;
  assign n11129 = n11128 ^ n11123;
  assign n11130 = ~n11125 & ~n11129;
  assign n11131 = n11130 ^ n11123;
  assign n11132 = ~n10425 & ~n11131;
  assign n11133 = n11132 ^ n11123;
  assign n11134 = n11121 & n11133;
  assign n11135 = n10383 & ~n10438;
  assign n11136 = ~n10428 & ~n10431;
  assign n11137 = ~n10425 & n11136;
  assign n11138 = n10429 & ~n11116;
  assign n11139 = ~n10417 & n11138;
  assign n11140 = ~n10399 & n11139;
  assign n11141 = ~n11137 & ~n11140;
  assign n11142 = ~n10449 & ~n11141;
  assign n11143 = ~n10426 & ~n11142;
  assign n11144 = ~n11135 & ~n11143;
  assign n11145 = n11134 & n11144;
  assign n11146 = ~n10419 & n11145;
  assign n11147 = n11115 & n11146;
  assign n11148 = n10407 & n11147;
  assign n11149 = n11148 ^ n9433;
  assign n11150 = n11149 ^ x480;
  assign n11151 = n11109 & ~n11150;
  assign n11152 = n10988 & n11151;
  assign n11153 = n10821 & n11152;
  assign n11154 = ~n10951 & n10987;
  assign n11155 = n11150 & n11154;
  assign n11156 = ~n11109 & n11155;
  assign n11157 = ~n10777 & ~n10820;
  assign n11158 = n11156 & n11157;
  assign n11159 = n10777 & n10820;
  assign n11160 = n10951 & ~n10987;
  assign n11161 = n11151 & n11160;
  assign n11162 = n11159 & n11161;
  assign n11163 = ~n11158 & ~n11162;
  assign n11164 = n11151 & n11154;
  assign n11165 = n11157 & n11164;
  assign n11166 = ~n11109 & ~n11150;
  assign n11167 = n10988 & n11166;
  assign n11168 = n10821 & n11167;
  assign n11169 = ~n11165 & ~n11168;
  assign n11170 = n11109 & n11150;
  assign n11171 = n10988 & n11170;
  assign n11172 = ~n11167 & ~n11171;
  assign n11173 = n11157 & ~n11172;
  assign n11174 = n10777 & ~n10820;
  assign n11175 = n11109 & n11155;
  assign n11176 = ~n11109 & n11150;
  assign n11177 = n10988 & n11176;
  assign n11178 = ~n11152 & ~n11177;
  assign n11179 = ~n11175 & n11178;
  assign n11180 = ~n11167 & n11179;
  assign n11181 = n11174 & ~n11180;
  assign n11182 = n10987 ^ n10951;
  assign n11183 = n11182 ^ n11150;
  assign n11184 = n11150 ^ n11109;
  assign n11185 = n11109 ^ n10987;
  assign n11186 = n11185 ^ n11109;
  assign n11187 = n11184 & n11186;
  assign n11188 = n11187 ^ n11109;
  assign n11189 = n11183 & ~n11188;
  assign n11190 = n11189 ^ n10951;
  assign n11191 = n10821 & ~n11190;
  assign n11192 = n11154 & n11166;
  assign n11193 = ~n10951 & ~n10987;
  assign n11194 = n11176 & n11193;
  assign n11195 = n11160 & n11170;
  assign n11196 = ~n11194 & ~n11195;
  assign n11197 = ~n11161 & n11196;
  assign n11198 = ~n11174 & n11197;
  assign n11199 = n11160 & n11176;
  assign n11200 = n11170 & n11193;
  assign n11201 = n11151 & n11193;
  assign n11202 = ~n11200 & ~n11201;
  assign n11203 = ~n11199 & n11202;
  assign n11204 = ~n11157 & n11203;
  assign n11205 = ~n11198 & ~n11204;
  assign n11206 = ~n11192 & ~n11205;
  assign n11207 = n11206 ^ n10777;
  assign n11208 = n11207 ^ n11206;
  assign n11209 = ~n11156 & ~n11164;
  assign n11210 = n11160 & n11166;
  assign n11211 = ~n11195 & ~n11210;
  assign n11212 = ~n11192 & n11211;
  assign n11213 = n11209 & n11212;
  assign n11214 = ~n11177 & n11213;
  assign n11215 = ~n11194 & n11214;
  assign n11216 = n11215 ^ n11206;
  assign n11217 = n11216 ^ n11206;
  assign n11218 = n11208 & ~n11217;
  assign n11219 = n11218 ^ n11206;
  assign n11220 = n10820 & ~n11219;
  assign n11221 = n11220 ^ n11206;
  assign n11222 = ~n11191 & n11221;
  assign n11223 = ~n11181 & n11222;
  assign n11224 = ~n11173 & n11223;
  assign n11225 = n11169 & n11224;
  assign n11226 = n11163 & n11225;
  assign n11227 = ~n11153 & n11226;
  assign n11228 = n11227 ^ n9499;
  assign n11229 = n11228 ^ x502;
  assign n11230 = n10736 & ~n11229;
  assign n11231 = n10986 ^ x477;
  assign n11232 = ~n11047 & ~n11064;
  assign n11233 = n11053 & ~n11232;
  assign n11234 = ~n11056 & ~n11085;
  assign n11235 = n10991 & ~n11234;
  assign n11236 = ~n11233 & ~n11235;
  assign n11237 = ~n11061 & n11068;
  assign n11238 = ~n11043 & n11071;
  assign n11239 = ~n11063 & ~n11238;
  assign n11240 = ~n11055 & ~n11080;
  assign n11241 = n11078 & n11240;
  assign n11242 = n11068 & ~n11241;
  assign n11243 = n11036 ^ n11018;
  assign n11244 = n11035 ^ n11018;
  assign n11245 = n11244 ^ n11019;
  assign n11246 = n11245 ^ n11019;
  assign n11247 = n11246 ^ n11245;
  assign n11248 = n11245 ^ n11036;
  assign n11249 = ~n11247 & ~n11248;
  assign n11250 = n11249 ^ n11245;
  assign n11251 = n11243 & ~n11250;
  assign n11252 = n11251 ^ n11245;
  assign n11253 = n11040 & ~n11252;
  assign n11254 = ~n11242 & ~n11253;
  assign n11255 = ~n11051 & n11254;
  assign n11256 = ~n11239 & n11255;
  assign n11257 = ~n11237 & n11256;
  assign n11258 = n11236 & n11257;
  assign n11259 = ~n11039 & n11258;
  assign n11260 = n10990 ^ n10989;
  assign n11261 = n11076 ^ n10990;
  assign n11262 = n11261 ^ n11076;
  assign n11263 = n11076 ^ n11073;
  assign n11264 = n11262 & ~n11263;
  assign n11265 = n11264 ^ n11076;
  assign n11266 = n11260 & n11265;
  assign n11267 = n11259 & ~n11266;
  assign n11268 = ~n11106 & n11267;
  assign n11269 = n11064 ^ n10990;
  assign n11270 = n11269 ^ n11064;
  assign n11271 = n11077 ^ n11064;
  assign n11272 = n11270 & n11271;
  assign n11273 = n11272 ^ n11064;
  assign n11274 = ~n11260 & n11273;
  assign n11275 = n11268 & ~n11274;
  assign n11276 = n11275 ^ n9139;
  assign n11277 = n11276 ^ x472;
  assign n11278 = n11231 & n11277;
  assign n11279 = ~n10215 & ~n10224;
  assign n11280 = n10237 & ~n11279;
  assign n11281 = ~n10234 & ~n10259;
  assign n11282 = n10127 & ~n11281;
  assign n11283 = ~n10212 & ~n10222;
  assign n11284 = n10220 & ~n11283;
  assign n11285 = ~n11282 & ~n11284;
  assign n11286 = ~n11280 & n11285;
  assign n11287 = ~n10248 & ~n10260;
  assign n11288 = ~n10126 & ~n11287;
  assign n11289 = ~n10228 & ~n10240;
  assign n11290 = ~n10234 & n11289;
  assign n11291 = ~n10254 & n11290;
  assign n11292 = n10220 & ~n11291;
  assign n11293 = ~n11288 & ~n11292;
  assign n11294 = ~n10222 & ~n10230;
  assign n11295 = n10264 & n11294;
  assign n11296 = ~n10255 & n11295;
  assign n11297 = n10237 & ~n11296;
  assign n11298 = ~n10228 & ~n10255;
  assign n11299 = ~n10127 & n11298;
  assign n11300 = ~n10230 & ~n10236;
  assign n11301 = ~n10218 & n11300;
  assign n11302 = ~n11299 & ~n11301;
  assign n11303 = n11279 & ~n11302;
  assign n11304 = n11303 ^ n10245;
  assign n11305 = n11303 ^ n10238;
  assign n11306 = n11303 & n11305;
  assign n11307 = n11306 ^ n11303;
  assign n11308 = n11304 & n11307;
  assign n11309 = n11308 ^ n11306;
  assign n11310 = n11309 ^ n11303;
  assign n11311 = n11310 ^ n10238;
  assign n11312 = ~n11297 & n11311;
  assign n11313 = n11312 ^ n11297;
  assign n11314 = n11293 & ~n11313;
  assign n11315 = n11286 & n11314;
  assign n11316 = n11315 ^ n9235;
  assign n11317 = n11316 ^ x475;
  assign n11318 = n10824 & n10894;
  assign n11319 = n10906 & n10910;
  assign n11320 = ~n11318 & ~n11319;
  assign n11321 = n10822 & ~n10923;
  assign n11322 = n10888 ^ n10884;
  assign n11323 = n10887 & n11322;
  assign n11324 = ~n11321 & ~n11323;
  assign n11325 = n10894 & n10910;
  assign n11326 = ~n10913 & ~n10916;
  assign n11327 = n11326 ^ n10914;
  assign n11328 = n10823 ^ n10822;
  assign n11329 = n11328 ^ n10823;
  assign n11330 = n11326 ^ n10823;
  assign n11331 = ~n11329 & n11330;
  assign n11332 = n11331 ^ n10823;
  assign n11333 = n11327 & n11332;
  assign n11334 = n11333 ^ n10914;
  assign n11335 = ~n10885 & n11334;
  assign n11336 = ~n10889 & n11335;
  assign n11337 = n11336 ^ n10823;
  assign n11338 = n11337 ^ n11336;
  assign n11339 = ~n10902 & ~n10921;
  assign n11340 = ~n10912 & n11339;
  assign n11341 = n10929 & n11340;
  assign n11342 = ~n10937 & n11341;
  assign n11343 = n11342 ^ n11336;
  assign n11344 = n11343 ^ n11336;
  assign n11345 = n11338 & ~n11344;
  assign n11346 = n11345 ^ n11336;
  assign n11347 = ~n10822 & ~n11346;
  assign n11348 = n11347 ^ n11336;
  assign n11349 = ~n11325 & n11348;
  assign n11350 = n11324 & n11349;
  assign n11351 = n10905 & n11350;
  assign n11352 = ~n10896 & n11351;
  assign n11353 = n11320 & n11352;
  assign n11354 = n11353 ^ n9205;
  assign n11355 = n11354 ^ x473;
  assign n11356 = n11317 & ~n11355;
  assign n11357 = n10776 ^ x476;
  assign n11358 = n9719 & n9728;
  assign n11359 = n9725 ^ n9500;
  assign n11360 = n11359 ^ n9725;
  assign n11361 = n9725 ^ n9714;
  assign n11362 = n11360 & n11361;
  assign n11363 = n11362 ^ n9725;
  assign n11364 = n9532 & n11363;
  assign n11365 = ~n11358 & ~n11364;
  assign n11366 = n9728 & n9733;
  assign n11367 = ~n9730 & ~n9749;
  assign n11368 = n9704 & ~n11367;
  assign n11369 = ~n11366 & ~n11368;
  assign n11370 = n9738 & ~n9750;
  assign n11371 = n9533 & n9736;
  assign n11372 = ~n11370 & ~n11371;
  assign n11373 = ~n9707 & ~n9738;
  assign n11374 = n9716 & ~n11373;
  assign n11375 = ~n9725 & n11367;
  assign n11376 = ~n9733 & n11375;
  assign n11377 = n9533 & ~n11376;
  assign n11378 = n9744 & ~n9749;
  assign n11379 = ~n9714 & n11378;
  assign n11380 = n9716 & ~n11379;
  assign n11381 = n9701 & n9705;
  assign n11382 = ~n9736 & ~n11381;
  assign n11383 = n9704 & ~n11382;
  assign n11384 = n9624 & n9724;
  assign n11385 = ~n11381 & ~n11384;
  assign n11386 = ~n9714 & ~n9746;
  assign n11387 = n11385 & n11386;
  assign n11388 = n9728 & ~n11387;
  assign n11389 = ~n11383 & ~n11388;
  assign n11390 = ~n11380 & n11389;
  assign n11391 = ~n11377 & n11390;
  assign n11392 = ~n9727 & n11391;
  assign n11393 = ~n11374 & n11392;
  assign n11394 = n11372 & n11393;
  assign n11395 = n11369 & n11394;
  assign n11396 = n11365 & n11395;
  assign n11397 = ~n9729 & n11396;
  assign n11398 = n9712 & n11397;
  assign n11399 = n11398 ^ n9175;
  assign n11400 = n11399 ^ x474;
  assign n11401 = ~n11357 & n11400;
  assign n11402 = n11356 & n11401;
  assign n11403 = n11278 & n11402;
  assign n11404 = ~n11231 & n11277;
  assign n11405 = ~n11317 & n11355;
  assign n11406 = ~n11357 & ~n11400;
  assign n11407 = n11405 & n11406;
  assign n11408 = n11404 & n11407;
  assign n11409 = ~n11231 & ~n11277;
  assign n11410 = n11357 & n11400;
  assign n11411 = n11405 & n11410;
  assign n11412 = n11317 & n11355;
  assign n11413 = n11401 & n11412;
  assign n11414 = ~n11411 & ~n11413;
  assign n11415 = n11409 & ~n11414;
  assign n11416 = ~n11408 & ~n11415;
  assign n11417 = n11357 & ~n11400;
  assign n11418 = n11405 & n11417;
  assign n11419 = n11412 & n11417;
  assign n11420 = ~n11413 & ~n11419;
  assign n11421 = ~n11418 & n11420;
  assign n11422 = n11404 & ~n11421;
  assign n11423 = n11231 & ~n11277;
  assign n11424 = n11356 & n11406;
  assign n11425 = ~n11317 & ~n11355;
  assign n11426 = n11417 & n11425;
  assign n11427 = n11356 & n11410;
  assign n11428 = n11406 & n11425;
  assign n11429 = ~n11427 & ~n11428;
  assign n11430 = ~n11426 & n11429;
  assign n11431 = ~n11424 & n11430;
  assign n11432 = n11423 & ~n11431;
  assign n11433 = n11410 & n11412;
  assign n11434 = n11406 & n11412;
  assign n11435 = ~n11433 & ~n11434;
  assign n11436 = n11409 & ~n11435;
  assign n11437 = ~n11407 & ~n11434;
  assign n11438 = ~n11411 & n11437;
  assign n11439 = n11278 & ~n11438;
  assign n11440 = n11401 & n11405;
  assign n11441 = ~n11419 & n11435;
  assign n11442 = ~n11440 & n11441;
  assign n11443 = n11423 & ~n11442;
  assign n11444 = ~n11439 & ~n11443;
  assign n11445 = ~n11436 & n11444;
  assign n11446 = n11401 & n11425;
  assign n11447 = n11410 & n11425;
  assign n11448 = ~n11424 & ~n11447;
  assign n11449 = ~n11446 & n11448;
  assign n11450 = ~n11402 & n11449;
  assign n11451 = n11404 & ~n11450;
  assign n11452 = ~n11278 & ~n11409;
  assign n11453 = n11356 & n11417;
  assign n11454 = ~n11426 & ~n11446;
  assign n11455 = ~n11453 & n11454;
  assign n11456 = ~n11409 & n11455;
  assign n11457 = ~n11428 & n11456;
  assign n11458 = n11429 & ~n11446;
  assign n11459 = ~n11418 & n11458;
  assign n11460 = ~n11278 & n11459;
  assign n11461 = ~n11457 & ~n11460;
  assign n11462 = ~n11452 & n11461;
  assign n11463 = ~n11451 & ~n11462;
  assign n11464 = n11445 & n11463;
  assign n11465 = ~n11432 & n11464;
  assign n11466 = ~n11422 & n11465;
  assign n11467 = n11416 & n11466;
  assign n11468 = ~n11403 & n11467;
  assign n11469 = n11468 ^ n9699;
  assign n11470 = n11469 ^ x506;
  assign n11471 = n11108 ^ x484;
  assign n11472 = n10127 & n10222;
  assign n11473 = n10212 & n10218;
  assign n11474 = n10224 & n10238;
  assign n11475 = ~n11473 & ~n11474;
  assign n11476 = ~n10126 & n10236;
  assign n11477 = n10220 & n10240;
  assign n11478 = ~n11476 & ~n11477;
  assign n11479 = ~n10243 & n11287;
  assign n11480 = ~n10254 & n11479;
  assign n11481 = n10237 & ~n11480;
  assign n11482 = n10249 & n10261;
  assign n11483 = n10127 & ~n11482;
  assign n11484 = ~n10222 & n10245;
  assign n11485 = ~n10234 & n11484;
  assign n11486 = n10218 & ~n11485;
  assign n11487 = ~n11483 & ~n11486;
  assign n11488 = n10126 ^ n10087;
  assign n11491 = n10256 & ~n10259;
  assign n11492 = ~n10248 & n11491;
  assign n11489 = ~n10230 & n11289;
  assign n11490 = ~n10255 & n11489;
  assign n11493 = n11492 ^ n11490;
  assign n11494 = n11492 ^ n10126;
  assign n11495 = n11494 ^ n11492;
  assign n11496 = n11493 & n11495;
  assign n11497 = n11496 ^ n11492;
  assign n11498 = n11488 & ~n11497;
  assign n11499 = n11487 & ~n11498;
  assign n11500 = ~n11481 & n11499;
  assign n11501 = n11478 & n11500;
  assign n11502 = n11475 & n11501;
  assign n11503 = ~n11472 & n11502;
  assign n11504 = n10227 & n11503;
  assign n11505 = ~n10217 & n11504;
  assign n11506 = n11505 ^ n7993;
  assign n11507 = n11506 ^ x489;
  assign n11508 = n11471 & n11507;
  assign n11509 = n9343 & ~n10744;
  assign n11510 = n9314 & ~n10750;
  assign n11511 = ~n11509 & ~n11510;
  assign n11512 = n9329 & ~n10762;
  assign n11513 = n8460 & ~n10770;
  assign n11514 = ~n11512 & ~n11513;
  assign n11515 = n11511 & n11514;
  assign n11516 = n11515 ^ n6744;
  assign n11517 = n11516 ^ x486;
  assign n11518 = ~n9717 & ~n9733;
  assign n11519 = n9704 & ~n11518;
  assign n11520 = n9702 & n9728;
  assign n11521 = n9709 & n9716;
  assign n11522 = n9533 & ~n11385;
  assign n11523 = ~n11521 & ~n11522;
  assign n11524 = ~n11520 & n11523;
  assign n11525 = n9533 & n9733;
  assign n11526 = n9728 & n9736;
  assign n11527 = ~n11525 & ~n11526;
  assign n11528 = ~n9500 & n9707;
  assign n11529 = n9716 & ~n11367;
  assign n11530 = ~n11528 & ~n11529;
  assign n11531 = ~n9737 & ~n9746;
  assign n11532 = ~n9750 & ~n11531;
  assign n11533 = ~n9730 & n11385;
  assign n11534 = ~n9709 & n11533;
  assign n11535 = ~n9725 & n11534;
  assign n11536 = n9704 & ~n11535;
  assign n11537 = ~n11532 & ~n11536;
  assign n11538 = n11530 & n11537;
  assign n11539 = n11527 & n11538;
  assign n11540 = n11372 & n11539;
  assign n11541 = n11524 & n11540;
  assign n11542 = n11365 & n11541;
  assign n11543 = ~n11519 & n11542;
  assign n11544 = n9723 & n11543;
  assign n11545 = ~n9729 & n11544;
  assign n11546 = n11545 ^ n7679;
  assign n11547 = n11546 ^ x488;
  assign n11548 = ~n11517 & n11547;
  assign n11549 = n10505 & ~n10617;
  assign n11550 = n10585 & ~n10627;
  assign n11551 = ~n11549 & ~n11550;
  assign n11552 = n10632 & ~n10641;
  assign n11553 = n10615 & ~n11552;
  assign n11554 = n10953 & n10968;
  assign n11555 = n10590 & ~n11554;
  assign n11556 = ~n11553 & ~n11555;
  assign n11557 = n11551 & n11556;
  assign n11558 = n10652 ^ n10612;
  assign n11559 = n10652 ^ n10504;
  assign n11560 = n11559 ^ n10504;
  assign n11561 = n10974 ^ n10504;
  assign n11562 = ~n11560 & n11561;
  assign n11563 = n11562 ^ n10504;
  assign n11564 = ~n11558 & n11563;
  assign n11565 = n11564 ^ n10652;
  assign n11566 = n11557 & ~n11565;
  assign n11567 = n10611 & n11566;
  assign n11568 = n10960 & n11567;
  assign n11569 = n10955 & n11568;
  assign n11570 = ~n10580 & n11569;
  assign n11571 = n11570 ^ n7407;
  assign n11572 = n11571 ^ x487;
  assign n11573 = n10819 ^ x485;
  assign n11574 = n11572 & n11573;
  assign n11575 = n11548 & n11574;
  assign n11576 = n11508 & n11575;
  assign n11577 = ~n11471 & ~n11507;
  assign n11578 = n11517 & ~n11547;
  assign n11579 = ~n11572 & ~n11573;
  assign n11580 = n11578 & n11579;
  assign n11581 = n11548 & n11579;
  assign n11582 = ~n11580 & ~n11581;
  assign n11583 = n11577 & ~n11582;
  assign n11584 = ~n11576 & ~n11583;
  assign n11585 = ~n11572 & n11573;
  assign n11586 = n11548 & n11585;
  assign n11587 = n11508 & n11586;
  assign n11588 = n11574 & n11578;
  assign n11589 = n11471 & n11588;
  assign n11590 = ~n11517 & ~n11547;
  assign n11591 = n11585 & n11590;
  assign n11592 = ~n11471 & n11507;
  assign n11593 = n11471 & ~n11507;
  assign n11594 = ~n11592 & ~n11593;
  assign n11595 = n11591 & n11594;
  assign n11596 = ~n11589 & ~n11595;
  assign n11597 = n11517 & n11547;
  assign n11598 = n11572 & ~n11573;
  assign n11599 = n11597 & n11598;
  assign n11600 = n11577 & n11599;
  assign n11601 = n11574 & n11590;
  assign n11602 = n11592 & n11601;
  assign n11603 = ~n11580 & ~n11599;
  assign n11604 = n11508 & ~n11603;
  assign n11605 = n11574 & n11597;
  assign n11606 = ~n11601 & ~n11605;
  assign n11607 = n11578 & n11585;
  assign n11608 = ~n11575 & ~n11607;
  assign n11609 = n11606 & n11608;
  assign n11610 = n11577 & ~n11609;
  assign n11611 = n11590 & n11598;
  assign n11612 = ~n11581 & ~n11611;
  assign n11613 = n11508 & ~n11612;
  assign n11614 = ~n11610 & ~n11613;
  assign n11615 = n11579 & n11590;
  assign n11616 = n11548 & n11598;
  assign n11617 = n11585 & n11597;
  assign n11618 = ~n11586 & ~n11617;
  assign n11619 = n11578 & n11598;
  assign n11620 = n11579 & n11597;
  assign n11621 = ~n11611 & ~n11620;
  assign n11622 = ~n11619 & n11621;
  assign n11623 = n11618 & n11622;
  assign n11624 = ~n11616 & n11623;
  assign n11625 = ~n11615 & n11624;
  assign n11626 = ~n11594 & ~n11625;
  assign n11627 = n11614 & ~n11626;
  assign n11628 = ~n11604 & n11627;
  assign n11629 = ~n11602 & n11628;
  assign n11630 = ~n11600 & n11629;
  assign n11631 = n11596 & n11630;
  assign n11632 = ~n11587 & n11631;
  assign n11633 = n11584 & n11632;
  assign n11634 = n11633 ^ n9574;
  assign n11635 = n11634 ^ x505;
  assign n11636 = ~n11470 & ~n11635;
  assign n11637 = n9354 ^ x495;
  assign n11638 = n11546 ^ x490;
  assign n11639 = ~n11637 & ~n11638;
  assign n11640 = ~n10889 & n10929;
  assign n11641 = n10824 & ~n11640;
  assign n11642 = n10908 & ~n10937;
  assign n11643 = n10910 & ~n11642;
  assign n11644 = ~n11641 & ~n11643;
  assign n11645 = ~n10922 & n11339;
  assign n11646 = n10898 & ~n11645;
  assign n11647 = ~n10913 & n11640;
  assign n11648 = n10910 & ~n11647;
  assign n11649 = ~n10916 & ~n10937;
  assign n11650 = n10914 & n11649;
  assign n11651 = n10898 & ~n11650;
  assign n11652 = ~n11648 & ~n11651;
  assign n11653 = n10887 & ~n10939;
  assign n11654 = ~n10894 & n10930;
  assign n11655 = ~n10922 & n11654;
  assign n11656 = n10824 & ~n11655;
  assign n11657 = ~n11653 & ~n11656;
  assign n11658 = n11652 & n11657;
  assign n11659 = ~n10890 & n11658;
  assign n11660 = ~n11646 & n11659;
  assign n11661 = n10894 ^ n10823;
  assign n11662 = n11661 ^ n10894;
  assign n11663 = n10903 & n10923;
  assign n11664 = n11663 ^ n10894;
  assign n11665 = n11664 ^ n10894;
  assign n11666 = ~n11662 & ~n11665;
  assign n11667 = n11666 ^ n10894;
  assign n11668 = ~n10822 & n11667;
  assign n11669 = n11668 ^ n10894;
  assign n11670 = n11660 & ~n11669;
  assign n11671 = n11644 & n11670;
  assign n11672 = ~n10886 & n11671;
  assign n11673 = n11672 ^ n8958;
  assign n11674 = n11673 ^ x493;
  assign n11675 = n10991 & n11079;
  assign n11676 = ~n11057 & n11063;
  assign n11677 = ~n11675 & ~n11676;
  assign n11678 = n11047 & ~n11063;
  assign n11679 = ~n11080 & ~n11085;
  assign n11680 = n11053 & ~n11679;
  assign n11681 = ~n11678 & ~n11680;
  assign n11682 = ~n11070 & ~n11072;
  assign n11683 = ~n11077 & n11682;
  assign n11684 = n11063 & ~n11683;
  assign n11685 = ~n11038 & n11065;
  assign n11686 = n11068 & ~n11685;
  assign n11687 = ~n11684 & ~n11686;
  assign n11688 = n11040 & n11080;
  assign n11689 = n11071 & n11078;
  assign n11690 = n10991 & ~n11689;
  assign n11691 = ~n11688 & ~n11690;
  assign n11692 = n11687 & n11691;
  assign n11693 = n11681 & n11692;
  assign n11694 = n11677 & n11693;
  assign n11695 = n11059 & n11694;
  assign n11696 = ~n11106 & n11695;
  assign n11697 = ~n11274 & n11696;
  assign n11698 = n11697 ^ n8997;
  assign n11699 = n11698 ^ x492;
  assign n11700 = n10468 ^ x494;
  assign n11701 = ~n11699 & n11700;
  assign n11702 = n11506 ^ x491;
  assign n11703 = n11701 & ~n11702;
  assign n11704 = ~n11674 & n11703;
  assign n11705 = n11699 & ~n11702;
  assign n11706 = ~n11700 & n11705;
  assign n11707 = ~n11674 & n11706;
  assign n11708 = ~n11704 & ~n11707;
  assign n11709 = n11639 & ~n11708;
  assign n11710 = n11637 & ~n11638;
  assign n11711 = n11674 & n11700;
  assign n11712 = n11705 & n11711;
  assign n11713 = ~n11699 & ~n11700;
  assign n11714 = n11674 & n11702;
  assign n11715 = n11713 & n11714;
  assign n11716 = ~n11674 & n11702;
  assign n11717 = n11699 & n11716;
  assign n11718 = ~n11700 & n11717;
  assign n11719 = n11699 & n11714;
  assign n11720 = n11700 & n11719;
  assign n11721 = ~n11718 & ~n11720;
  assign n11722 = ~n11715 & n11721;
  assign n11723 = ~n11712 & n11722;
  assign n11724 = n11710 & ~n11723;
  assign n11725 = n11713 & n11716;
  assign n11726 = n11725 ^ n11638;
  assign n11727 = n11726 ^ n11725;
  assign n11728 = n11700 & n11717;
  assign n11729 = n11728 ^ n11725;
  assign n11730 = ~n11727 & n11729;
  assign n11731 = n11730 ^ n11725;
  assign n11732 = ~n11637 & n11731;
  assign n11733 = ~n11724 & ~n11732;
  assign n11734 = ~n11637 & n11638;
  assign n11735 = ~n11702 & n11713;
  assign n11736 = n11674 & n11735;
  assign n11737 = n11734 & n11736;
  assign n11738 = n11637 & n11638;
  assign n11739 = n11701 & n11714;
  assign n11740 = ~n11700 & n11719;
  assign n11741 = ~n11739 & ~n11740;
  assign n11742 = n11738 & ~n11741;
  assign n11743 = ~n11737 & ~n11742;
  assign n11744 = n11700 ^ n11674;
  assign n11745 = n11705 & n11744;
  assign n11746 = n11710 & n11745;
  assign n11747 = n11701 & n11716;
  assign n11748 = ~n11728 & ~n11747;
  assign n11749 = n11734 & ~n11748;
  assign n11750 = ~n11746 & ~n11749;
  assign n11751 = n11734 & n11740;
  assign n11752 = ~n11674 & n11735;
  assign n11753 = ~n11639 & n11752;
  assign n11754 = ~n11751 & ~n11753;
  assign n11755 = n11639 & ~n11722;
  assign n11756 = n11708 & ~n11718;
  assign n11757 = ~n11728 & n11756;
  assign n11758 = n11738 & ~n11757;
  assign n11759 = ~n11755 & ~n11758;
  assign n11760 = n11638 ^ n11637;
  assign n11761 = n11674 & n11703;
  assign n11762 = n11761 ^ n11638;
  assign n11763 = n11762 ^ n11761;
  assign n11764 = n11761 ^ n11747;
  assign n11765 = n11764 ^ n11761;
  assign n11766 = ~n11763 & n11765;
  assign n11767 = n11766 ^ n11761;
  assign n11768 = n11760 & n11767;
  assign n11769 = n11768 ^ n11761;
  assign n11770 = n11759 & ~n11769;
  assign n11771 = n11754 & n11770;
  assign n11772 = n11750 & n11771;
  assign n11773 = n11743 & n11772;
  assign n11774 = n11734 ^ n11712;
  assign n11775 = n11712 ^ n11639;
  assign n11776 = n11775 ^ n11639;
  assign n11777 = n11761 ^ n11639;
  assign n11778 = ~n11776 & ~n11777;
  assign n11779 = n11778 ^ n11639;
  assign n11780 = n11774 & n11779;
  assign n11781 = n11780 ^ n11734;
  assign n11782 = n11773 & ~n11781;
  assign n11783 = n11733 & n11782;
  assign n11784 = ~n11709 & n11783;
  assign n11785 = n11784 ^ n9622;
  assign n11786 = n11785 ^ x503;
  assign n11787 = ~n9312 & n9329;
  assign n11788 = ~n9318 & n9341;
  assign n11789 = ~n9308 & n9317;
  assign n11790 = ~n11788 & ~n11789;
  assign n11791 = ~n9073 & n9315;
  assign n11792 = ~n9344 & ~n11791;
  assign n11793 = n11790 & n11792;
  assign n11794 = n9314 & ~n11793;
  assign n11795 = ~n11787 & ~n11794;
  assign n11796 = n9326 & n9343;
  assign n11797 = n8460 & ~n9339;
  assign n11798 = ~n11796 & ~n11797;
  assign n11799 = n11795 & n11798;
  assign n11800 = n11799 ^ n8818;
  assign n11801 = n11800 ^ x462;
  assign n11802 = n10426 & n11116;
  assign n11803 = ~n10354 & ~n10437;
  assign n11804 = ~n11802 & ~n11803;
  assign n11805 = n10317 & n10396;
  assign n11806 = ~n10410 & ~n11805;
  assign n11807 = n10399 & ~n11806;
  assign n11808 = n10429 & n11122;
  assign n11809 = n10448 & ~n11808;
  assign n11810 = ~n11807 & ~n11809;
  assign n11811 = n11804 & n11810;
  assign n11812 = ~n10401 & n10432;
  assign n11813 = n11812 ^ n10382;
  assign n11814 = n11813 ^ n11812;
  assign n11815 = n11812 ^ n10460;
  assign n11816 = ~n11814 & ~n11815;
  assign n11817 = n11816 ^ n11812;
  assign n11818 = n10354 & ~n11817;
  assign n11819 = n11811 & ~n11818;
  assign n11820 = n10420 & n11819;
  assign n11821 = n11115 & n11820;
  assign n11822 = n11821 ^ n8804;
  assign n11823 = n11822 ^ x464;
  assign n11824 = ~n11801 & n11823;
  assign n11825 = n10218 & ~n10261;
  assign n11826 = n10249 & ~n10259;
  assign n11827 = ~n10238 & ~n11826;
  assign n11828 = ~n11825 & ~n11827;
  assign n11829 = n10243 ^ n10087;
  assign n11830 = n11829 ^ n10243;
  assign n11831 = n10255 ^ n10243;
  assign n11832 = n11831 ^ n10243;
  assign n11833 = n11830 & n11832;
  assign n11834 = n11833 ^ n10243;
  assign n11835 = n10126 & n11834;
  assign n11836 = n11835 ^ n10243;
  assign n11837 = n11828 & ~n11836;
  assign n11838 = n10220 & ~n11279;
  assign n11839 = ~n10260 & n11289;
  assign n11840 = n10237 & ~n11839;
  assign n11841 = ~n11838 & ~n11840;
  assign n11842 = ~n10218 & n11294;
  assign n11843 = n11300 & ~n11472;
  assign n11844 = n10250 & n11843;
  assign n11845 = ~n11842 & ~n11844;
  assign n11846 = n10238 & ~n11845;
  assign n11847 = ~n10254 & n11846;
  assign n11848 = n11847 ^ n10238;
  assign n11849 = n11841 & ~n11848;
  assign n11850 = n11837 & n11849;
  assign n11851 = n11286 & n11850;
  assign n11852 = ~n10217 & n11851;
  assign n11853 = n11852 ^ n8851;
  assign n11854 = n11853 ^ x463;
  assign n11855 = n10824 & n10916;
  assign n11856 = ~n10893 & n11642;
  assign n11857 = n10887 & ~n11856;
  assign n11858 = n10887 & ~n10914;
  assign n11859 = ~n10928 & n11340;
  assign n11860 = ~n10889 & n11859;
  assign n11861 = ~n10922 & n11860;
  assign n11862 = n10910 & ~n11861;
  assign n11863 = ~n11858 & ~n11862;
  assign n11864 = ~n10900 & n11339;
  assign n11865 = ~n10893 & n11864;
  assign n11866 = n10824 & ~n11865;
  assign n11868 = ~n10907 & n10924;
  assign n11867 = ~n10913 & n10938;
  assign n11869 = n11868 ^ n11867;
  assign n11870 = n11868 ^ n10898;
  assign n11871 = n11868 & n11870;
  assign n11872 = n11871 ^ n11868;
  assign n11873 = n11869 & n11872;
  assign n11874 = n11873 ^ n11871;
  assign n11875 = n11874 ^ n11868;
  assign n11876 = n11875 ^ n10898;
  assign n11877 = ~n11866 & n11876;
  assign n11878 = n11877 ^ n11866;
  assign n11879 = n11863 & ~n11878;
  assign n11880 = ~n10890 & n11879;
  assign n11881 = ~n10915 & n11880;
  assign n11882 = ~n11857 & n11881;
  assign n11883 = ~n11855 & n11882;
  assign n11884 = n11320 & n11883;
  assign n11885 = ~n10886 & n11884;
  assign n11886 = n11885 ^ n8685;
  assign n11887 = n11886 ^ x461;
  assign n11888 = n11854 & n11887;
  assign n11889 = n11824 & n11888;
  assign n11890 = n9739 ^ n9725;
  assign n11891 = n11890 ^ n9725;
  assign n11892 = n9725 ^ n9532;
  assign n11893 = n11892 ^ n9725;
  assign n11894 = ~n11891 & ~n11893;
  assign n11895 = n11894 ^ n9725;
  assign n11896 = n9750 & n11895;
  assign n11897 = n11896 ^ n9725;
  assign n11898 = n9719 ^ n9533;
  assign n11899 = n9719 ^ n9717;
  assign n11900 = n11899 ^ n9717;
  assign n11901 = n9717 ^ n9500;
  assign n11902 = n11900 & n11901;
  assign n11903 = n11902 ^ n9717;
  assign n11904 = n11898 & ~n11903;
  assign n11905 = n11904 ^ n9533;
  assign n11906 = ~n11897 & ~n11905;
  assign n11907 = n9728 & n11381;
  assign n11908 = ~n11384 & n11386;
  assign n11909 = n9716 & ~n11908;
  assign n11910 = ~n11907 & ~n11909;
  assign n11911 = n11906 & n11910;
  assign n11912 = n9732 & n11911;
  assign n11913 = ~n11374 & n11912;
  assign n11914 = n11527 & n11913;
  assign n11915 = ~n11364 & n11914;
  assign n11916 = n11524 & n11915;
  assign n11917 = n11369 & n11916;
  assign n11918 = ~n11519 & n11917;
  assign n11919 = n9712 & n11918;
  assign n11920 = n11919 ^ n8777;
  assign n11921 = n11920 ^ x465;
  assign n11922 = n10029 & n10063;
  assign n11923 = n10041 ^ n9804;
  assign n11924 = n11923 ^ n10041;
  assign n11925 = n10056 ^ n10041;
  assign n11926 = ~n11924 & ~n11925;
  assign n11927 = n11926 ^ n10041;
  assign n11928 = n10798 & n11927;
  assign n11929 = ~n11922 & ~n11928;
  assign n11930 = n10018 & n10022;
  assign n11931 = ~n10036 & ~n10053;
  assign n11932 = ~n11930 & ~n11931;
  assign n11933 = n10029 & n10055;
  assign n11934 = ~n10043 & ~n10062;
  assign n11935 = ~n10033 & n11934;
  assign n11936 = n10015 & ~n11935;
  assign n11937 = n9768 & n10031;
  assign n11938 = ~n10025 & n10039;
  assign n11939 = ~n10013 & n11938;
  assign n11940 = n10022 & ~n11939;
  assign n11941 = ~n11937 & ~n11940;
  assign n11942 = ~n10019 & n10786;
  assign n11943 = n10015 & ~n11942;
  assign n11944 = n10026 & ~n10041;
  assign n11945 = ~n10029 & n11944;
  assign n11946 = ~n10018 & ~n10043;
  assign n11947 = ~n10025 & n11946;
  assign n11948 = ~n9805 & n11947;
  assign n11949 = ~n11945 & ~n11948;
  assign n11950 = ~n10062 & ~n11949;
  assign n11951 = ~n10036 & ~n11950;
  assign n11952 = ~n11943 & ~n11951;
  assign n11953 = n11941 & n11952;
  assign n11954 = ~n11936 & n11953;
  assign n11955 = ~n11933 & n11954;
  assign n11956 = n11932 & n11955;
  assign n11957 = n11929 & n11956;
  assign n11958 = ~n10014 & n11957;
  assign n11959 = n11958 ^ n8555;
  assign n11960 = n11959 ^ x460;
  assign n11961 = ~n11921 & n11960;
  assign n11962 = n11889 & n11961;
  assign n11963 = ~n11854 & n11887;
  assign n11964 = n11824 & n11963;
  assign n11965 = n11921 & n11960;
  assign n11966 = n11964 & n11965;
  assign n11967 = ~n11962 & ~n11966;
  assign n11968 = n11801 & n11823;
  assign n11969 = n11888 & n11968;
  assign n11970 = n11960 ^ n11921;
  assign n11971 = n11969 & ~n11970;
  assign n11972 = n11801 & ~n11823;
  assign n11973 = n11963 & n11972;
  assign n11974 = ~n11921 & n11973;
  assign n11975 = ~n11854 & ~n11887;
  assign n11976 = n11972 & n11975;
  assign n11977 = n11854 & ~n11887;
  assign n11978 = n11968 & n11977;
  assign n11979 = ~n11976 & ~n11978;
  assign n11980 = n11824 & n11975;
  assign n11981 = ~n11801 & ~n11823;
  assign n11982 = n11977 & n11981;
  assign n11983 = ~n11980 & ~n11982;
  assign n11984 = n11979 & n11983;
  assign n11985 = n11961 & ~n11984;
  assign n11986 = n11823 ^ n11801;
  assign n11987 = n11963 & ~n11986;
  assign n11988 = n11921 & ~n11960;
  assign n11989 = n11987 & ~n11988;
  assign n11990 = ~n11985 & ~n11989;
  assign n11991 = n11887 ^ n11801;
  assign n11992 = n11991 ^ n11854;
  assign n11993 = n11992 ^ n11887;
  assign n11994 = ~n11823 & ~n11993;
  assign n11995 = n11994 ^ n11991;
  assign n11996 = n11988 & n11995;
  assign n11997 = n11972 & n11977;
  assign n11998 = ~n11980 & ~n11997;
  assign n11999 = n11824 & n11977;
  assign n12000 = n11982 ^ n11976;
  assign n12001 = ~n11921 & ~n11960;
  assign n12002 = n12001 ^ n11965;
  assign n12003 = n11982 ^ n11965;
  assign n12004 = n12003 ^ n11965;
  assign n12005 = ~n12002 & n12004;
  assign n12006 = n12005 ^ n11965;
  assign n12007 = n12000 & ~n12006;
  assign n12008 = n12007 ^ n11976;
  assign n12009 = ~n11999 & ~n12008;
  assign n12010 = n11998 & n12009;
  assign n12011 = ~n11970 & ~n12010;
  assign n12012 = ~n11996 & ~n12011;
  assign n12013 = n11990 & n12012;
  assign n12014 = ~n11974 & n12013;
  assign n12015 = ~n11971 & n12014;
  assign n12016 = n11967 & n12015;
  assign n12017 = n12016 ^ n9662;
  assign n12018 = n12017 ^ x504;
  assign n12019 = n11786 & ~n12018;
  assign n12020 = n11636 & n12019;
  assign n12021 = n11230 & n12020;
  assign n12022 = ~n11470 & n11635;
  assign n12023 = n11786 & n12018;
  assign n12024 = n12022 & n12023;
  assign n12025 = n11230 & n12024;
  assign n12026 = n10736 & n11229;
  assign n12027 = n11470 & ~n11635;
  assign n12028 = ~n11786 & ~n12018;
  assign n12029 = n12027 & n12028;
  assign n12030 = n12026 & n12029;
  assign n12031 = ~n12025 & ~n12030;
  assign n12032 = ~n12021 & n12031;
  assign n12033 = n11636 & n12028;
  assign n12034 = n12026 & n12033;
  assign n12035 = n11470 & n11635;
  assign n12036 = ~n11786 & n12018;
  assign n12037 = n12035 & n12036;
  assign n12038 = n12022 & n12028;
  assign n12039 = ~n12037 & ~n12038;
  assign n12040 = n11230 & ~n12039;
  assign n12041 = ~n12034 & ~n12040;
  assign n12042 = ~n10736 & n11229;
  assign n12043 = n11636 & n12023;
  assign n12044 = n12019 & n12027;
  assign n12045 = ~n12043 & ~n12044;
  assign n12046 = n12042 & ~n12045;
  assign n12047 = n12019 & n12035;
  assign n12048 = ~n12024 & ~n12047;
  assign n12049 = n12026 & ~n12048;
  assign n12050 = ~n12046 & ~n12049;
  assign n12051 = ~n12033 & n12039;
  assign n12052 = n12042 & ~n12051;
  assign n12053 = ~n10736 & ~n11229;
  assign n12054 = ~n12024 & ~n12044;
  assign n12055 = n12053 & ~n12054;
  assign n12056 = n12018 ^ n11635;
  assign n12057 = n11786 ^ n11470;
  assign n12058 = n12057 ^ n11470;
  assign n12059 = n12018 ^ n11470;
  assign n12060 = ~n12058 & n12059;
  assign n12061 = n12060 ^ n11470;
  assign n12062 = n12056 & n12061;
  assign n12063 = n11230 & n12062;
  assign n12064 = n11636 & n12036;
  assign n12065 = n12028 & n12035;
  assign n12066 = ~n12064 & ~n12065;
  assign n12067 = n12026 & ~n12066;
  assign n12068 = n11229 ^ n10736;
  assign n12069 = n12023 & n12027;
  assign n12070 = n12019 & n12022;
  assign n12071 = ~n12069 & ~n12070;
  assign n12072 = ~n12068 & ~n12071;
  assign n12073 = n12027 & n12036;
  assign n12074 = n12023 & n12035;
  assign n12075 = ~n12070 & ~n12074;
  assign n12076 = ~n12073 & n12075;
  assign n12077 = n12042 & ~n12076;
  assign n12078 = n12022 & n12036;
  assign n12079 = ~n12065 & ~n12078;
  assign n12080 = ~n12033 & n12079;
  assign n12081 = ~n12029 & n12080;
  assign n12082 = n12053 & ~n12081;
  assign n12083 = ~n12077 & ~n12082;
  assign n12084 = ~n12072 & n12083;
  assign n12085 = ~n12067 & n12084;
  assign n12086 = ~n12063 & n12085;
  assign n12087 = ~n12055 & n12086;
  assign n12088 = ~n12052 & n12087;
  assign n12089 = n12050 & n12088;
  assign n12090 = n12041 & n12089;
  assign n12091 = n12032 & n12090;
  assign n12092 = n12091 ^ n11920;
  assign n12093 = n12092 ^ x561;
  assign n12094 = n11982 & n12001;
  assign n12095 = n11975 & n11981;
  assign n12096 = ~n11999 & ~n12095;
  assign n12097 = ~n11970 & ~n12096;
  assign n12098 = ~n11973 & ~n11997;
  assign n12099 = n11965 & ~n12098;
  assign n12100 = n11888 & n11972;
  assign n12101 = n11963 & n11981;
  assign n12102 = n11888 & n11981;
  assign n12103 = ~n11969 & ~n12102;
  assign n12104 = ~n12101 & n12103;
  assign n12105 = ~n12100 & n12104;
  assign n12106 = n11988 & ~n12105;
  assign n12107 = ~n12099 & ~n12106;
  assign n12108 = n11968 & n11975;
  assign n12109 = ~n11976 & ~n12108;
  assign n12110 = n11998 & n12109;
  assign n12111 = n11961 & ~n12110;
  assign n12112 = n11978 & n12001;
  assign n12113 = ~n11889 & n12104;
  assign n12114 = n11961 & ~n12113;
  assign n12115 = n11983 & n12109;
  assign n12116 = n11988 & ~n12115;
  assign n12117 = ~n12114 & ~n12116;
  assign n12118 = ~n11889 & ~n12100;
  assign n12119 = n11963 & n11968;
  assign n12120 = ~n11964 & ~n12119;
  assign n12121 = n12118 & n12120;
  assign n12122 = n12121 ^ n11960;
  assign n12123 = n12122 ^ n12121;
  assign n12124 = ~n12100 & n12120;
  assign n12125 = ~n11969 & n12124;
  assign n12126 = n12125 ^ n12121;
  assign n12127 = ~n12123 & n12126;
  assign n12128 = n12127 ^ n12121;
  assign n12129 = ~n11970 & ~n12128;
  assign n12130 = n12117 & ~n12129;
  assign n12131 = ~n12112 & n12130;
  assign n12132 = ~n12111 & n12131;
  assign n12133 = n12107 & n12132;
  assign n12134 = ~n12097 & n12133;
  assign n12135 = ~n12094 & n12134;
  assign n12136 = n12135 ^ n8917;
  assign n12137 = n12136 ^ x520;
  assign n12138 = n11700 & n11705;
  assign n12139 = ~n11674 & n12138;
  assign n12140 = ~n11752 & ~n12139;
  assign n12141 = n11738 & ~n12140;
  assign n12142 = n11715 & n11734;
  assign n12143 = n11710 & n11728;
  assign n12144 = n11639 & ~n11741;
  assign n12145 = ~n12143 & ~n12144;
  assign n12146 = n11736 & ~n11760;
  assign n12147 = n11637 & n11707;
  assign n12148 = n11712 & n11734;
  assign n12149 = ~n11720 & ~n11745;
  assign n12150 = ~n11747 & n12149;
  assign n12151 = n11734 & ~n12150;
  assign n12154 = ~n11725 & ~n11761;
  assign n12152 = n11674 & n11706;
  assign n12153 = ~n11747 & ~n12152;
  assign n12155 = n12154 ^ n12153;
  assign n12156 = n12155 ^ n12154;
  assign n12157 = n12154 ^ n11637;
  assign n12158 = n12157 ^ n12154;
  assign n12159 = ~n12156 & n12158;
  assign n12160 = n12159 ^ n12154;
  assign n12161 = n11638 & ~n12160;
  assign n12162 = n12161 ^ n12154;
  assign n12163 = ~n12151 & n12162;
  assign n12164 = n11743 & n12163;
  assign n12165 = ~n12148 & n12164;
  assign n12166 = ~n12147 & n12165;
  assign n12167 = ~n12146 & n12166;
  assign n12168 = n12145 & n12167;
  assign n12169 = n11733 & n12168;
  assign n12170 = ~n12142 & n12169;
  assign n12171 = ~n12141 & n12170;
  assign n12172 = ~n11709 & n12171;
  assign n12173 = n12172 ^ n9803;
  assign n12174 = n12173 ^ x525;
  assign n12175 = n12137 & ~n12174;
  assign n12176 = n11822 ^ x466;
  assign n12177 = n11354 ^ x471;
  assign n12178 = ~n12176 & ~n12177;
  assign n12179 = n11920 ^ x467;
  assign n12180 = n10020 & n10026;
  assign n12181 = ~n10033 & n12180;
  assign n12182 = n9805 & ~n12181;
  assign n12183 = n10010 ^ n9970;
  assign n12184 = n12183 ^ n9940;
  assign n12185 = ~n10011 & n12184;
  assign n12186 = n10029 & n12185;
  assign n12187 = ~n12182 & ~n12186;
  assign n12188 = n10022 & ~n11947;
  assign n12189 = n10031 & ~n10036;
  assign n12190 = ~n9804 & ~n10053;
  assign n12191 = ~n12189 & ~n12190;
  assign n12192 = n10056 & n11947;
  assign n12193 = n10039 & n12192;
  assign n12194 = n10015 & ~n12193;
  assign n12195 = n12191 & ~n12194;
  assign n12196 = ~n12188 & n12195;
  assign n12197 = n12187 & n12196;
  assign n12198 = n11929 & n12197;
  assign n12199 = n10779 & n12198;
  assign n12200 = ~n10064 & n12199;
  assign n12201 = n12200 ^ n9846;
  assign n12202 = n12201 ^ x468;
  assign n12203 = n11276 ^ x470;
  assign n12205 = ~n12202 & ~n12203;
  assign n12204 = n12202 & ~n12203;
  assign n12206 = n12205 ^ n12204;
  assign n12207 = ~n12179 & n12206;
  assign n12208 = n12207 ^ n12205;
  assign n12209 = n10505 & n10624;
  assign n12210 = ~n10634 & n10653;
  assign n12211 = n10615 & ~n12210;
  assign n12212 = ~n12209 & ~n12211;
  assign n12213 = ~n10504 & n10974;
  assign n12214 = ~n10604 & n10617;
  assign n12215 = n10590 & ~n12214;
  assign n12216 = ~n10621 & n10632;
  assign n12217 = ~n10579 & n12216;
  assign n12218 = ~n10600 & n12217;
  assign n12219 = ~n10597 & n12218;
  assign n12220 = n10585 & ~n12219;
  assign n12221 = ~n10974 & n12210;
  assign n12222 = n10590 & ~n12221;
  assign n12223 = ~n10584 & n12214;
  assign n12224 = ~n10583 & ~n10592;
  assign n12225 = ~n10615 & n12224;
  assign n12226 = ~n12223 & ~n12225;
  assign n12227 = ~n10588 & ~n12226;
  assign n12228 = ~n10612 & ~n12227;
  assign n12229 = ~n12222 & ~n12228;
  assign n12230 = ~n12220 & n12229;
  assign n12231 = ~n10580 & n12230;
  assign n12232 = ~n12215 & n12231;
  assign n12233 = ~n12213 & n12232;
  assign n12234 = n12212 & n12233;
  assign n12235 = n10963 & n12234;
  assign n12236 = ~n10954 & n12235;
  assign n12237 = n12236 ^ n9879;
  assign n12238 = n12237 ^ x469;
  assign n12239 = n12238 ^ n12179;
  assign n12240 = n12202 & n12203;
  assign n12241 = n12240 ^ n12203;
  assign n12242 = n12238 ^ n12203;
  assign n12243 = n12242 ^ n12203;
  assign n12244 = ~n12241 & ~n12243;
  assign n12245 = n12244 ^ n12203;
  assign n12246 = n12239 & n12245;
  assign n12247 = ~n12208 & ~n12246;
  assign n12248 = n12178 & ~n12247;
  assign n12249 = n12176 & ~n12177;
  assign n12250 = n12179 & n12238;
  assign n12251 = n12204 & n12250;
  assign n12252 = ~n12202 & n12203;
  assign n12253 = ~n12179 & n12238;
  assign n12254 = n12252 & n12253;
  assign n12255 = ~n12179 & ~n12238;
  assign n12256 = n12205 & n12255;
  assign n12257 = ~n12254 & ~n12256;
  assign n12258 = n12179 & ~n12238;
  assign n12259 = n12203 & n12258;
  assign n12260 = n12240 ^ n12238;
  assign n12261 = n12260 ^ n12240;
  assign n12262 = n12240 ^ n12205;
  assign n12263 = n12261 & n12262;
  assign n12264 = n12263 ^ n12240;
  assign n12265 = ~n12259 & ~n12264;
  assign n12266 = n12257 & n12265;
  assign n12267 = ~n12251 & n12266;
  assign n12268 = n12249 & ~n12267;
  assign n12269 = ~n12248 & ~n12268;
  assign n12270 = n12176 & n12177;
  assign n12271 = n12203 ^ n12202;
  assign n12272 = n12271 ^ n12203;
  assign n12273 = n12202 ^ n12179;
  assign n12274 = n12273 ^ n12203;
  assign n12275 = n12274 ^ n12203;
  assign n12276 = n12275 ^ n12203;
  assign n12277 = ~n12272 & ~n12276;
  assign n12278 = n12277 ^ n12203;
  assign n12279 = ~n12238 & ~n12278;
  assign n12280 = n12279 ^ n12274;
  assign n12281 = n12270 & ~n12280;
  assign n12282 = ~n12176 & n12177;
  assign n12283 = n12202 & n12258;
  assign n12284 = n12252 & n12255;
  assign n12285 = ~n12179 & ~n12203;
  assign n12286 = ~n12205 & ~n12285;
  assign n12287 = ~n12240 & n12286;
  assign n12288 = n12238 & ~n12287;
  assign n12289 = ~n12284 & ~n12288;
  assign n12290 = ~n12283 & n12289;
  assign n12291 = n12282 & ~n12290;
  assign n12292 = ~n12281 & ~n12291;
  assign n12293 = n12269 & n12292;
  assign n12294 = n12293 ^ n9939;
  assign n12295 = n12294 ^ x524;
  assign n12296 = n11886 ^ x459;
  assign n12297 = n10278 ^ x454;
  assign n12298 = ~n12296 & ~n12297;
  assign n12299 = ~n11111 & n11127;
  assign n12300 = n10383 & ~n12299;
  assign n12301 = ~n10410 & ~n10458;
  assign n12302 = n10425 & ~n12301;
  assign n12303 = ~n12300 & ~n12302;
  assign n12304 = ~n10414 & ~n11126;
  assign n12305 = n10429 & n12304;
  assign n12306 = n12305 ^ n10382;
  assign n12307 = n12306 ^ n12305;
  assign n12308 = ~n10417 & n11812;
  assign n12309 = n12308 ^ n12305;
  assign n12310 = n12307 & n12309;
  assign n12311 = n12310 ^ n12305;
  assign n12312 = ~n10354 & ~n12311;
  assign n12313 = n10440 & ~n11111;
  assign n12314 = n12313 ^ n10426;
  assign n12315 = n12314 ^ n12313;
  assign n12316 = n10450 & ~n11116;
  assign n12317 = n12316 ^ n12313;
  assign n12318 = n12315 & n12317;
  assign n12319 = n12318 ^ n12313;
  assign n12320 = ~n12312 & n12319;
  assign n12321 = n12303 & n12320;
  assign n12322 = n10424 & n12321;
  assign n12323 = n12322 ^ n8533;
  assign n12324 = n12323 ^ x457;
  assign n12325 = n10663 ^ x455;
  assign n12326 = n12324 & ~n12325;
  assign n12327 = ~n11038 & ~n11098;
  assign n12328 = n11053 & ~n12327;
  assign n12329 = ~n11070 & n11679;
  assign n12330 = ~n11079 & n12329;
  assign n12331 = n11068 & ~n12330;
  assign n12332 = ~n12328 & ~n12331;
  assign n12333 = ~n11060 & ~n11098;
  assign n12334 = n11040 & ~n12333;
  assign n12335 = ~n11064 & n11240;
  assign n12336 = ~n10991 & n12335;
  assign n12337 = ~n11077 & n11679;
  assign n12338 = ~n11053 & n12337;
  assign n12339 = ~n12336 & ~n12338;
  assign n12340 = n11682 & ~n12339;
  assign n12341 = ~n11063 & ~n12340;
  assign n12342 = ~n12334 & ~n12341;
  assign n12343 = n12332 & n12342;
  assign n12344 = n11052 & n12343;
  assign n12345 = n11677 & n12344;
  assign n12346 = ~n11266 & n12345;
  assign n12347 = n11045 & n12346;
  assign n12348 = ~n11274 & n12347;
  assign n12349 = n12348 ^ n8496;
  assign n12350 = n12349 ^ x456;
  assign n12351 = n11959 ^ x458;
  assign n12352 = n12350 & n12351;
  assign n12353 = n12326 & n12352;
  assign n12354 = ~n12350 & ~n12351;
  assign n12355 = n12326 & n12354;
  assign n12356 = ~n12353 & ~n12355;
  assign n12357 = n12298 & ~n12356;
  assign n12358 = n12296 & ~n12297;
  assign n12359 = ~n12324 & n12325;
  assign n12360 = ~n12350 & n12351;
  assign n12361 = n12359 & n12360;
  assign n12362 = n12358 & n12361;
  assign n12363 = ~n12296 & n12297;
  assign n12364 = ~n12324 & ~n12325;
  assign n12365 = n12352 & n12364;
  assign n12366 = n12354 & n12364;
  assign n12367 = ~n12365 & ~n12366;
  assign n12368 = n12363 & ~n12367;
  assign n12369 = ~n12362 & ~n12368;
  assign n12370 = ~n12357 & n12369;
  assign n12371 = n12360 & n12364;
  assign n12372 = n12350 & ~n12351;
  assign n12373 = n12364 & n12372;
  assign n12374 = ~n12371 & ~n12373;
  assign n12375 = n12363 & ~n12374;
  assign n12376 = n12354 & n12359;
  assign n12377 = n12324 & n12325;
  assign n12378 = n12360 & n12377;
  assign n12379 = n12359 & n12372;
  assign n12380 = ~n12378 & ~n12379;
  assign n12381 = ~n12376 & n12380;
  assign n12382 = n12358 & ~n12381;
  assign n12383 = ~n12375 & ~n12382;
  assign n12384 = n12326 & n12360;
  assign n12385 = ~n12373 & ~n12384;
  assign n12386 = n12298 & ~n12385;
  assign n12387 = n12296 & n12297;
  assign n12388 = n12326 & n12372;
  assign n12389 = ~n12353 & ~n12388;
  assign n12390 = ~n12355 & ~n12371;
  assign n12391 = n12389 & n12390;
  assign n12392 = n12387 & ~n12391;
  assign n12393 = n12372 & n12377;
  assign n12394 = ~n12361 & ~n12393;
  assign n12395 = n12380 & n12394;
  assign n12396 = n12387 & ~n12395;
  assign n12397 = n12352 & n12377;
  assign n12398 = n12352 & n12359;
  assign n12399 = n12354 & n12377;
  assign n12400 = ~n12398 & ~n12399;
  assign n12401 = ~n12379 & n12400;
  assign n12402 = ~n12397 & n12401;
  assign n12403 = n12298 & ~n12402;
  assign n12404 = ~n12396 & ~n12403;
  assign n12405 = n12394 & ~n12399;
  assign n12406 = ~n12378 & n12405;
  assign n12407 = n12363 & ~n12406;
  assign n12408 = ~n12365 & n12389;
  assign n12409 = ~n12355 & n12408;
  assign n12410 = n12358 & ~n12409;
  assign n12411 = ~n12407 & ~n12410;
  assign n12412 = n12404 & n12411;
  assign n12413 = ~n12392 & n12412;
  assign n12414 = ~n12386 & n12413;
  assign n12415 = n12383 & n12414;
  assign n12416 = n12370 & n12415;
  assign n12417 = n12416 ^ n9969;
  assign n12418 = n12417 ^ x522;
  assign n12419 = ~n12295 & n12418;
  assign n12420 = n11161 & n11174;
  assign n12421 = ~n11175 & ~n11177;
  assign n12422 = n11159 & ~n12421;
  assign n12423 = ~n12420 & ~n12422;
  assign n12424 = n11166 & n11193;
  assign n12425 = ~n11195 & ~n12424;
  assign n12426 = n11157 & ~n12425;
  assign n12427 = n10821 & n11200;
  assign n12428 = ~n11194 & ~n11201;
  assign n12429 = ~n11195 & n12428;
  assign n12430 = ~n11167 & n12429;
  assign n12431 = ~n11164 & n12430;
  assign n12432 = n11159 & ~n12431;
  assign n12433 = ~n12427 & ~n12432;
  assign n12434 = n11199 ^ n11164;
  assign n12435 = n12434 ^ n11199;
  assign n12436 = n11199 ^ n10777;
  assign n12437 = n12436 ^ n11199;
  assign n12438 = n12435 & n12437;
  assign n12439 = n12438 ^ n11199;
  assign n12440 = ~n10820 & n12439;
  assign n12441 = n12440 ^ n11199;
  assign n12442 = n12433 & ~n12441;
  assign n12443 = ~n10821 & ~n11174;
  assign n12444 = ~n12428 & ~n12443;
  assign n12445 = n11172 & ~n11192;
  assign n12446 = ~n11192 & n12443;
  assign n12447 = ~n10821 & n11172;
  assign n12448 = ~n11157 & n12447;
  assign n12449 = ~n12446 & ~n12448;
  assign n12450 = ~n12445 & n12449;
  assign n12451 = n12421 & ~n12450;
  assign n12452 = n12451 ^ n11157;
  assign n12453 = ~n11161 & ~n11210;
  assign n12454 = n12453 ^ n12451;
  assign n12455 = n12454 ^ n12453;
  assign n12456 = ~n11174 & n12445;
  assign n12457 = ~n12443 & ~n12456;
  assign n12458 = n12457 ^ n12453;
  assign n12459 = ~n12455 & n12458;
  assign n12460 = n12459 ^ n12453;
  assign n12461 = ~n12452 & n12460;
  assign n12462 = n12461 ^ n11157;
  assign n12463 = ~n12444 & ~n12462;
  assign n12464 = n12442 & n12463;
  assign n12465 = ~n12426 & n12464;
  assign n12466 = ~n11158 & n12465;
  assign n12467 = n12423 & n12466;
  assign n12468 = ~n11153 & n12467;
  assign n12469 = n12468 ^ n10009;
  assign n12470 = n12469 ^ x523;
  assign n12471 = n10665 & n10677;
  assign n12472 = ~n10281 & ~n10711;
  assign n12473 = n10675 & ~n12472;
  assign n12474 = ~n12471 & ~n12473;
  assign n12475 = n10670 & n10677;
  assign n12476 = n10681 & n10692;
  assign n12477 = n10675 & n10701;
  assign n12478 = ~n12476 & ~n12477;
  assign n12479 = ~n12475 & n12478;
  assign n12480 = n10692 & n10705;
  assign n12481 = n10670 & n10694;
  assign n12482 = ~n12480 & ~n12481;
  assign n12483 = ~n10665 & n10693;
  assign n12484 = n10679 & ~n12483;
  assign n12485 = ~n10665 & ~n10701;
  assign n12486 = n10690 & n12485;
  assign n12487 = ~n10699 & n12486;
  assign n12488 = ~n10687 & n10700;
  assign n12489 = ~n10701 & n12488;
  assign n12490 = n10665 & ~n12489;
  assign n12491 = ~n10692 & ~n12490;
  assign n12492 = ~n12487 & ~n12491;
  assign n12494 = ~n10281 & n10690;
  assign n12493 = n10684 & ~n10695;
  assign n12495 = n12494 ^ n12493;
  assign n12496 = n12493 ^ n10670;
  assign n12497 = n12496 ^ n10670;
  assign n12498 = ~n10675 & ~n10695;
  assign n12499 = n12498 ^ n10670;
  assign n12500 = ~n12497 & n12499;
  assign n12501 = n12500 ^ n10670;
  assign n12502 = n12495 & ~n12501;
  assign n12503 = n12502 ^ n12494;
  assign n12504 = ~n10469 & ~n12503;
  assign n12505 = ~n12492 & ~n12504;
  assign n12506 = ~n10678 & n12505;
  assign n12507 = ~n12484 & n12506;
  assign n12508 = n12482 & n12507;
  assign n12509 = n10672 ^ n10664;
  assign n12510 = n12509 ^ n10672;
  assign n12511 = n10698 ^ n10672;
  assign n12512 = n12511 ^ n10672;
  assign n12513 = n12510 & n12512;
  assign n12514 = n12513 ^ n10672;
  assign n12515 = ~n10469 & n12514;
  assign n12516 = n12515 ^ n10672;
  assign n12517 = n12508 & ~n12516;
  assign n12518 = n12479 & n12517;
  assign n12519 = n12474 & n12518;
  assign n12520 = n10674 & n12519;
  assign n12521 = n12520 ^ n8458;
  assign n12522 = n12521 ^ x521;
  assign n12523 = ~n12470 & n12522;
  assign n12524 = n12419 & n12523;
  assign n12525 = n12175 & n12524;
  assign n12526 = n12137 & n12174;
  assign n12527 = ~n12470 & ~n12522;
  assign n12528 = n12419 & n12527;
  assign n12529 = n12526 & n12528;
  assign n12530 = ~n12137 & n12174;
  assign n12531 = n12295 & n12418;
  assign n12532 = n12527 & n12531;
  assign n12533 = n12530 & n12532;
  assign n12534 = n12295 & ~n12418;
  assign n12535 = n12470 & ~n12522;
  assign n12536 = n12534 & n12535;
  assign n12537 = n12175 & n12536;
  assign n12538 = ~n12533 & ~n12537;
  assign n12539 = ~n12529 & n12538;
  assign n12540 = ~n12525 & n12539;
  assign n12541 = n12530 & n12536;
  assign n12542 = ~n12137 & ~n12174;
  assign n12543 = n12532 & n12542;
  assign n12544 = ~n12541 & ~n12543;
  assign n12545 = ~n12295 & ~n12418;
  assign n12546 = n12470 & n12522;
  assign n12547 = n12545 & n12546;
  assign n12548 = n12542 & n12547;
  assign n12549 = n12535 & n12545;
  assign n12550 = n12530 & n12549;
  assign n12551 = ~n12548 & ~n12550;
  assign n12552 = n12534 & n12546;
  assign n12553 = n12552 ^ n12536;
  assign n12554 = n12553 ^ n12552;
  assign n12555 = n12552 ^ n12174;
  assign n12556 = n12555 ^ n12552;
  assign n12557 = n12554 & n12556;
  assign n12558 = n12557 ^ n12552;
  assign n12559 = n12137 & n12558;
  assign n12560 = n12559 ^ n12552;
  assign n12561 = n12551 & ~n12560;
  assign n12562 = n12531 & n12535;
  assign n12563 = ~n12137 & n12562;
  assign n12564 = n12523 & n12545;
  assign n12565 = n12523 & n12531;
  assign n12566 = n12527 & n12534;
  assign n12567 = n12419 & n12535;
  assign n12568 = ~n12566 & ~n12567;
  assign n12569 = ~n12565 & n12568;
  assign n12570 = ~n12564 & n12569;
  assign n12571 = n12542 & ~n12570;
  assign n12572 = ~n12563 & ~n12571;
  assign n12573 = n12523 & n12534;
  assign n12574 = n12419 & n12546;
  assign n12575 = ~n12573 & ~n12574;
  assign n12576 = ~n12565 & n12575;
  assign n12577 = ~n12528 & ~n12562;
  assign n12578 = ~n12547 & n12577;
  assign n12579 = n12576 & n12578;
  assign n12580 = n12175 & ~n12579;
  assign n12581 = n12527 & n12545;
  assign n12582 = n12575 & ~n12581;
  assign n12583 = n12530 & ~n12582;
  assign n12584 = n12531 & n12546;
  assign n12585 = ~n12524 & ~n12573;
  assign n12586 = ~n12564 & n12585;
  assign n12587 = ~n12566 & n12586;
  assign n12588 = ~n12549 & n12587;
  assign n12589 = ~n12584 & n12588;
  assign n12590 = n12526 & ~n12589;
  assign n12591 = ~n12583 & ~n12590;
  assign n12592 = ~n12580 & n12591;
  assign n12593 = n12572 & n12592;
  assign n12594 = n12561 & n12593;
  assign n12595 = n12544 & n12594;
  assign n12596 = n12540 & n12595;
  assign n12597 = n12596 ^ n11959;
  assign n12598 = n12597 ^ x556;
  assign n12599 = n12093 & ~n12598;
  assign n12600 = ~n11588 & ~n11617;
  assign n12601 = n11508 & ~n12600;
  assign n12602 = ~n11586 & ~n11607;
  assign n12603 = n11592 & ~n12602;
  assign n12604 = ~n12601 & ~n12603;
  assign n12605 = n11508 & n11601;
  assign n12606 = ~n11581 & ~n11619;
  assign n12607 = n11592 & ~n12606;
  assign n12608 = ~n12605 & ~n12607;
  assign n12609 = n11606 & ~n11617;
  assign n12610 = n11577 & ~n12609;
  assign n12611 = ~n11588 & ~n11599;
  assign n12612 = n11592 & ~n12611;
  assign n12613 = ~n12610 & ~n12612;
  assign n12614 = ~n11580 & ~n11616;
  assign n12615 = n11508 & ~n12614;
  assign n12616 = ~n11591 & n12606;
  assign n12617 = n11594 & ~n12616;
  assign n12618 = ~n12615 & ~n12617;
  assign n12619 = n12613 & n12618;
  assign n12620 = n11547 ^ n11517;
  assign n12621 = n12620 ^ n11573;
  assign n12622 = n12621 ^ n11572;
  assign n12623 = n12622 ^ n11547;
  assign n12624 = n12623 ^ n11573;
  assign n12625 = n11573 ^ n11547;
  assign n12626 = n11572 ^ n11547;
  assign n12627 = n12626 ^ n11547;
  assign n12628 = n12625 & ~n12627;
  assign n12629 = n12628 ^ n11547;
  assign n12630 = ~n12624 & n12629;
  assign n12631 = n12630 ^ n12621;
  assign n12632 = n12631 ^ n11621;
  assign n12633 = n12632 ^ n11621;
  assign n12634 = n11621 ^ n11507;
  assign n12635 = n12634 ^ n11621;
  assign n12636 = ~n12633 & ~n12635;
  assign n12637 = n12636 ^ n11621;
  assign n12638 = n11471 & ~n12637;
  assign n12639 = n12638 ^ n11621;
  assign n12640 = n12619 & n12639;
  assign n12641 = n12608 & n12640;
  assign n12642 = n12604 & n12641;
  assign n12643 = n12642 ^ n8065;
  assign n12644 = n12643 ^ x514;
  assign n12645 = n12521 ^ x519;
  assign n12646 = ~n12644 & ~n12645;
  assign n12647 = n11638 & n11718;
  assign n12648 = n11738 & n11740;
  assign n12649 = ~n12647 & ~n12648;
  assign n12650 = ~n11708 & n11710;
  assign n12651 = ~n11715 & ~n11739;
  assign n12652 = n11639 & ~n12651;
  assign n12653 = ~n11720 & ~n11725;
  assign n12654 = ~n11760 & ~n12653;
  assign n12655 = ~n11736 & ~n11761;
  assign n12656 = n11738 & ~n12655;
  assign n12657 = ~n12654 & ~n12656;
  assign n12658 = n11639 & n11745;
  assign n12659 = n11700 ^ n11699;
  assign n12660 = n11699 ^ n11674;
  assign n12661 = n12659 & ~n12660;
  assign n12662 = ~n11702 & n12661;
  assign n12663 = ~n11752 & ~n12662;
  assign n12664 = n11734 & ~n12663;
  assign n12665 = ~n11720 & ~n11728;
  assign n12666 = n12651 & n12665;
  assign n12667 = n11710 & ~n12666;
  assign n12668 = ~n12664 & ~n12667;
  assign n12669 = ~n12658 & n12668;
  assign n12670 = n12657 & n12669;
  assign n12671 = ~n12141 & n12670;
  assign n12672 = ~n11709 & n12671;
  assign n12673 = ~n12148 & n12672;
  assign n12674 = ~n12652 & n12673;
  assign n12675 = ~n12650 & n12674;
  assign n12676 = n12649 & n12675;
  assign n12677 = n11750 & n12676;
  assign n12678 = ~n12142 & n12677;
  assign n12679 = n12678 ^ n9072;
  assign n12680 = n12679 ^ x517;
  assign n12714 = n11407 & n11409;
  assign n12715 = ~n11427 & n11448;
  assign n12716 = n11423 & ~n12715;
  assign n12717 = ~n12714 & ~n12716;
  assign n12718 = ~n11427 & n11454;
  assign n12719 = ~n11418 & n12718;
  assign n12720 = n11404 & ~n12719;
  assign n12721 = n11421 & n11454;
  assign n12722 = n11423 & ~n12721;
  assign n12723 = ~n12720 & ~n12722;
  assign n12724 = ~n11428 & ~n11453;
  assign n12725 = ~n11447 & n12724;
  assign n12726 = ~n11402 & n12725;
  assign n12727 = n11409 & ~n12726;
  assign n12728 = ~n11446 & ~n11453;
  assign n12729 = ~n11424 & n12728;
  assign n12730 = ~n11418 & ~n11440;
  assign n12731 = ~n11433 & n12730;
  assign n12732 = ~n11407 & n12731;
  assign n12733 = n12729 & n12732;
  assign n12734 = n11278 & ~n12733;
  assign n12736 = n11414 & ~n11434;
  assign n12737 = ~n11419 & n12736;
  assign n12735 = ~n11411 & n11435;
  assign n12738 = n12737 ^ n12735;
  assign n12739 = n12737 ^ n11277;
  assign n12740 = n12739 ^ n12737;
  assign n12741 = n12738 & ~n12740;
  assign n12742 = n12741 ^ n12737;
  assign n12743 = ~n11231 & ~n12742;
  assign n12744 = ~n12734 & ~n12743;
  assign n12745 = ~n12727 & n12744;
  assign n12746 = n12723 & n12745;
  assign n12747 = n12717 & n12746;
  assign n12748 = ~n11403 & n12747;
  assign n12749 = n12748 ^ n9307;
  assign n12750 = n12749 ^ x516;
  assign n12681 = n12358 & ~n12367;
  assign n12682 = n12298 & ~n12400;
  assign n12683 = ~n12681 & ~n12682;
  assign n12684 = n12358 & n12397;
  assign n12685 = n12384 & n12387;
  assign n12686 = ~n12684 & ~n12685;
  assign n12687 = ~n12371 & n12394;
  assign n12688 = n12298 & ~n12687;
  assign n12689 = ~n12379 & ~n12399;
  assign n12690 = ~n12384 & n12689;
  assign n12691 = ~n12355 & n12690;
  assign n12692 = n12358 & ~n12691;
  assign n12693 = ~n12688 & ~n12692;
  assign n12694 = ~n12356 & n12363;
  assign n12695 = n12297 ^ n12296;
  assign n12696 = ~n12373 & n12389;
  assign n12697 = ~n12695 & ~n12696;
  assign n12698 = ~n12387 & ~n12393;
  assign n12699 = ~n12398 & n12698;
  assign n12700 = ~n12378 & n12699;
  assign n12701 = ~n12376 & n12700;
  assign n12702 = ~n12361 & n12401;
  assign n12703 = ~n12363 & n12702;
  assign n12704 = ~n12701 & ~n12703;
  assign n12705 = n12297 & n12704;
  assign n12706 = ~n12697 & ~n12705;
  assign n12707 = ~n12694 & n12706;
  assign n12708 = n12693 & n12707;
  assign n12709 = n12686 & n12708;
  assign n12710 = n12683 & n12709;
  assign n12711 = n12369 & n12710;
  assign n12712 = n12711 ^ n8750;
  assign n12713 = n12712 ^ x515;
  assign n12751 = n12750 ^ n12713;
  assign n12752 = n12751 ^ n12713;
  assign n12753 = n12136 ^ x518;
  assign n12754 = n12753 ^ n12750;
  assign n12755 = n12754 ^ n12713;
  assign n12756 = n12755 ^ n12713;
  assign n12757 = n12756 ^ n12713;
  assign n12758 = n12752 & n12757;
  assign n12759 = n12758 ^ n12713;
  assign n12760 = ~n12680 & n12759;
  assign n12761 = n12760 ^ n12755;
  assign n12762 = n12646 & ~n12761;
  assign n12763 = ~n12644 & n12645;
  assign n12764 = ~n12680 & n12753;
  assign n12765 = ~n12713 & n12750;
  assign n12766 = n12764 & n12765;
  assign n12767 = ~n12713 & ~n12750;
  assign n12768 = n12680 & n12767;
  assign n12769 = ~n12766 & ~n12768;
  assign n12770 = n12713 & n12764;
  assign n12771 = n12680 & n12713;
  assign n12772 = ~n12767 & ~n12771;
  assign n12773 = ~n12753 & ~n12772;
  assign n12774 = ~n12770 & ~n12773;
  assign n12775 = n12769 & n12774;
  assign n12776 = n12763 & ~n12775;
  assign n12777 = ~n12762 & ~n12776;
  assign n12778 = n12644 & ~n12645;
  assign n12779 = n12713 & ~n12750;
  assign n12780 = ~n12765 & ~n12779;
  assign n12781 = ~n12680 & ~n12780;
  assign n12782 = n12753 ^ n12680;
  assign n12783 = n12782 ^ n12771;
  assign n12784 = n12783 ^ n12782;
  assign n12785 = n12782 ^ n12680;
  assign n12786 = n12784 & ~n12785;
  assign n12787 = n12786 ^ n12782;
  assign n12788 = n12750 & ~n12787;
  assign n12789 = n12788 ^ n12782;
  assign n12790 = ~n12781 & n12789;
  assign n12791 = n12778 & n12790;
  assign n12792 = n12644 & n12645;
  assign n12793 = n12764 & n12779;
  assign n12794 = n12680 & n12753;
  assign n12795 = ~n12713 & n12794;
  assign n12796 = ~n12680 & ~n12753;
  assign n12797 = n12750 & n12796;
  assign n12798 = ~n12753 & ~n12780;
  assign n12799 = ~n12797 & ~n12798;
  assign n12800 = ~n12795 & n12799;
  assign n12801 = ~n12793 & n12800;
  assign n12802 = n12792 & ~n12801;
  assign n12803 = ~n12791 & ~n12802;
  assign n12804 = n12777 & n12803;
  assign n12805 = n12804 ^ n11800;
  assign n12806 = n12805 ^ x558;
  assign n12807 = n12298 & n12376;
  assign n12808 = n12363 & ~n12389;
  assign n12809 = ~n12807 & ~n12808;
  assign n12810 = ~n12366 & ~n12388;
  assign n12811 = n12387 & ~n12810;
  assign n12812 = ~n12358 & ~n12363;
  assign n12813 = ~n12358 & n12689;
  assign n12814 = ~n12361 & n12813;
  assign n12815 = ~n12388 & n12390;
  assign n12816 = ~n12363 & n12815;
  assign n12817 = ~n12814 & ~n12816;
  assign n12818 = ~n12376 & ~n12817;
  assign n12819 = ~n12812 & ~n12818;
  assign n12820 = ~n12811 & ~n12819;
  assign n12821 = n12397 ^ n12393;
  assign n12822 = n12393 ^ n12298;
  assign n12823 = n12822 ^ n12298;
  assign n12824 = n12387 ^ n12298;
  assign n12825 = ~n12823 & ~n12824;
  assign n12826 = n12825 ^ n12298;
  assign n12827 = n12821 & n12826;
  assign n12828 = n12827 ^ n12397;
  assign n12829 = n12380 & ~n12828;
  assign n12830 = ~n12398 & n12829;
  assign n12831 = ~n12371 & n12830;
  assign n12832 = n12831 ^ n12297;
  assign n12833 = n12832 ^ n12831;
  assign n12834 = n12831 ^ n12400;
  assign n12835 = n12834 ^ n12831;
  assign n12836 = ~n12833 & ~n12835;
  assign n12837 = n12836 ^ n12831;
  assign n12838 = n12695 & ~n12837;
  assign n12839 = n12838 ^ n12831;
  assign n12840 = n12820 & n12839;
  assign n12841 = n12809 & n12840;
  assign n12842 = n12686 & n12841;
  assign n12843 = n12370 & n12842;
  assign n12844 = n12843 ^ n10849;
  assign n12845 = n12844 ^ x498;
  assign n12846 = n11404 & ~n12729;
  assign n12847 = ~n11231 & n11427;
  assign n12848 = ~n11413 & ~n11426;
  assign n12849 = n11435 & n12848;
  assign n12850 = ~n11407 & n12849;
  assign n12851 = n11278 & ~n12850;
  assign n12852 = n11409 & ~n12737;
  assign n12853 = n11437 & n12730;
  assign n12854 = n11404 & ~n12853;
  assign n12855 = ~n12852 & ~n12854;
  assign n12856 = ~n12851 & n12855;
  assign n12857 = ~n11448 & ~n11452;
  assign n12858 = n11357 ^ n11355;
  assign n12859 = n12858 ^ n11317;
  assign n12860 = n12859 ^ n11355;
  assign n12861 = n12860 ^ n11400;
  assign n12862 = n11400 ^ n11317;
  assign n12863 = n11355 ^ n11317;
  assign n12864 = n12863 ^ n11317;
  assign n12865 = n12862 & n12864;
  assign n12866 = n12865 ^ n11317;
  assign n12867 = n12861 & n12866;
  assign n12868 = n12867 ^ n12858;
  assign n12869 = n11423 & ~n12868;
  assign n12870 = ~n12857 & ~n12869;
  assign n12871 = n12856 & n12870;
  assign n12872 = ~n12847 & n12871;
  assign n12873 = ~n12846 & n12872;
  assign n12874 = ~n12714 & n12873;
  assign n12875 = ~n11403 & n12874;
  assign n12876 = n12875 ^ n10882;
  assign n12877 = n12876 ^ x499;
  assign n12878 = n12204 & n12255;
  assign n12879 = ~n12251 & ~n12878;
  assign n12880 = ~n12239 & n12252;
  assign n12881 = n12179 & n12240;
  assign n12882 = n12257 & ~n12881;
  assign n12883 = ~n12880 & n12882;
  assign n12884 = n12249 & ~n12883;
  assign n12885 = n12240 & n12253;
  assign n12886 = n12265 & ~n12885;
  assign n12887 = n12178 & ~n12886;
  assign n12888 = ~n12884 & ~n12887;
  assign n12889 = ~n12238 & n12240;
  assign n12890 = n12206 & n12253;
  assign n12891 = n12890 ^ n12205;
  assign n12892 = ~n12889 & ~n12891;
  assign n12893 = ~n12880 & n12892;
  assign n12894 = n12270 & n12893;
  assign n12895 = n12240 & n12258;
  assign n12896 = ~n12208 & ~n12895;
  assign n12897 = ~n12880 & n12896;
  assign n12898 = ~n12251 & n12897;
  assign n12899 = n12282 & ~n12898;
  assign n12900 = ~n12894 & ~n12899;
  assign n12901 = n12888 & n12900;
  assign n12902 = n12879 & n12901;
  assign n12903 = n12902 ^ n10503;
  assign n12904 = n12903 ^ x497;
  assign n12905 = n11228 ^ x500;
  assign n12906 = n12904 & ~n12905;
  assign n12907 = ~n12877 & n12906;
  assign n12908 = n12845 & n12907;
  assign n12909 = n11592 & ~n12614;
  assign n12910 = ~n11587 & ~n12909;
  assign n12911 = ~n11615 & ~n11620;
  assign n12912 = n11471 & ~n12911;
  assign n12913 = ~n11607 & ~n11617;
  assign n12914 = n12606 & n12913;
  assign n12915 = n11593 & ~n12914;
  assign n12916 = ~n12912 & ~n12915;
  assign n12917 = n12910 & n12916;
  assign n12918 = ~n11594 & ~n11606;
  assign n12919 = n11577 & ~n12631;
  assign n12920 = ~n12918 & ~n12919;
  assign n12921 = n12917 & n12920;
  assign n12922 = ~n11604 & n12921;
  assign n12923 = n12608 & n12922;
  assign n12924 = n12604 & n12923;
  assign n12925 = n12924 ^ n10528;
  assign n12926 = n12925 ^ x496;
  assign n12927 = n11785 ^ x501;
  assign n12928 = n12926 & n12927;
  assign n12929 = n12877 & n12904;
  assign n12930 = n12845 & n12905;
  assign n12931 = n12929 & n12930;
  assign n12932 = n12928 & n12931;
  assign n12933 = n12926 & ~n12927;
  assign n12934 = n12904 & n12930;
  assign n12935 = ~n12877 & n12934;
  assign n12936 = n12933 & n12935;
  assign n12937 = ~n12932 & ~n12936;
  assign n12938 = ~n12905 & n12929;
  assign n12939 = ~n12845 & n12938;
  assign n12940 = n12928 & n12939;
  assign n12941 = ~n12845 & ~n12877;
  assign n12942 = n12906 & n12941;
  assign n12943 = n12928 & n12942;
  assign n12944 = ~n12926 & n12927;
  assign n12945 = ~n12904 & ~n12905;
  assign n12946 = n12877 & n12945;
  assign n12947 = ~n12845 & n12946;
  assign n12948 = ~n12904 & n12930;
  assign n12949 = n12877 & n12948;
  assign n12950 = ~n12947 & ~n12949;
  assign n12951 = n12944 & ~n12950;
  assign n12952 = ~n12943 & ~n12951;
  assign n12953 = n12941 & n12945;
  assign n12954 = n12944 & n12953;
  assign n12955 = n12905 ^ n12877;
  assign n12956 = n12905 ^ n12845;
  assign n12957 = n12955 & n12956;
  assign n12958 = n12904 & n12957;
  assign n12959 = n12933 & n12958;
  assign n12960 = ~n12954 & ~n12959;
  assign n12961 = ~n12926 & ~n12927;
  assign n12962 = n12939 & n12961;
  assign n12963 = ~n12877 & n12948;
  assign n12964 = n12944 & n12963;
  assign n12965 = ~n12962 & ~n12964;
  assign n12966 = n12931 & n12944;
  assign n12967 = n12928 & n12963;
  assign n12968 = ~n12966 & ~n12967;
  assign n12969 = ~n12904 & n12905;
  assign n12970 = n12877 & n12969;
  assign n12971 = ~n12845 & n12970;
  assign n12972 = ~n12927 & n12971;
  assign n12973 = ~n12928 & ~n12961;
  assign n12974 = ~n12944 & n12973;
  assign n12975 = n12941 & n12969;
  assign n12976 = ~n12974 & n12975;
  assign n12977 = ~n12972 & ~n12976;
  assign n12978 = n12845 & n12938;
  assign n12979 = ~n12935 & ~n12978;
  assign n12980 = ~n12942 & n12979;
  assign n12981 = n12961 & ~n12980;
  assign n12982 = n12977 & ~n12981;
  assign n12983 = n12845 & n12946;
  assign n12984 = ~n12973 & n12983;
  assign n12985 = n12905 & n12929;
  assign n12986 = ~n12845 & n12985;
  assign n12987 = n12944 & n12986;
  assign n12988 = ~n12984 & ~n12987;
  assign n12989 = ~n12877 & n12945;
  assign n12990 = n12845 & n12989;
  assign n12991 = n12926 & n12990;
  assign n12992 = n12933 & ~n12950;
  assign n12993 = ~n12991 & ~n12992;
  assign n12994 = n12988 & n12993;
  assign n12995 = n12982 & n12994;
  assign n12996 = n12968 & n12995;
  assign n12997 = n12965 & n12996;
  assign n12998 = n12960 & n12997;
  assign n12999 = n12952 & n12998;
  assign n13000 = ~n12940 & n12999;
  assign n13001 = n12937 & n13000;
  assign n13002 = ~n12908 & n13001;
  assign n13003 = n13002 ^ n11886;
  assign n13004 = n13003 ^ x557;
  assign n13005 = ~n12806 & n13004;
  assign n13006 = n11965 & ~n11979;
  assign n13007 = n11988 & ~n12118;
  assign n13008 = ~n13006 & ~n13007;
  assign n13009 = ~n11921 & n12108;
  assign n13010 = n11980 & n12001;
  assign n13011 = ~n13009 & ~n13010;
  assign n13012 = ~n11973 & ~n11982;
  assign n13013 = n11988 & ~n13012;
  assign n13014 = ~n11987 & ~n11999;
  assign n13015 = n12118 & n13014;
  assign n13016 = ~n11997 & n13015;
  assign n13017 = ~n11982 & n13016;
  assign n13018 = n11961 & ~n13017;
  assign n13019 = ~n13013 & ~n13018;
  assign n13022 = ~n11964 & ~n11973;
  assign n13023 = n12103 & n13022;
  assign n13020 = n11998 & ~n12095;
  assign n13021 = ~n12108 & n13020;
  assign n13024 = n13023 ^ n13021;
  assign n13025 = n13024 ^ n13023;
  assign n13026 = n13023 ^ n11960;
  assign n13027 = n13026 ^ n13023;
  assign n13028 = ~n13025 & ~n13027;
  assign n13029 = n13028 ^ n13023;
  assign n13030 = n11970 & ~n13029;
  assign n13031 = n13030 ^ n13023;
  assign n13032 = n13019 & n13031;
  assign n13033 = n13011 & n13032;
  assign n13034 = ~n12097 & n13033;
  assign n13035 = n13008 & n13034;
  assign n13036 = n13035 ^ n10154;
  assign n13037 = n13036 ^ x532;
  assign n13038 = n10820 & ~n12421;
  assign n13039 = ~n11171 & n11209;
  assign n13040 = ~n12424 & n13039;
  assign n13041 = ~n11199 & n13040;
  assign n13042 = n11159 & ~n13041;
  assign n13043 = ~n13038 & ~n13042;
  assign n13044 = ~n11200 & ~n11210;
  assign n13045 = n12429 & n13044;
  assign n13046 = n12445 & n13045;
  assign n13047 = n11174 & ~n13046;
  assign n13048 = n11178 & ~n11200;
  assign n13049 = ~n11194 & n13048;
  assign n13050 = n11157 & ~n13049;
  assign n13051 = n11212 & n12428;
  assign n13052 = n10821 & ~n13051;
  assign n13053 = ~n13050 & ~n13052;
  assign n13054 = ~n13047 & n13053;
  assign n13055 = n13043 & n13054;
  assign n13056 = ~n12426 & n13055;
  assign n13057 = n11169 & n13056;
  assign n13058 = n11163 & n13057;
  assign n13059 = n13058 ^ n10381;
  assign n13060 = n13059 ^ x537;
  assign n13061 = n13037 & n13060;
  assign n13062 = n12249 & ~n12280;
  assign n13063 = n12178 & ~n12290;
  assign n13064 = ~n13062 & ~n13063;
  assign n13065 = n12247 ^ n12176;
  assign n13066 = n13065 ^ n12247;
  assign n13067 = n12267 ^ n12247;
  assign n13068 = n13066 & n13067;
  assign n13069 = n13068 ^ n12247;
  assign n13070 = n12177 & n13069;
  assign n13071 = n13064 & ~n13070;
  assign n13072 = n13071 ^ n10393;
  assign n13073 = n13072 ^ x534;
  assign n13074 = n11639 & n11736;
  assign n13075 = ~n11760 & n12662;
  assign n13076 = ~n13074 & ~n13075;
  assign n13077 = ~n11708 & n11734;
  assign n13078 = n11721 & n11741;
  assign n13079 = n11710 & ~n13078;
  assign n13080 = n11734 & ~n12665;
  assign n13081 = ~n11715 & ~n11725;
  assign n13082 = ~n11747 & n13081;
  assign n13083 = n11639 & ~n13082;
  assign n13084 = ~n13080 & ~n13083;
  assign n13085 = n11722 & ~n11739;
  assign n13086 = n11738 & ~n13085;
  assign n13087 = ~n11707 & n12140;
  assign n13088 = ~n11761 & n13087;
  assign n13089 = n11710 & ~n13088;
  assign n13090 = ~n13086 & ~n13089;
  assign n13091 = n13084 & n13090;
  assign n13092 = ~n11732 & n13091;
  assign n13093 = ~n12142 & n13092;
  assign n13094 = ~n13079 & n13093;
  assign n13095 = ~n13077 & n13094;
  assign n13096 = n13076 & n13095;
  assign n13097 = ~n11781 & n13096;
  assign n13098 = ~n12141 & n13097;
  assign n13099 = n13098 ^ n10351;
  assign n13100 = n13099 ^ x535;
  assign n13101 = ~n13073 & ~n13100;
  assign n13102 = n11277 & ~n11441;
  assign n13103 = ~n11402 & n11456;
  assign n13104 = ~n11424 & n12724;
  assign n13105 = ~n11418 & n13104;
  assign n13106 = ~n11404 & n13105;
  assign n13107 = ~n13103 & ~n13106;
  assign n13108 = n13107 ^ n11277;
  assign n13109 = n13108 ^ n13107;
  assign n13110 = ~n11402 & n12732;
  assign n13111 = n13110 ^ n13107;
  assign n13112 = n13111 ^ n13107;
  assign n13113 = ~n13109 & ~n13112;
  assign n13114 = n13113 ^ n13107;
  assign n13115 = n11231 & n13114;
  assign n13116 = n13115 ^ n13107;
  assign n13117 = ~n13102 & ~n13116;
  assign n13118 = n11440 ^ n11278;
  assign n13119 = n11440 ^ n11409;
  assign n13120 = n13119 ^ n11409;
  assign n13121 = n12725 ^ n11409;
  assign n13122 = ~n13120 & n13121;
  assign n13123 = n13122 ^ n11409;
  assign n13124 = n13118 & n13123;
  assign n13125 = n13124 ^ n11278;
  assign n13126 = n13117 & ~n13125;
  assign n13127 = n12717 & n13126;
  assign n13128 = n11416 & n13127;
  assign n13129 = ~n11403 & n13128;
  assign n13130 = n13129 ^ n10125;
  assign n13131 = n13130 ^ x533;
  assign n13132 = n12297 & n12379;
  assign n13133 = n12394 & ~n12398;
  assign n13134 = n12363 & ~n13133;
  assign n13135 = ~n13132 & ~n13134;
  assign n13136 = n12353 & n12387;
  assign n13137 = ~n12361 & ~n12388;
  assign n13138 = n12358 & ~n13137;
  assign n13139 = ~n12376 & ~n12397;
  assign n13140 = ~n12695 & ~n13139;
  assign n13141 = ~n12393 & n12400;
  assign n13142 = ~n12378 & n13141;
  assign n13143 = n12358 & ~n13142;
  assign n13144 = ~n12365 & n12815;
  assign n13145 = n12298 & ~n13144;
  assign n13146 = ~n13143 & ~n13145;
  assign n13147 = ~n13140 & n13146;
  assign n13148 = n12385 ^ n12297;
  assign n13149 = n12390 ^ n12296;
  assign n13150 = n13149 ^ n12390;
  assign n13151 = ~n12353 & ~n12366;
  assign n13152 = n13151 ^ n12390;
  assign n13153 = ~n13150 & n13152;
  assign n13154 = n13153 ^ n12390;
  assign n13155 = n13154 ^ n12385;
  assign n13156 = n13148 & n13155;
  assign n13157 = n13156 ^ n13153;
  assign n13158 = n13157 ^ n12390;
  assign n13159 = n13158 ^ n12297;
  assign n13160 = n12385 & n13159;
  assign n13161 = n13160 ^ n12385;
  assign n13162 = n13161 ^ n12297;
  assign n13163 = n13147 & ~n13162;
  assign n13164 = ~n13138 & n13163;
  assign n13165 = ~n13136 & n13164;
  assign n13166 = n13135 & n13165;
  assign n13167 = n12683 & n13166;
  assign n13168 = n13167 ^ n10316;
  assign n13169 = n13168 ^ x536;
  assign n13170 = n13131 & n13169;
  assign n13171 = n13101 & n13170;
  assign n13172 = ~n13073 & n13100;
  assign n13173 = n13131 & ~n13169;
  assign n13174 = n13172 & n13173;
  assign n13175 = ~n13171 & ~n13174;
  assign n13176 = n13061 & ~n13175;
  assign n13177 = ~n13037 & n13060;
  assign n13178 = n13073 & ~n13100;
  assign n13179 = n13170 & n13178;
  assign n13180 = n13101 & n13173;
  assign n13181 = ~n13179 & ~n13180;
  assign n13182 = n13177 & ~n13181;
  assign n13183 = ~n13176 & ~n13182;
  assign n13184 = ~n13131 & n13169;
  assign n13185 = n13178 & n13184;
  assign n13186 = ~n13131 & ~n13169;
  assign n13187 = n13172 & n13186;
  assign n13188 = ~n13185 & ~n13187;
  assign n13189 = n13061 & ~n13188;
  assign n13190 = n13172 & n13184;
  assign n13191 = n13177 & n13190;
  assign n13192 = ~n13037 & ~n13060;
  assign n13193 = n13173 & n13178;
  assign n13194 = ~n13171 & ~n13193;
  assign n13195 = n13192 & ~n13194;
  assign n13196 = ~n13191 & ~n13195;
  assign n13197 = ~n13189 & n13196;
  assign n13198 = n13174 & n13177;
  assign n13199 = n13170 & n13172;
  assign n13200 = n13073 & n13100;
  assign n13201 = n13173 & n13200;
  assign n13202 = ~n13199 & ~n13201;
  assign n13203 = n13192 & ~n13202;
  assign n13204 = ~n13198 & ~n13203;
  assign n13205 = n13037 & ~n13060;
  assign n13206 = n13184 & n13200;
  assign n13207 = n13131 ^ n13100;
  assign n13208 = n13207 ^ n13169;
  assign n13209 = n13131 ^ n13073;
  assign n13210 = ~n13208 & ~n13209;
  assign n13211 = ~n13206 & ~n13210;
  assign n13212 = n13188 & n13211;
  assign n13213 = ~n13171 & n13212;
  assign n13214 = n13205 & n13213;
  assign n13215 = n13101 & n13184;
  assign n13216 = n13186 & n13200;
  assign n13217 = ~n13215 & ~n13216;
  assign n13218 = n13188 & n13217;
  assign n13219 = ~n13037 & ~n13218;
  assign n13220 = n13101 & n13186;
  assign n13221 = ~n13206 & ~n13220;
  assign n13222 = ~n13201 & n13221;
  assign n13223 = ~n13193 & n13222;
  assign n13224 = n13061 & ~n13223;
  assign n13225 = ~n13219 & ~n13224;
  assign n13226 = ~n13214 & n13225;
  assign n13227 = n13204 & n13226;
  assign n13228 = n13197 & n13227;
  assign n13229 = n13183 & n13228;
  assign n13230 = n13229 ^ n11822;
  assign n13231 = n13230 ^ x560;
  assign n13232 = n12294 ^ x526;
  assign n13233 = n13130 ^ x531;
  assign n13234 = n13232 & n13233;
  assign n13235 = n13036 ^ x530;
  assign n13236 = n12173 ^ x527;
  assign n13237 = ~n13235 & ~n13236;
  assign n13238 = ~n11611 & ~n11616;
  assign n13239 = n11577 & ~n13238;
  assign n13240 = ~n11593 & n12606;
  assign n13241 = ~n11622 & ~n13240;
  assign n13242 = ~n11615 & n12606;
  assign n13243 = n11508 & ~n13242;
  assign n13244 = ~n13241 & ~n13243;
  assign n13245 = ~n11599 & n13244;
  assign n13246 = n11471 & ~n13245;
  assign n13247 = ~n13239 & ~n13246;
  assign n13248 = n11508 & n11607;
  assign n13249 = ~n11591 & n11606;
  assign n13250 = ~n11586 & n13249;
  assign n13251 = n11593 & ~n13250;
  assign n13252 = ~n13248 & ~n13251;
  assign n13253 = ~n11605 & ~n11617;
  assign n13254 = n11592 & ~n13253;
  assign n13255 = n11591 ^ n11471;
  assign n13256 = ~n11575 & n12600;
  assign n13257 = n13256 ^ n11507;
  assign n13258 = n13257 ^ n13256;
  assign n13259 = ~n11599 & n13238;
  assign n13260 = n13259 ^ n13256;
  assign n13261 = n13258 & n13260;
  assign n13262 = n13261 ^ n13256;
  assign n13263 = n13262 ^ n11591;
  assign n13264 = n13255 & ~n13263;
  assign n13265 = n13264 ^ n13261;
  assign n13266 = n13265 ^ n13256;
  assign n13267 = n13266 ^ n11471;
  assign n13268 = ~n11591 & ~n13267;
  assign n13269 = n13268 ^ n11591;
  assign n13270 = n13269 ^ n11471;
  assign n13271 = ~n13254 & ~n13270;
  assign n13272 = n13252 & n13271;
  assign n13273 = n13247 & n13272;
  assign n13274 = n11584 & n13273;
  assign n13275 = n12604 & n13274;
  assign n13276 = n13275 ^ n10181;
  assign n13277 = n13276 ^ x528;
  assign n13278 = ~n10687 & ~n10701;
  assign n13279 = n10670 & ~n13278;
  assign n13280 = ~n10678 & ~n13279;
  assign n13281 = ~n10668 & ~n10705;
  assign n13282 = ~n10693 & ~n13281;
  assign n13283 = n10700 & n10707;
  assign n13284 = ~n10689 & n13283;
  assign n13285 = ~n10281 & n13284;
  assign n13286 = n10665 & ~n13285;
  assign n13287 = n10675 & ~n12488;
  assign n13288 = ~n10692 & n10707;
  assign n13289 = ~n10698 & n12498;
  assign n13290 = ~n10687 & n13289;
  assign n13291 = ~n13288 & ~n13290;
  assign n13292 = ~n10679 & ~n13291;
  assign n13293 = n10664 & ~n13292;
  assign n13294 = ~n13287 & ~n13293;
  assign n13295 = ~n13286 & n13294;
  assign n13296 = ~n13282 & n13295;
  assign n13297 = n10694 ^ n10664;
  assign n13298 = n13297 ^ n10694;
  assign n13299 = n12472 ^ n10694;
  assign n13300 = n13299 ^ n10694;
  assign n13301 = ~n13298 & ~n13300;
  assign n13302 = n13301 ^ n10694;
  assign n13303 = ~n10469 & n13302;
  assign n13304 = n13303 ^ n10694;
  assign n13305 = n13296 & ~n13304;
  assign n13306 = n13280 & n13305;
  assign n13307 = n12479 & n13306;
  assign n13308 = n10674 & n13307;
  assign n13309 = n13308 ^ n10208;
  assign n13310 = n13309 ^ x529;
  assign n13311 = n13277 & n13310;
  assign n13312 = n13237 & n13311;
  assign n13313 = n13235 & ~n13236;
  assign n13314 = n13277 & ~n13310;
  assign n13315 = n13313 & n13314;
  assign n13316 = ~n13312 & ~n13315;
  assign n13317 = n13234 & ~n13316;
  assign n13318 = n13235 & n13236;
  assign n13319 = n13311 & n13318;
  assign n13320 = n13234 & n13319;
  assign n13321 = ~n13232 & ~n13233;
  assign n13322 = ~n13277 & ~n13310;
  assign n13323 = n13318 & n13322;
  assign n13324 = n13321 & n13323;
  assign n13325 = ~n13320 & ~n13324;
  assign n13326 = ~n13235 & n13236;
  assign n13327 = n13314 & n13326;
  assign n13328 = n13234 & n13327;
  assign n13329 = ~n13232 & n13233;
  assign n13330 = n13237 & n13322;
  assign n13331 = ~n13315 & ~n13330;
  assign n13332 = n13329 & ~n13331;
  assign n13333 = ~n13328 & ~n13332;
  assign n13334 = n13232 & ~n13233;
  assign n13335 = ~n13277 & n13310;
  assign n13336 = n13313 & n13335;
  assign n13337 = ~n13330 & ~n13336;
  assign n13338 = ~n13327 & n13337;
  assign n13339 = n13334 & ~n13338;
  assign n13340 = n13326 & n13335;
  assign n13341 = ~n13319 & ~n13340;
  assign n13342 = n13334 & ~n13341;
  assign n13343 = n13311 & n13313;
  assign n13344 = n13237 & n13314;
  assign n13345 = ~n13343 & ~n13344;
  assign n13346 = n13329 & ~n13345;
  assign n13347 = ~n13234 & ~n13321;
  assign n13348 = n13237 & n13335;
  assign n13349 = ~n13347 & n13348;
  assign n13350 = n13236 ^ n13235;
  assign n13351 = n13310 ^ n13236;
  assign n13352 = n13351 ^ n13236;
  assign n13353 = n13310 ^ n13277;
  assign n13354 = n13353 ^ n13236;
  assign n13355 = ~n13352 & ~n13354;
  assign n13356 = n13355 ^ n13236;
  assign n13357 = ~n13350 & n13356;
  assign n13358 = n13357 ^ n13353;
  assign n13359 = n13321 & ~n13358;
  assign n13360 = ~n13349 & ~n13359;
  assign n13361 = n13322 & n13326;
  assign n13362 = n13314 & n13318;
  assign n13363 = ~n13361 & ~n13362;
  assign n13364 = ~n13336 & n13363;
  assign n13365 = n13234 & ~n13364;
  assign n13366 = n13318 & n13335;
  assign n13367 = n13316 & ~n13366;
  assign n13368 = n13334 & ~n13367;
  assign n13369 = ~n13323 & ~n13340;
  assign n13370 = ~n13319 & n13369;
  assign n13371 = ~n13327 & n13370;
  assign n13372 = n13329 & ~n13371;
  assign n13373 = ~n13368 & ~n13372;
  assign n13374 = ~n13365 & n13373;
  assign n13375 = n13360 & n13374;
  assign n13376 = ~n13346 & n13375;
  assign n13377 = ~n13342 & n13376;
  assign n13378 = ~n13339 & n13377;
  assign n13379 = n13333 & n13378;
  assign n13380 = n13325 & n13379;
  assign n13381 = ~n13317 & n13380;
  assign n13382 = n13381 ^ n11853;
  assign n13383 = n13382 ^ x559;
  assign n13384 = ~n13231 & n13383;
  assign n13385 = n13005 & n13384;
  assign n13386 = n12806 & ~n13004;
  assign n13387 = n13384 & n13386;
  assign n13388 = n13231 & ~n13383;
  assign n13389 = n13386 & n13388;
  assign n13390 = ~n13387 & ~n13389;
  assign n13391 = ~n13385 & n13390;
  assign n13392 = n12599 & ~n13391;
  assign n13393 = ~n12093 & n12598;
  assign n13394 = ~n13231 & ~n13383;
  assign n13395 = n13386 & n13394;
  assign n13396 = ~n13389 & ~n13395;
  assign n13397 = n13393 & ~n13396;
  assign n13398 = ~n12093 & ~n12598;
  assign n13399 = n13231 & n13383;
  assign n13400 = ~n12806 & ~n13004;
  assign n13401 = n13399 & n13400;
  assign n13402 = n13384 & n13400;
  assign n13403 = ~n13401 & ~n13402;
  assign n13404 = n13386 & n13399;
  assign n13405 = n13394 & n13400;
  assign n13406 = ~n13404 & ~n13405;
  assign n13407 = n13403 & n13406;
  assign n13408 = n13398 & ~n13407;
  assign n13409 = n12806 & n13004;
  assign n13410 = n13399 & n13409;
  assign n13411 = n12599 & n13410;
  assign n13412 = n13005 & n13399;
  assign n13413 = n13393 & n13412;
  assign n13414 = n13005 & n13388;
  assign n13415 = n13005 & n13394;
  assign n13416 = ~n13410 & ~n13415;
  assign n13417 = ~n13414 & n13416;
  assign n13418 = n13393 & ~n13417;
  assign n13419 = n13388 & n13409;
  assign n13420 = ~n13415 & ~n13419;
  assign n13421 = ~n13412 & n13420;
  assign n13422 = n12599 & ~n13421;
  assign n13423 = ~n13418 & ~n13422;
  assign n13424 = n13384 & n13409;
  assign n13425 = n13394 & n13409;
  assign n13426 = ~n13424 & ~n13425;
  assign n13427 = ~n13414 & n13426;
  assign n13428 = ~n13419 & n13427;
  assign n13429 = n13398 & ~n13428;
  assign n13431 = ~n13395 & n13403;
  assign n13432 = ~n13404 & n13431;
  assign n13430 = ~n13415 & n13427;
  assign n13433 = n13432 ^ n13430;
  assign n13434 = n12093 & n12598;
  assign n13435 = n13434 ^ n13432;
  assign n13436 = n13432 & n13435;
  assign n13437 = n13436 ^ n13432;
  assign n13438 = n13433 & n13437;
  assign n13439 = n13438 ^ n13436;
  assign n13440 = n13439 ^ n13432;
  assign n13441 = n13440 ^ n13434;
  assign n13442 = ~n13429 & n13441;
  assign n13443 = n13442 ^ n13429;
  assign n13444 = n13423 & ~n13443;
  assign n13445 = ~n13413 & n13444;
  assign n13446 = ~n13411 & n13445;
  assign n13447 = ~n13408 & n13446;
  assign n13448 = n12598 ^ n12093;
  assign n13449 = n13405 ^ n12598;
  assign n13450 = n13449 ^ n13405;
  assign n13451 = n13388 & n13400;
  assign n13452 = ~n13387 & ~n13451;
  assign n13453 = n13452 ^ n13405;
  assign n13454 = n13450 & ~n13453;
  assign n13455 = n13454 ^ n13405;
  assign n13456 = n13448 & n13455;
  assign n13457 = n13447 & ~n13456;
  assign n13458 = ~n13397 & n13457;
  assign n13459 = ~n13392 & n13458;
  assign n13460 = n13459 ^ n12136;
  assign n13461 = n13460 ^ x614;
  assign n13462 = n12282 & ~n12886;
  assign n13463 = n12249 & ~n12893;
  assign n13464 = n12270 & ~n12883;
  assign n13465 = ~n13463 & ~n13464;
  assign n13466 = ~n13462 & n13465;
  assign n13467 = n12898 ^ n12879;
  assign n13468 = n13467 ^ n12879;
  assign n13469 = n12879 ^ n12176;
  assign n13470 = n13469 ^ n12879;
  assign n13471 = n13468 & ~n13470;
  assign n13472 = n13471 ^ n12879;
  assign n13473 = ~n12177 & ~n13472;
  assign n13474 = n13473 ^ n12879;
  assign n13475 = n13466 & n13474;
  assign n13476 = n13475 ^ n11034;
  assign n13477 = n13476 ^ x510;
  assign n13478 = n10735 ^ x509;
  assign n13479 = n13477 & ~n13478;
  assign n13480 = n12643 ^ x512;
  assign n13481 = ~n11199 & n13044;
  assign n13482 = n11174 & ~n13481;
  assign n13483 = n11211 & n12428;
  assign n13484 = n11157 & ~n13483;
  assign n13485 = ~n13482 & ~n13484;
  assign n13486 = ~n11201 & n11211;
  assign n13487 = ~n11199 & n13486;
  assign n13488 = n10821 & ~n13487;
  assign n13489 = ~n11152 & ~n11192;
  assign n13490 = n11159 & ~n13489;
  assign n13491 = ~n11155 & n11172;
  assign n13492 = n11174 & ~n13491;
  assign n13493 = ~n12424 & n12428;
  assign n13494 = ~n11161 & n13493;
  assign n13495 = n11159 & ~n13494;
  assign n13496 = ~n13492 & ~n13495;
  assign n13497 = n11192 ^ n10777;
  assign n13498 = ~n11171 & n11178;
  assign n13499 = n13498 ^ n11209;
  assign n13500 = n11209 ^ n10820;
  assign n13501 = n13500 ^ n11209;
  assign n13502 = n13499 & ~n13501;
  assign n13503 = n13502 ^ n11209;
  assign n13504 = n13503 ^ n11192;
  assign n13505 = n13497 & ~n13504;
  assign n13506 = n13505 ^ n13502;
  assign n13507 = n13506 ^ n11209;
  assign n13508 = n13507 ^ n10777;
  assign n13509 = ~n11192 & ~n13508;
  assign n13510 = n13509 ^ n11192;
  assign n13511 = n13510 ^ n10777;
  assign n13512 = n13496 & ~n13511;
  assign n13513 = ~n11153 & n13512;
  assign n13514 = ~n13490 & n13513;
  assign n13515 = ~n13488 & n13514;
  assign n13516 = n13485 & n13515;
  assign n13517 = n12423 & n13516;
  assign n13518 = n13517 ^ n11017;
  assign n13519 = n13518 ^ x511;
  assign n13520 = ~n13480 & ~n13519;
  assign n13521 = n13479 & n13520;
  assign n13522 = n11469 ^ x508;
  assign n13523 = n12712 ^ x513;
  assign n13524 = ~n13522 & ~n13523;
  assign n13525 = n13521 & n13524;
  assign n13526 = n13522 & n13523;
  assign n13527 = n13521 & n13526;
  assign n13528 = ~n13477 & n13478;
  assign n13529 = n13480 & n13519;
  assign n13530 = n13528 & n13529;
  assign n13531 = ~n13522 & n13523;
  assign n13532 = n13530 & n13531;
  assign n13533 = ~n13477 & ~n13478;
  assign n13534 = n13529 & n13533;
  assign n13535 = n13526 & n13534;
  assign n13536 = ~n13532 & ~n13535;
  assign n13537 = ~n13527 & n13536;
  assign n13538 = n13477 & n13478;
  assign n13539 = n13520 & n13538;
  assign n13540 = n13480 & ~n13519;
  assign n13541 = n13528 & n13540;
  assign n13542 = ~n13539 & ~n13541;
  assign n13543 = n13526 & ~n13542;
  assign n13544 = n13522 & ~n13523;
  assign n13545 = ~n13531 & ~n13544;
  assign n13546 = n13521 & ~n13545;
  assign n13547 = ~n13543 & ~n13546;
  assign n13548 = n13519 ^ n13480;
  assign n13549 = n13480 ^ n13477;
  assign n13550 = n13549 ^ n13519;
  assign n13551 = n13550 ^ n13480;
  assign n13552 = ~n13548 & ~n13551;
  assign n13553 = n13552 ^ n13480;
  assign n13554 = n13478 & n13553;
  assign n13555 = n13554 ^ n13550;
  assign n13556 = n13531 & ~n13555;
  assign n13557 = ~n13480 & n13519;
  assign n13558 = n13538 & n13557;
  assign n13559 = n13529 & n13538;
  assign n13560 = n13533 & n13540;
  assign n13561 = n13479 & n13529;
  assign n13562 = n13542 & ~n13561;
  assign n13563 = ~n13560 & n13562;
  assign n13564 = ~n13559 & n13563;
  assign n13565 = ~n13530 & n13564;
  assign n13566 = ~n13558 & n13565;
  assign n13567 = n13544 & ~n13566;
  assign n13568 = ~n13556 & ~n13567;
  assign n13569 = n13523 ^ n13522;
  assign n13570 = n13528 & n13557;
  assign n13571 = ~n13559 & ~n13570;
  assign n13572 = n13479 & n13557;
  assign n13573 = n13479 & n13540;
  assign n13574 = ~n13572 & ~n13573;
  assign n13575 = n13571 & n13574;
  assign n13576 = n13575 ^ n13523;
  assign n13577 = n13576 ^ n13575;
  assign n13578 = n13538 & n13540;
  assign n13579 = n13571 & ~n13578;
  assign n13580 = ~n13560 & n13579;
  assign n13581 = n13533 & n13557;
  assign n13582 = n13574 & ~n13581;
  assign n13583 = n13580 & n13582;
  assign n13584 = n13583 ^ n13575;
  assign n13585 = ~n13577 & n13584;
  assign n13586 = n13585 ^ n13575;
  assign n13587 = ~n13569 & ~n13586;
  assign n13588 = n13568 & ~n13587;
  assign n13589 = n13547 & n13588;
  assign n13590 = n13537 & n13589;
  assign n13591 = ~n13525 & n13590;
  assign n13592 = n13591 ^ n11698;
  assign n13593 = n13592 ^ x588;
  assign n13594 = n13329 & n13348;
  assign n13595 = n13311 & n13326;
  assign n13596 = ~n13366 & ~n13595;
  assign n13597 = n13321 & ~n13596;
  assign n13598 = ~n13594 & ~n13597;
  assign n13599 = n13321 & n13336;
  assign n13600 = n13327 & ~n13347;
  assign n13601 = ~n13599 & ~n13600;
  assign n13602 = n13313 & n13322;
  assign n13603 = n13337 & n13363;
  assign n13604 = ~n13602 & n13603;
  assign n13605 = n13334 & ~n13604;
  assign n13606 = ~n13366 & n13369;
  assign n13607 = ~n13361 & n13606;
  assign n13608 = n13329 & ~n13607;
  assign n13609 = ~n13605 & ~n13608;
  assign n13610 = n13369 & ~n13595;
  assign n13611 = n13234 & ~n13610;
  assign n13612 = n13233 ^ n13232;
  assign n13613 = ~n13312 & n13331;
  assign n13614 = ~n13602 & n13613;
  assign n13615 = n13614 ^ n13337;
  assign n13616 = n13337 ^ n13233;
  assign n13617 = n13616 ^ n13337;
  assign n13618 = n13615 & ~n13617;
  assign n13619 = n13618 ^ n13337;
  assign n13620 = ~n13612 & ~n13619;
  assign n13621 = ~n13611 & ~n13620;
  assign n13622 = n13609 & n13621;
  assign n13623 = n13601 & n13622;
  assign n13624 = ~n13346 & n13623;
  assign n13625 = n13598 & n13624;
  assign n13626 = ~n13342 & n13625;
  assign n13627 = n13362 ^ n13233;
  assign n13628 = n13627 ^ n13362;
  assign n13629 = n13362 ^ n13344;
  assign n13630 = ~n13628 & n13629;
  assign n13631 = n13630 ^ n13362;
  assign n13632 = n13612 & n13631;
  assign n13633 = n13626 & ~n13632;
  assign n13634 = ~n13317 & n13633;
  assign n13635 = n13634 ^ n11506;
  assign n13636 = n13635 ^ x587;
  assign n13637 = ~n13593 & n13636;
  assign n13638 = ~n13171 & ~n13180;
  assign n13639 = n13205 & ~n13638;
  assign n13640 = n13060 ^ n13037;
  assign n13641 = n13188 & n13202;
  assign n13642 = n13640 & ~n13641;
  assign n13643 = ~n13639 & ~n13642;
  assign n13644 = n13177 & ~n13221;
  assign n13645 = n13061 & n13210;
  assign n13646 = ~n13644 & ~n13645;
  assign n13647 = n13643 & n13646;
  assign n13648 = n13178 & n13186;
  assign n13649 = ~n13215 & ~n13648;
  assign n13650 = n13037 & ~n13649;
  assign n13651 = n13192 & n13213;
  assign n13652 = ~n13650 & ~n13651;
  assign n13653 = n13647 & n13652;
  assign n13654 = n13183 & n13653;
  assign n13655 = n13654 ^ n10468;
  assign n13656 = n13655 ^ x590;
  assign n13657 = ~n12949 & ~n12990;
  assign n13658 = n12928 & ~n13657;
  assign n13659 = ~n12975 & ~n12990;
  assign n13660 = n12961 & ~n13659;
  assign n13661 = ~n13658 & ~n13660;
  assign n13662 = n12928 & n12935;
  assign n13663 = ~n12964 & ~n13662;
  assign n13664 = ~n12908 & ~n12958;
  assign n13665 = n12944 & ~n13664;
  assign n13666 = ~n12927 & n12939;
  assign n13667 = ~n12949 & n12979;
  assign n13668 = ~n12953 & n13667;
  assign n13669 = n12961 & ~n13668;
  assign n13670 = ~n13666 & ~n13669;
  assign n13671 = n12933 & n12963;
  assign n13672 = ~n12947 & ~n12986;
  assign n13673 = ~n12942 & n13672;
  assign n13674 = n12928 & ~n13673;
  assign n13675 = n12933 & n12942;
  assign n13676 = n12908 & n12933;
  assign n13677 = ~n12971 & ~n12990;
  assign n13678 = n12944 & ~n13677;
  assign n13679 = ~n13676 & ~n13678;
  assign n13680 = n12960 & n13679;
  assign n13681 = ~n13675 & n13680;
  assign n13682 = ~n13674 & n13681;
  assign n13683 = ~n13671 & n13682;
  assign n13684 = n13670 & n13683;
  assign n13685 = n12968 & n13684;
  assign n13686 = ~n13665 & n13685;
  assign n13687 = n12931 ^ n12926;
  assign n13688 = n13687 ^ n12931;
  assign n13689 = ~n12971 & ~n12983;
  assign n13690 = n13689 ^ n12931;
  assign n13691 = n13688 & ~n13690;
  assign n13692 = n13691 ^ n12931;
  assign n13693 = ~n12927 & n13692;
  assign n13694 = n13686 & ~n13693;
  assign n13695 = n13663 & n13694;
  assign n13696 = n13661 & n13695;
  assign n13697 = ~n12940 & n13696;
  assign n13698 = n13697 ^ n11673;
  assign n13699 = n13698 ^ x589;
  assign n13700 = n13656 & ~n13699;
  assign n13701 = n13637 & n13700;
  assign n13702 = ~n12790 & n12792;
  assign n13703 = n12761 & n12763;
  assign n13704 = ~n13702 & ~n13703;
  assign n13705 = n12775 ^ n12644;
  assign n13706 = n13705 ^ n12775;
  assign n13707 = n12800 ^ n12775;
  assign n13708 = n13706 & n13707;
  assign n13709 = n13708 ^ n12775;
  assign n13710 = ~n12645 & ~n13709;
  assign n13711 = n13704 & ~n13710;
  assign n13712 = ~n12793 & n13711;
  assign n13713 = n13712 ^ n9354;
  assign n13714 = n13713 ^ x591;
  assign n13715 = n12020 & n12026;
  assign n13716 = ~n12020 & n12071;
  assign n13717 = n12053 & ~n13716;
  assign n13718 = n12053 & n12074;
  assign n13719 = ~n12047 & ~n12070;
  assign n13720 = n12054 & n13719;
  assign n13721 = n12042 & ~n13720;
  assign n13722 = n12026 & n12078;
  assign n13723 = n11230 & ~n12071;
  assign n13724 = ~n13722 & ~n13723;
  assign n13725 = ~n12024 & n12045;
  assign n13726 = ~n12029 & n13725;
  assign n13727 = n11230 & ~n13726;
  assign n13728 = ~n12037 & n12066;
  assign n13729 = ~n12033 & n13728;
  assign n13730 = n12042 & ~n13729;
  assign n13731 = ~n13727 & ~n13730;
  assign n13732 = ~n12047 & ~n12074;
  assign n13733 = n12026 & ~n13732;
  assign n13734 = ~n12053 & n12066;
  assign n13735 = ~n12038 & ~n12067;
  assign n13736 = ~n12078 & n13735;
  assign n13737 = ~n12029 & n13736;
  assign n13738 = ~n13734 & ~n13737;
  assign n13739 = ~n12073 & ~n13738;
  assign n13740 = ~n12068 & ~n13739;
  assign n13741 = ~n13733 & ~n13740;
  assign n13742 = n13731 & n13741;
  assign n13743 = n13724 & n13742;
  assign n13744 = ~n13721 & n13743;
  assign n13745 = ~n13718 & n13744;
  assign n13746 = n12041 & n13745;
  assign n13747 = ~n13717 & n13746;
  assign n13748 = ~n13715 & n13747;
  assign n13749 = n13748 ^ n11546;
  assign n13750 = n13749 ^ x586;
  assign n13751 = n13714 & ~n13750;
  assign n13752 = n13701 & n13751;
  assign n13753 = ~n13593 & ~n13636;
  assign n13754 = n13656 & n13699;
  assign n13755 = n13753 & n13754;
  assign n13756 = n13593 & ~n13636;
  assign n13757 = ~n13656 & ~n13699;
  assign n13758 = n13756 & n13757;
  assign n13759 = ~n13755 & ~n13758;
  assign n13760 = ~n13714 & ~n13750;
  assign n13761 = ~n13759 & n13760;
  assign n13762 = ~n13752 & ~n13761;
  assign n13763 = ~n13656 & n13699;
  assign n13764 = n13753 & n13763;
  assign n13765 = ~n13714 & n13750;
  assign n13766 = n13764 & n13765;
  assign n13767 = n13700 & n13756;
  assign n13768 = n13765 & n13767;
  assign n13769 = n13714 & n13750;
  assign n13770 = n13764 & n13769;
  assign n13771 = ~n13768 & ~n13770;
  assign n13772 = ~n13766 & n13771;
  assign n13773 = n13756 & n13763;
  assign n13774 = n13760 & n13773;
  assign n13775 = n13637 & n13757;
  assign n13776 = n13751 & n13775;
  assign n13777 = ~n13774 & ~n13776;
  assign n13778 = ~n13759 & n13765;
  assign n13779 = n13636 ^ n13593;
  assign n13780 = n13779 ^ n13656;
  assign n13781 = n13780 ^ n13779;
  assign n13782 = n13779 ^ n13636;
  assign n13783 = n13782 ^ n13779;
  assign n13784 = ~n13781 & n13783;
  assign n13785 = n13784 ^ n13779;
  assign n13786 = n13699 & ~n13785;
  assign n13787 = n13786 ^ n13779;
  assign n13788 = n13769 & ~n13787;
  assign n13789 = ~n13778 & ~n13788;
  assign n13790 = n13754 & n13756;
  assign n13791 = ~n13760 & ~n13769;
  assign n13792 = n13790 & ~n13791;
  assign n13793 = n13593 & n13636;
  assign n13794 = n13700 & n13793;
  assign n13795 = n13754 & n13793;
  assign n13796 = n13759 & ~n13790;
  assign n13797 = ~n13773 & n13796;
  assign n13798 = ~n13795 & n13797;
  assign n13799 = ~n13794 & n13798;
  assign n13800 = n13751 & ~n13799;
  assign n13801 = n13765 ^ n13760;
  assign n13806 = n13763 & n13793;
  assign n13807 = n13637 & n13754;
  assign n13808 = ~n13775 & ~n13807;
  assign n13809 = ~n13795 & n13808;
  assign n13810 = ~n13806 & n13809;
  assign n13802 = n13637 & n13763;
  assign n13803 = ~n13775 & ~n13794;
  assign n13804 = ~n13802 & n13803;
  assign n13805 = ~n13701 & n13804;
  assign n13811 = n13810 ^ n13805;
  assign n13812 = n13810 ^ n13760;
  assign n13813 = n13812 ^ n13810;
  assign n13814 = ~n13811 & n13813;
  assign n13815 = n13814 ^ n13810;
  assign n13816 = n13801 & n13815;
  assign n13817 = n13816 ^ n13765;
  assign n13818 = ~n13800 & ~n13817;
  assign n13819 = ~n13792 & n13818;
  assign n13820 = n13789 & n13819;
  assign n13821 = n13777 & n13820;
  assign n13822 = n13772 & n13821;
  assign n13823 = n13762 & n13822;
  assign n13824 = n13823 ^ n12679;
  assign n13825 = n13824 ^ x613;
  assign n13826 = ~n13190 & ~n13220;
  assign n13827 = ~n13185 & n13826;
  assign n13828 = ~n13216 & n13827;
  assign n13829 = n13061 & ~n13828;
  assign n13830 = ~n13179 & ~n13187;
  assign n13831 = ~n13171 & n13830;
  assign n13832 = ~n13201 & n13831;
  assign n13833 = n13177 & ~n13832;
  assign n13834 = ~n13193 & n13827;
  assign n13835 = n13192 & ~n13834;
  assign n13836 = ~n13833 & ~n13835;
  assign n13841 = ~n13174 & n13831;
  assign n13837 = n13170 & n13200;
  assign n13838 = ~n13174 & ~n13837;
  assign n13839 = ~n13179 & n13838;
  assign n13840 = ~n13193 & n13839;
  assign n13842 = n13841 ^ n13840;
  assign n13843 = n13841 ^ n13060;
  assign n13844 = n13843 ^ n13841;
  assign n13845 = n13842 & n13844;
  assign n13846 = n13845 ^ n13841;
  assign n13847 = n13037 & ~n13846;
  assign n13848 = n13836 & ~n13847;
  assign n13849 = ~n13829 & n13848;
  assign n13850 = ~n13206 & ~n13216;
  assign n13851 = n13649 & n13850;
  assign n13852 = n13851 ^ n13060;
  assign n13853 = n13852 ^ n13851;
  assign n13854 = ~n13180 & ~n13837;
  assign n13855 = n13202 & n13854;
  assign n13856 = n13855 ^ n13851;
  assign n13857 = n13856 ^ n13851;
  assign n13858 = ~n13853 & ~n13857;
  assign n13859 = n13858 ^ n13851;
  assign n13860 = ~n13640 & ~n13859;
  assign n13861 = n13860 ^ n13851;
  assign n13862 = n13849 & n13861;
  assign n13863 = n13862 ^ n12323;
  assign n13864 = n13863 ^ x553;
  assign n13865 = n13544 & n13560;
  assign n13866 = n13524 & ~n13571;
  assign n13867 = ~n13865 & ~n13866;
  assign n13868 = n13520 & n13533;
  assign n13869 = ~n13558 & ~n13578;
  assign n13870 = n13571 & n13869;
  assign n13871 = ~n13868 & n13870;
  assign n13872 = n13544 & ~n13871;
  assign n13873 = n13524 & ~n13555;
  assign n13874 = ~n13872 & ~n13873;
  assign n13875 = ~n13572 & n13580;
  assign n13876 = ~n13530 & n13875;
  assign n13877 = n13531 & ~n13876;
  assign n13878 = n13534 & ~n13545;
  assign n13879 = n13520 & n13528;
  assign n13880 = n13582 & ~n13879;
  assign n13881 = ~n13561 & n13880;
  assign n13882 = ~n13530 & n13881;
  assign n13883 = n13526 & ~n13882;
  assign n13884 = ~n13878 & ~n13883;
  assign n13885 = ~n13877 & n13884;
  assign n13886 = n13874 & n13885;
  assign n13887 = n13867 & n13886;
  assign n13888 = n13547 & n13887;
  assign n13889 = n13888 ^ n12349;
  assign n13890 = n13889 ^ x552;
  assign n13891 = ~n13864 & n13890;
  assign n13892 = n12903 ^ x543;
  assign n13893 = n13168 ^ x538;
  assign n13894 = ~n13892 & n13893;
  assign n13895 = n11965 & ~n11998;
  assign n13896 = n11987 & n11988;
  assign n13897 = ~n13895 & ~n13896;
  assign n13898 = n11979 & ~n12095;
  assign n13899 = n11961 & ~n13898;
  assign n13900 = ~n11973 & ~n11999;
  assign n13901 = ~n12108 & n13900;
  assign n13902 = n12001 & ~n13901;
  assign n13903 = ~n11889 & n13022;
  assign n13904 = ~n11982 & n13903;
  assign n13905 = n11965 & ~n13904;
  assign n13906 = n12001 & ~n12121;
  assign n13907 = ~n13905 & ~n13906;
  assign n13908 = ~n11969 & n13014;
  assign n13909 = n11961 & ~n13908;
  assign n13910 = n11979 & n11998;
  assign n13911 = n11988 & ~n13910;
  assign n13912 = ~n13909 & ~n13911;
  assign n13913 = n13907 & n13912;
  assign n13914 = ~n13902 & n13913;
  assign n13915 = ~n13899 & n13914;
  assign n13916 = n13897 & n13915;
  assign n13917 = n13008 & n13916;
  assign n13918 = ~n11997 & n13917;
  assign n13919 = n13918 ^ n10555;
  assign n13920 = n13919 ^ x540;
  assign n13921 = n13059 ^ x539;
  assign n13922 = n12925 ^ x542;
  assign n13923 = n10689 & n10692;
  assign n13924 = ~n10679 & n13281;
  assign n13925 = n10675 & ~n13924;
  assign n13926 = ~n13923 & ~n13925;
  assign n13927 = n10469 & n10699;
  assign n13928 = ~n10695 & ~n10698;
  assign n13929 = ~n10693 & ~n13928;
  assign n13930 = n10675 & n10687;
  assign n13931 = n10696 & n10702;
  assign n13932 = n12472 & n13931;
  assign n13933 = n10665 & ~n13932;
  assign n13934 = ~n13930 & ~n13933;
  assign n13935 = ~n10677 & ~n10683;
  assign n13936 = ~n10670 & n13935;
  assign n13937 = ~n10672 & n10706;
  assign n13938 = ~n10692 & n13937;
  assign n13939 = ~n13936 & ~n13938;
  assign n13940 = ~n10679 & ~n13939;
  assign n13941 = ~n10693 & ~n13940;
  assign n13942 = n13934 & ~n13941;
  assign n13943 = n12478 & n13942;
  assign n13944 = n12474 & n13943;
  assign n13945 = ~n13929 & n13944;
  assign n13946 = ~n13927 & n13945;
  assign n13947 = n13926 & n13946;
  assign n13948 = n13280 & n13947;
  assign n13949 = n13948 ^ n10576;
  assign n13950 = n13949 ^ x541;
  assign n13951 = ~n13922 & n13950;
  assign n13952 = n13921 & n13951;
  assign n13953 = ~n13920 & n13952;
  assign n13954 = n13894 & n13953;
  assign n13955 = n13892 & ~n13893;
  assign n13956 = n13920 & n13952;
  assign n13957 = n13921 & n13922;
  assign n13958 = n13920 & ~n13950;
  assign n13959 = n13957 & n13958;
  assign n13960 = ~n13956 & ~n13959;
  assign n13961 = n13955 & ~n13960;
  assign n13962 = ~n13954 & ~n13961;
  assign n13963 = ~n13892 & ~n13893;
  assign n13964 = ~n13920 & ~n13921;
  assign n13965 = n13922 & n13964;
  assign n13966 = ~n13950 & n13965;
  assign n13967 = n13950 & n13965;
  assign n13968 = n13920 & ~n13921;
  assign n13969 = n13951 & n13968;
  assign n13970 = ~n13967 & ~n13969;
  assign n13971 = ~n13966 & n13970;
  assign n13972 = n13963 & ~n13971;
  assign n13973 = ~n13920 & n13921;
  assign n13974 = ~n13922 & n13973;
  assign n13975 = ~n13950 & n13974;
  assign n13976 = ~n13921 & n13958;
  assign n13977 = n13922 & n13976;
  assign n13978 = ~n13975 & ~n13977;
  assign n13979 = n13955 & ~n13978;
  assign n13980 = ~n13972 & ~n13979;
  assign n13981 = n13962 & n13980;
  assign n13982 = n13920 & n13957;
  assign n13983 = n13950 & n13982;
  assign n13984 = n13894 & n13983;
  assign n13985 = n13922 & n13968;
  assign n13986 = n13950 & n13985;
  assign n13987 = n13955 & n13986;
  assign n13988 = ~n13984 & ~n13987;
  assign n13989 = ~n13920 & n13957;
  assign n13990 = n13950 & n13989;
  assign n13991 = n13894 & n13990;
  assign n13992 = ~n13922 & n13976;
  assign n13993 = n13955 & n13992;
  assign n13994 = ~n13991 & ~n13993;
  assign n13995 = n13988 & n13994;
  assign n13996 = n13951 & n13964;
  assign n13997 = n13955 & n13996;
  assign n13998 = n13894 & n13966;
  assign n13999 = n13892 & n13893;
  assign n14000 = ~n13950 & n13989;
  assign n14001 = n13999 & n14000;
  assign n14002 = ~n13998 & ~n14001;
  assign n14003 = ~n13997 & n14002;
  assign n14004 = ~n13922 & n13964;
  assign n14005 = ~n13950 & n14004;
  assign n14006 = n13894 & n14005;
  assign n14007 = ~n13971 & n13999;
  assign n14008 = ~n14006 & ~n14007;
  assign n14009 = ~n13959 & ~n13975;
  assign n14010 = ~n13956 & n14009;
  assign n14011 = n13963 & ~n14010;
  assign n14012 = n13921 & n13958;
  assign n14013 = ~n13922 & n14012;
  assign n14014 = ~n13996 & ~n14013;
  assign n14015 = n13893 & ~n14014;
  assign n14016 = ~n14011 & ~n14015;
  assign n14017 = n13893 ^ n13892;
  assign n14018 = n13990 ^ n13983;
  assign n14019 = n14018 ^ n13983;
  assign n14020 = n13983 ^ n13893;
  assign n14021 = n14020 ^ n13983;
  assign n14022 = n14019 & ~n14021;
  assign n14023 = n14022 ^ n13983;
  assign n14024 = n14017 & n14023;
  assign n14025 = n14024 ^ n13983;
  assign n14026 = n14016 & ~n14025;
  assign n14027 = n14008 & n14026;
  assign n14028 = n13977 ^ n13893;
  assign n14029 = n14028 ^ n13977;
  assign n14030 = n13977 ^ n13956;
  assign n14031 = n14030 ^ n13977;
  assign n14032 = n14029 & n14031;
  assign n14033 = n14032 ^ n13977;
  assign n14034 = n13892 & n14033;
  assign n14035 = n14034 ^ n13977;
  assign n14036 = n14027 & ~n14035;
  assign n14037 = n14003 & n14036;
  assign n14038 = n13995 & n14037;
  assign n14039 = n13981 & n14038;
  assign n14040 = n14039 ^ n10663;
  assign n14041 = n14040 ^ x551;
  assign n14042 = n12597 ^ x554;
  assign n14043 = n14041 & n14042;
  assign n14044 = n13891 & n14043;
  assign n14045 = n13864 & ~n13890;
  assign n14046 = n14041 & ~n14042;
  assign n14047 = n14045 & n14046;
  assign n14048 = ~n14044 & ~n14047;
  assign n14049 = n13003 ^ x555;
  assign n14050 = n13334 & n13343;
  assign n14051 = ~n13347 & n13602;
  assign n14052 = ~n14050 & ~n14051;
  assign n14053 = n13234 & n13344;
  assign n14054 = ~n13315 & ~n13348;
  assign n14055 = ~n13327 & n14054;
  assign n14056 = n13321 & ~n14055;
  assign n14057 = n13334 & ~n13596;
  assign n14058 = ~n13363 & n13612;
  assign n14059 = ~n14057 & ~n14058;
  assign n14060 = ~n13312 & ~n13343;
  assign n14061 = ~n13327 & n14060;
  assign n14062 = ~n13340 & n14061;
  assign n14063 = n13337 & n14062;
  assign n14064 = n13329 & ~n14063;
  assign n14065 = ~n13234 & n13341;
  assign n14066 = ~n13323 & ~n13361;
  assign n14067 = ~n13321 & n14066;
  assign n14068 = ~n14065 & ~n14067;
  assign n14069 = ~n13595 & ~n14068;
  assign n14070 = ~n13347 & ~n14069;
  assign n14071 = ~n14064 & ~n14070;
  assign n14072 = n14059 & n14071;
  assign n14073 = n13325 & n14072;
  assign n14074 = ~n14056 & n14073;
  assign n14075 = ~n14053 & n14074;
  assign n14076 = n14052 & n14075;
  assign n14077 = ~n13339 & n14076;
  assign n14078 = ~n13317 & n14077;
  assign n14079 = n14078 ^ n10278;
  assign n14080 = n14079 ^ x550;
  assign n14081 = ~n14049 & ~n14080;
  assign n14082 = ~n14048 & n14081;
  assign n14083 = n13864 & n13890;
  assign n14084 = ~n14041 & n14042;
  assign n14085 = n14083 & n14084;
  assign n14086 = ~n14041 & ~n14042;
  assign n14087 = n14045 & n14086;
  assign n14088 = ~n14085 & ~n14087;
  assign n14089 = n14049 & ~n14080;
  assign n14090 = ~n14088 & n14089;
  assign n14091 = ~n14082 & ~n14090;
  assign n14092 = n14046 & n14083;
  assign n14093 = n14089 & n14092;
  assign n14094 = n14083 & n14086;
  assign n14095 = n14081 & n14094;
  assign n14096 = ~n14093 & ~n14095;
  assign n14097 = ~n14049 & n14080;
  assign n14098 = ~n13864 & ~n13890;
  assign n14099 = n14086 & n14098;
  assign n14100 = ~n14085 & ~n14099;
  assign n14101 = n14097 & ~n14100;
  assign n14102 = n14087 & n14097;
  assign n14103 = n13891 & n14084;
  assign n14104 = n14089 & n14103;
  assign n14105 = ~n14102 & ~n14104;
  assign n14106 = ~n14101 & n14105;
  assign n14107 = n13891 & n14086;
  assign n14108 = n14049 & n14080;
  assign n14109 = n14107 & n14108;
  assign n14110 = n14046 & n14098;
  assign n14111 = n14089 & n14110;
  assign n14112 = ~n14109 & ~n14111;
  assign n14113 = n14043 & n14098;
  assign n14114 = ~n14092 & ~n14113;
  assign n14115 = n14081 & ~n14114;
  assign n14116 = n14043 & n14045;
  assign n14117 = ~n14044 & ~n14107;
  assign n14118 = ~n14116 & n14117;
  assign n14119 = n14089 & ~n14118;
  assign n14120 = ~n14115 & ~n14119;
  assign n14121 = n14097 & n14103;
  assign n14122 = n14080 ^ n14049;
  assign n14123 = n14084 & n14098;
  assign n14124 = n14045 & n14084;
  assign n14125 = ~n14099 & ~n14124;
  assign n14126 = ~n14123 & n14125;
  assign n14127 = ~n14122 & ~n14126;
  assign n14131 = n14048 & ~n14116;
  assign n14132 = ~n14092 & n14131;
  assign n14128 = n13890 ^ n13864;
  assign n14129 = n14128 ^ n14042;
  assign n14130 = n14041 & n14129;
  assign n14133 = n14132 ^ n14130;
  assign n14134 = n14130 ^ n14049;
  assign n14135 = n14134 ^ n14130;
  assign n14136 = ~n14133 & n14135;
  assign n14137 = n14136 ^ n14130;
  assign n14138 = n14080 & n14137;
  assign n14139 = ~n14127 & ~n14138;
  assign n14140 = ~n14121 & n14139;
  assign n14141 = n14120 & n14140;
  assign n14142 = n14112 & n14141;
  assign n14143 = n14106 & n14142;
  assign n14144 = n14096 & n14143;
  assign n14145 = n14091 & n14144;
  assign n14146 = n14145 ^ n12712;
  assign n14147 = n14146 ^ x611;
  assign n14148 = n13530 & n13544;
  assign n14149 = ~n13561 & ~n13868;
  assign n14150 = n13526 & ~n14149;
  assign n14151 = ~n14148 & ~n14150;
  assign n14152 = n13526 & n13572;
  assign n14153 = ~n13545 & n13559;
  assign n14154 = ~n14152 & ~n14153;
  assign n14155 = n13531 & ~n13542;
  assign n14156 = ~n13539 & ~n13578;
  assign n14157 = n13544 & ~n14156;
  assign n14158 = ~n13534 & ~n13561;
  assign n14159 = ~n13480 & n13528;
  assign n14160 = ~n13578 & ~n14159;
  assign n14161 = n14158 & n14160;
  assign n14162 = ~n13541 & n14161;
  assign n14163 = ~n13572 & n14162;
  assign n14164 = n13524 & ~n14163;
  assign n14165 = ~n13560 & ~n13581;
  assign n14166 = ~n13573 & n14165;
  assign n14167 = ~n13868 & n14166;
  assign n14168 = n13544 & ~n14167;
  assign n14169 = ~n13539 & n14160;
  assign n14170 = n13526 & ~n14169;
  assign n14171 = ~n13521 & n14165;
  assign n14172 = ~n13558 & n14171;
  assign n14173 = n13531 & ~n14172;
  assign n14174 = ~n14170 & ~n14173;
  assign n14175 = ~n14168 & n14174;
  assign n14176 = ~n14164 & n14175;
  assign n14177 = ~n13525 & n14176;
  assign n14178 = ~n14157 & n14177;
  assign n14179 = ~n14155 & n14178;
  assign n14180 = n14154 & n14179;
  assign n14181 = n14151 & n14180;
  assign n14182 = n13536 & n14181;
  assign n14183 = n14182 ^ n11276;
  assign n14184 = n14183 ^ x568;
  assign n14185 = ~n13986 & ~n13996;
  assign n14186 = n13999 & ~n14185;
  assign n14187 = n13955 & n13966;
  assign n14188 = ~n13953 & ~n13983;
  assign n14189 = ~n14005 & n14188;
  assign n14190 = n13963 & ~n14189;
  assign n14191 = ~n14187 & ~n14190;
  assign n14192 = n13955 & n13969;
  assign n14193 = n13894 & n13975;
  assign n14194 = ~n14192 & ~n14193;
  assign n14195 = n13992 & n13999;
  assign n14196 = n14194 & ~n14195;
  assign n14197 = n13955 & ~n14188;
  assign n14198 = ~n14000 & ~n14013;
  assign n14199 = ~n14017 & ~n14198;
  assign n14200 = ~n14197 & ~n14199;
  assign n14201 = n13894 & n13959;
  assign n14202 = ~n13894 & ~n13969;
  assign n14203 = ~n13986 & ~n13992;
  assign n14204 = ~n13977 & n14203;
  assign n14205 = ~n13999 & n14204;
  assign n14206 = ~n14202 & ~n14205;
  assign n14207 = ~n13990 & ~n14206;
  assign n14208 = ~n14005 & n14207;
  assign n14209 = n13893 & ~n14208;
  assign n14210 = ~n14201 & ~n14209;
  assign n14211 = n14200 & n14210;
  assign n14212 = n14196 & n14211;
  assign n14213 = n14191 & n14212;
  assign n14214 = n13981 & n14213;
  assign n14215 = ~n14186 & n14214;
  assign n14216 = n14215 ^ n10986;
  assign n14217 = n14216 ^ x573;
  assign n14218 = n14184 & n14217;
  assign n14219 = n12753 & ~n12772;
  assign n14220 = n12796 ^ n12765;
  assign n14221 = n14220 ^ n12796;
  assign n14222 = n12680 & ~n12753;
  assign n14223 = n14222 ^ n12796;
  assign n14224 = n14221 & n14223;
  assign n14225 = n14224 ^ n12796;
  assign n14226 = ~n14219 & ~n14225;
  assign n14227 = n12778 & n14226;
  assign n14228 = n12750 & n12771;
  assign n14229 = ~n12713 & n12796;
  assign n14230 = ~n12771 & ~n12780;
  assign n14231 = n12753 & ~n14230;
  assign n14232 = ~n14229 & ~n14231;
  assign n14233 = ~n14228 & n14232;
  assign n14234 = n12646 & ~n14233;
  assign n14235 = ~n14227 & ~n14234;
  assign n14236 = ~n12764 & n12779;
  assign n14237 = ~n12713 & n14222;
  assign n14238 = ~n12764 & ~n14237;
  assign n14239 = n14238 ^ n12680;
  assign n14240 = n14239 ^ n14238;
  assign n14241 = n14238 ^ n12713;
  assign n14242 = n14241 ^ n14238;
  assign n14243 = ~n14240 & ~n14242;
  assign n14244 = n14243 ^ n14238;
  assign n14245 = ~n12750 & ~n14244;
  assign n14246 = n14245 ^ n14238;
  assign n14247 = ~n14236 & n14246;
  assign n14248 = n14247 ^ n12644;
  assign n14249 = n14248 ^ n14247;
  assign n14250 = n12779 ^ n12680;
  assign n14251 = n14250 ^ n12779;
  assign n14252 = n12780 ^ n12779;
  assign n14253 = ~n14251 & ~n14252;
  assign n14254 = n14253 ^ n12779;
  assign n14255 = ~n12782 & ~n14254;
  assign n14256 = n12769 & ~n14255;
  assign n14257 = ~n12793 & n14256;
  assign n14258 = n14257 ^ n14247;
  assign n14259 = n14249 & n14258;
  assign n14260 = n14259 ^ n14247;
  assign n14261 = n12645 & ~n14260;
  assign n14262 = n14235 & ~n14261;
  assign n14263 = n14262 ^ n10776;
  assign n14264 = n14263 ^ x572;
  assign n14265 = n13321 & n13340;
  assign n14266 = n13234 & ~n13596;
  assign n14267 = ~n14265 & ~n14266;
  assign n14268 = n13329 & n13595;
  assign n14269 = ~n13336 & n13369;
  assign n14270 = n13612 & ~n14269;
  assign n14271 = ~n14268 & ~n14270;
  assign n14272 = ~n13361 & n14061;
  assign n14273 = n13334 & ~n14272;
  assign n14274 = ~n13348 & ~n13602;
  assign n14275 = ~n13321 & n14274;
  assign n14276 = ~n13343 & ~n13362;
  assign n14277 = ~n13234 & n14276;
  assign n14278 = ~n14275 & ~n14277;
  assign n14279 = n13331 & ~n14278;
  assign n14280 = ~n13347 & ~n14279;
  assign n14281 = ~n14273 & ~n14280;
  assign n14282 = n14271 & n14281;
  assign n14283 = n14267 & n14282;
  assign n14284 = n13598 & n14283;
  assign n14285 = ~n13632 & n14284;
  assign n14286 = n13333 & n14285;
  assign n14287 = n13325 & n14286;
  assign n14288 = n14287 ^ n11316;
  assign n14289 = n14288 ^ x571;
  assign n14290 = n14264 & n14289;
  assign n14291 = ~n12029 & ~n12073;
  assign n14292 = n11230 & ~n14291;
  assign n14293 = ~n12024 & ~n12069;
  assign n14294 = n12042 & ~n14293;
  assign n14295 = ~n12033 & ~n12073;
  assign n14296 = ~n12068 & ~n14295;
  assign n14297 = ~n12047 & n12066;
  assign n14298 = n12053 & ~n14297;
  assign n14299 = n12039 & n12079;
  assign n14300 = n12042 & ~n14299;
  assign n14301 = ~n14298 & ~n14300;
  assign n14302 = ~n14296 & n14301;
  assign n14303 = n12026 & ~n12045;
  assign n14304 = ~n12043 & n13732;
  assign n14305 = ~n12038 & n14304;
  assign n14306 = ~n12033 & n14305;
  assign n14307 = n11230 & ~n14306;
  assign n14308 = ~n14303 & ~n14307;
  assign n14309 = n14302 & n14308;
  assign n14310 = ~n13722 & n14309;
  assign n14311 = ~n14294 & n14310;
  assign n14312 = n12031 & n14311;
  assign n14313 = n12050 & n14312;
  assign n14314 = ~n14292 & n14313;
  assign n14315 = ~n13717 & n14314;
  assign n14316 = n14315 ^ n11399;
  assign n14317 = n14316 ^ x570;
  assign n14318 = ~n12927 & n12931;
  assign n14319 = ~n12908 & ~n12983;
  assign n14320 = ~n12963 & n14319;
  assign n14321 = n12961 & ~n14320;
  assign n14322 = ~n14318 & ~n14321;
  assign n14323 = ~n12973 & n12986;
  assign n14324 = ~n12953 & ~n12975;
  assign n14325 = ~n12933 & n14324;
  assign n14326 = ~n12928 & ~n12963;
  assign n14327 = n13659 & n14326;
  assign n14328 = ~n12971 & n14327;
  assign n14329 = ~n14325 & ~n14328;
  assign n14330 = ~n12978 & ~n14329;
  assign n14331 = n14330 ^ n12927;
  assign n14332 = n14331 ^ n14330;
  assign n14333 = ~n12935 & ~n12939;
  assign n14334 = n14333 ^ n14330;
  assign n14335 = n14334 ^ n14330;
  assign n14336 = n14332 & ~n14335;
  assign n14337 = n14336 ^ n14330;
  assign n14338 = ~n12926 & ~n14337;
  assign n14339 = n14338 ^ n14330;
  assign n14340 = ~n14323 & n14339;
  assign n14341 = n14322 & n14340;
  assign n14342 = n12965 & n14341;
  assign n14343 = ~n13665 & n14342;
  assign n14344 = n13661 & n14343;
  assign n14345 = n12952 & n14344;
  assign n14346 = ~n13675 & n14345;
  assign n14347 = n12937 & n14346;
  assign n14348 = n14347 ^ n11354;
  assign n14349 = n14348 ^ x569;
  assign n14350 = ~n14317 & n14349;
  assign n14351 = n14290 & n14350;
  assign n14352 = n14218 & n14351;
  assign n14353 = ~n14184 & ~n14217;
  assign n14354 = n14351 & n14353;
  assign n14355 = n14184 & ~n14217;
  assign n14356 = ~n14264 & n14289;
  assign n14357 = ~n14317 & ~n14349;
  assign n14358 = n14356 & n14357;
  assign n14359 = n14355 & n14358;
  assign n14360 = ~n14354 & ~n14359;
  assign n14361 = n14317 & ~n14349;
  assign n14362 = n14290 & n14361;
  assign n14363 = n14355 & n14362;
  assign n14364 = n14264 & ~n14289;
  assign n14365 = n14350 & n14364;
  assign n14366 = n14218 & n14365;
  assign n14367 = n14361 & n14364;
  assign n14368 = n14353 & n14367;
  assign n14369 = ~n14366 & ~n14368;
  assign n14370 = ~n14363 & n14369;
  assign n14371 = n14290 & n14357;
  assign n14372 = n14353 & n14371;
  assign n14373 = n14217 ^ n14184;
  assign n14374 = n14357 & n14364;
  assign n14375 = ~n14264 & ~n14289;
  assign n14376 = n14361 & n14375;
  assign n14377 = ~n14374 & ~n14376;
  assign n14378 = n14373 & ~n14377;
  assign n14379 = ~n14372 & ~n14378;
  assign n14380 = n14356 & n14361;
  assign n14381 = ~n14184 & n14380;
  assign n14382 = ~n14184 & n14217;
  assign n14383 = n14357 & n14375;
  assign n14384 = n14382 & n14383;
  assign n14385 = ~n14381 & ~n14384;
  assign n14386 = n14317 & n14349;
  assign n14387 = n14375 & n14386;
  assign n14388 = n14290 & n14386;
  assign n14389 = ~n14387 & ~n14388;
  assign n14390 = n14350 & n14375;
  assign n14391 = ~n14365 & ~n14390;
  assign n14392 = n14389 & n14391;
  assign n14393 = n14353 & ~n14392;
  assign n14394 = n14350 & n14356;
  assign n14395 = n14364 & n14386;
  assign n14396 = ~n14390 & ~n14395;
  assign n14397 = ~n14394 & n14396;
  assign n14398 = ~n14388 & n14397;
  assign n14399 = n14355 & ~n14398;
  assign n14400 = n14356 & n14386;
  assign n14401 = ~n14395 & ~n14400;
  assign n14402 = ~n14394 & n14401;
  assign n14403 = ~n14351 & n14402;
  assign n14404 = n14382 & ~n14403;
  assign n14405 = ~n14399 & ~n14404;
  assign n14406 = ~n14393 & n14405;
  assign n14410 = ~n14367 & ~n14387;
  assign n14407 = ~n14371 & ~n14380;
  assign n14408 = ~n14362 & n14407;
  assign n14409 = ~n14383 & n14408;
  assign n14411 = n14410 ^ n14409;
  assign n14412 = n14410 ^ n14218;
  assign n14413 = n14410 & n14412;
  assign n14414 = n14413 ^ n14410;
  assign n14415 = n14411 & n14414;
  assign n14416 = n14415 ^ n14413;
  assign n14417 = n14416 ^ n14410;
  assign n14418 = n14417 ^ n14218;
  assign n14419 = n14406 & n14418;
  assign n14420 = n14419 ^ n14406;
  assign n14421 = n14385 & n14420;
  assign n14422 = n14379 & n14421;
  assign n14423 = n14370 & n14422;
  assign n14424 = n14360 & n14423;
  assign n14425 = ~n14352 & n14424;
  assign n14426 = n14425 ^ n12749;
  assign n14427 = n14426 ^ x612;
  assign n14428 = ~n14147 & n14427;
  assign n14429 = ~n13825 & n14428;
  assign n14430 = n13825 & n14427;
  assign n14431 = n14147 & n14430;
  assign n14432 = ~n14429 & ~n14431;
  assign n14433 = ~n13461 & ~n14432;
  assign n14434 = n13542 & ~n13581;
  assign n14435 = ~n13558 & n14434;
  assign n14436 = n13526 & ~n14435;
  assign n14437 = n13563 & ~n13868;
  assign n14438 = n13524 & ~n14437;
  assign n14439 = ~n14436 & ~n14438;
  assign n14441 = ~n13581 & n14158;
  assign n14440 = ~n13560 & n13582;
  assign n14442 = n14441 ^ n14440;
  assign n14443 = n14440 ^ n13523;
  assign n14444 = ~n13569 & n14443;
  assign n14445 = n14444 ^ n13523;
  assign n14446 = n14442 & n14445;
  assign n14447 = n14446 ^ n14441;
  assign n14448 = ~n13879 & n14447;
  assign n14449 = n13869 & n14448;
  assign n14450 = ~n13545 & ~n14449;
  assign n14451 = n14439 & ~n14450;
  assign n14452 = n14151 & n14451;
  assign n14453 = n13867 & n14452;
  assign n14454 = n13537 & n14453;
  assign n14455 = ~n13525 & n14454;
  assign n14456 = n14455 ^ n11108;
  assign n14457 = n14456 ^ x580;
  assign n14458 = n13635 ^ x585;
  assign n14459 = ~n14457 & n14458;
  assign n14460 = n14457 & ~n14458;
  assign n14461 = ~n14459 & ~n14460;
  assign n14462 = n12646 & ~n14247;
  assign n14463 = n12792 & ~n14226;
  assign n14464 = ~n14462 & ~n14463;
  assign n14465 = n12778 & ~n14257;
  assign n14466 = n12763 & n14233;
  assign n14467 = ~n14465 & ~n14466;
  assign n14468 = n14464 & n14467;
  assign n14469 = n14468 ^ n11516;
  assign n14470 = n14469 ^ x582;
  assign n14471 = n12524 & n12530;
  assign n14472 = n12526 & n12532;
  assign n14473 = ~n14471 & ~n14472;
  assign n14474 = n12530 & n12567;
  assign n14475 = ~n12566 & ~n12581;
  assign n14476 = ~n12574 & ~n12584;
  assign n14477 = ~n12547 & n14476;
  assign n14478 = ~n12565 & n14477;
  assign n14479 = n14475 & n14478;
  assign n14480 = ~n12552 & n14479;
  assign n14481 = n12175 & ~n14480;
  assign n14482 = ~n14474 & ~n14481;
  assign n14483 = ~n12549 & ~n12562;
  assign n14484 = n12542 & ~n14483;
  assign n14485 = n12470 ^ n12295;
  assign n14486 = n14485 ^ n12470;
  assign n14487 = n12470 ^ n12418;
  assign n14488 = n14487 ^ n12470;
  assign n14489 = ~n14486 & n14488;
  assign n14490 = n14489 ^ n12470;
  assign n14491 = n12522 & n14490;
  assign n14492 = n12568 & ~n14491;
  assign n14493 = n12526 & ~n14492;
  assign n14494 = n12581 ^ n12137;
  assign n14496 = ~n12573 & ~n12584;
  assign n14497 = ~n12564 & n14496;
  assign n14495 = ~n12552 & n12586;
  assign n14498 = n14497 ^ n14495;
  assign n14499 = n14497 ^ n12174;
  assign n14500 = n14499 ^ n14497;
  assign n14501 = n14498 & ~n14500;
  assign n14502 = n14501 ^ n14497;
  assign n14503 = n14502 ^ n12581;
  assign n14504 = n14494 & ~n14503;
  assign n14505 = n14504 ^ n14501;
  assign n14506 = n14505 ^ n14497;
  assign n14507 = n14506 ^ n12137;
  assign n14508 = ~n12581 & ~n14507;
  assign n14509 = n14508 ^ n12581;
  assign n14510 = n14509 ^ n12137;
  assign n14511 = ~n14493 & ~n14510;
  assign n14512 = ~n14484 & n14511;
  assign n14513 = n14482 & n14512;
  assign n14514 = n12539 & n14513;
  assign n14515 = n12544 & n14514;
  assign n14516 = n14473 & n14515;
  assign n14517 = n14516 ^ n10819;
  assign n14518 = n14517 ^ x581;
  assign n14519 = n14470 & n14518;
  assign n14520 = n13894 & n13969;
  assign n14521 = n13975 & ~n14017;
  assign n14522 = ~n14520 & ~n14521;
  assign n14523 = n13955 & ~n14198;
  assign n14524 = ~n13959 & ~n13967;
  assign n14525 = n13893 & ~n14524;
  assign n14526 = ~n13967 & ~n13992;
  assign n14527 = ~n13990 & n14526;
  assign n14528 = n13963 & ~n14527;
  assign n14529 = ~n14525 & ~n14528;
  assign n14530 = ~n14523 & n14529;
  assign n14531 = n14522 & n14530;
  assign n14532 = ~n14035 & n14531;
  assign n14533 = n13988 & n14532;
  assign n14534 = n14003 & n14533;
  assign n14535 = n14196 & n14534;
  assign n14536 = n13962 & n14535;
  assign n14537 = n14191 & n14536;
  assign n14538 = ~n14186 & n14537;
  assign n14539 = n14538 ^ n11571;
  assign n14540 = n14539 ^ x583;
  assign n14541 = n13749 ^ x584;
  assign n14542 = ~n14540 & ~n14541;
  assign n14543 = n14519 & n14542;
  assign n14544 = n14461 & n14543;
  assign n14545 = n14457 & n14458;
  assign n14546 = ~n14470 & n14518;
  assign n14547 = n14541 & n14546;
  assign n14548 = ~n14540 & n14547;
  assign n14549 = n14540 & ~n14541;
  assign n14550 = n14546 & n14549;
  assign n14551 = n14519 & n14549;
  assign n14552 = ~n14550 & ~n14551;
  assign n14553 = ~n14548 & n14552;
  assign n14554 = n14545 & ~n14553;
  assign n14555 = ~n14470 & ~n14518;
  assign n14556 = n14540 & n14541;
  assign n14557 = n14555 & n14556;
  assign n14558 = n14542 & n14546;
  assign n14559 = ~n14540 & n14541;
  assign n14560 = n14519 & n14559;
  assign n14561 = ~n14550 & ~n14560;
  assign n14562 = ~n14558 & n14561;
  assign n14563 = ~n14557 & n14562;
  assign n14564 = n14459 & ~n14563;
  assign n14565 = ~n14551 & ~n14560;
  assign n14566 = ~n14548 & n14565;
  assign n14567 = n14549 & n14555;
  assign n14568 = n14470 & ~n14518;
  assign n14569 = n14559 & n14568;
  assign n14570 = n14556 & n14568;
  assign n14571 = n14542 & n14555;
  assign n14572 = ~n14570 & ~n14571;
  assign n14573 = ~n14569 & n14572;
  assign n14574 = ~n14567 & n14573;
  assign n14575 = n14566 & n14574;
  assign n14576 = ~n14557 & n14575;
  assign n14577 = n14460 & n14576;
  assign n14578 = ~n14564 & ~n14577;
  assign n14579 = ~n14457 & ~n14458;
  assign n14580 = n14540 & n14547;
  assign n14581 = ~n14551 & ~n14580;
  assign n14582 = ~n14548 & n14581;
  assign n14583 = n14579 & ~n14582;
  assign n14584 = n14549 & n14568;
  assign n14585 = n14555 & n14559;
  assign n14586 = ~n14567 & ~n14585;
  assign n14587 = ~n14584 & n14586;
  assign n14588 = ~n14569 & n14587;
  assign n14589 = n14588 ^ n14458;
  assign n14590 = n14589 ^ n14588;
  assign n14591 = n14588 ^ n14574;
  assign n14592 = n14591 ^ n14588;
  assign n14593 = n14590 & ~n14592;
  assign n14594 = n14593 ^ n14588;
  assign n14595 = n14457 & ~n14594;
  assign n14596 = n14595 ^ n14588;
  assign n14597 = ~n14583 & n14596;
  assign n14598 = n14578 & n14597;
  assign n14599 = ~n14554 & n14598;
  assign n14600 = ~n14544 & n14599;
  assign n14601 = n14600 ^ n12643;
  assign n14602 = n14601 ^ x610;
  assign n14603 = n13655 ^ x544;
  assign n14604 = n14040 ^ x549;
  assign n14605 = n14603 & n14604;
  assign n14606 = ~n12552 & n12575;
  assign n14607 = n12175 & ~n14606;
  assign n14608 = n12577 & n14477;
  assign n14609 = ~n12564 & n14608;
  assign n14610 = n12526 & ~n14609;
  assign n14611 = n12577 & n14475;
  assign n14612 = ~n12584 & n14611;
  assign n14613 = n12542 & ~n14612;
  assign n14614 = ~n14610 & ~n14613;
  assign n14615 = ~n12137 & n12573;
  assign n14616 = ~n12532 & n12569;
  assign n14617 = n12530 & ~n14616;
  assign n14618 = ~n12528 & n12570;
  assign n14619 = n12175 & ~n14618;
  assign n14620 = ~n14617 & ~n14619;
  assign n14621 = ~n14615 & n14620;
  assign n14622 = n14614 & n14621;
  assign n14623 = ~n14607 & n14622;
  assign n14624 = n12561 & n14623;
  assign n14625 = n14473 & n14624;
  assign n14626 = n14625 ^ n10085;
  assign n14627 = n14626 ^ x547;
  assign n14628 = n12053 & ~n14295;
  assign n14629 = n12045 & ~n13715;
  assign n14630 = ~n12020 & ~n12043;
  assign n14631 = ~n12053 & n14630;
  assign n14632 = ~n14629 & ~n14631;
  assign n14633 = n13719 & ~n14632;
  assign n14634 = n14633 ^ n11229;
  assign n14635 = n14634 ^ n14633;
  assign n14636 = ~n12029 & n13732;
  assign n14637 = n14636 ^ n14633;
  assign n14638 = n14637 ^ n14633;
  assign n14639 = n14635 & ~n14638;
  assign n14640 = n14639 ^ n14633;
  assign n14641 = n12068 & ~n14640;
  assign n14642 = n14641 ^ n14633;
  assign n14643 = ~n14628 & n14642;
  assign n14644 = ~n12074 & ~n12078;
  assign n14645 = n14644 ^ n10736;
  assign n14646 = n14645 ^ n14644;
  assign n14647 = ~n12037 & ~n12064;
  assign n14648 = n14647 ^ n14644;
  assign n14649 = n14648 ^ n14644;
  assign n14650 = n14646 & ~n14649;
  assign n14651 = n14650 ^ n14644;
  assign n14652 = n11229 & ~n14651;
  assign n14653 = n14652 ^ n14644;
  assign n14654 = n14643 & n14653;
  assign n14655 = ~n14294 & n14654;
  assign n14656 = ~n12052 & n14655;
  assign n14657 = ~n14292 & n14656;
  assign n14658 = n12032 & n14657;
  assign n14659 = n13724 & n14658;
  assign n14660 = n14659 ^ n9765;
  assign n14661 = n14660 ^ x546;
  assign n14662 = ~n14627 & n14661;
  assign n14663 = n13713 ^ x545;
  assign n14664 = n14079 ^ x548;
  assign n14665 = ~n14663 & ~n14664;
  assign n14666 = n14662 & n14665;
  assign n14667 = n14605 & n14666;
  assign n14668 = ~n14603 & n14604;
  assign n14669 = ~n14663 & n14664;
  assign n14670 = n14662 & n14669;
  assign n14671 = n14668 & n14670;
  assign n14672 = n14603 & ~n14604;
  assign n14673 = n14627 & ~n14661;
  assign n14674 = n14669 & n14673;
  assign n14675 = ~n14666 & ~n14674;
  assign n14676 = n14672 & ~n14675;
  assign n14677 = ~n14671 & ~n14676;
  assign n14678 = ~n14603 & ~n14604;
  assign n14679 = ~n14627 & ~n14661;
  assign n14680 = n14669 & n14679;
  assign n14681 = ~n14666 & ~n14680;
  assign n14682 = n14678 & ~n14681;
  assign n14683 = n14627 & n14661;
  assign n14684 = n14669 & n14683;
  assign n14685 = n14665 & n14679;
  assign n14686 = ~n14684 & ~n14685;
  assign n14687 = n14605 & ~n14686;
  assign n14688 = n14665 & n14683;
  assign n14689 = ~n14670 & ~n14688;
  assign n14690 = n14678 & ~n14689;
  assign n14691 = ~n14687 & ~n14690;
  assign n14692 = n14663 & n14664;
  assign n14693 = n14662 & n14692;
  assign n14694 = n14663 & ~n14664;
  assign n14695 = n14683 & n14694;
  assign n14696 = ~n14693 & ~n14695;
  assign n14697 = n14683 & n14692;
  assign n14698 = n14679 & n14694;
  assign n14699 = ~n14697 & ~n14698;
  assign n14700 = n14696 & n14699;
  assign n14701 = ~n14670 & n14700;
  assign n14702 = n14672 & ~n14701;
  assign n14703 = n14673 & n14692;
  assign n14704 = n14662 & n14694;
  assign n14705 = n14673 & n14694;
  assign n14706 = ~n14704 & ~n14705;
  assign n14707 = ~n14605 & n14706;
  assign n14708 = ~n14697 & n14707;
  assign n14709 = ~n14703 & n14708;
  assign n14710 = ~n14695 & n14699;
  assign n14711 = ~n14703 & n14710;
  assign n14712 = n14605 & ~n14711;
  assign n14713 = ~n14678 & ~n14712;
  assign n14714 = ~n14709 & ~n14713;
  assign n14715 = ~n14702 & ~n14714;
  assign n14716 = n14680 ^ n14604;
  assign n14717 = n14716 ^ n14680;
  assign n14718 = n14679 & n14692;
  assign n14719 = n14665 & n14673;
  assign n14720 = ~n14684 & ~n14719;
  assign n14721 = ~n14718 & n14720;
  assign n14722 = n14696 & n14721;
  assign n14723 = n14706 & n14722;
  assign n14724 = n14723 ^ n14680;
  assign n14725 = n14724 ^ n14680;
  assign n14726 = n14717 & ~n14725;
  assign n14727 = n14726 ^ n14680;
  assign n14728 = ~n14603 & n14727;
  assign n14729 = n14728 ^ n14680;
  assign n14730 = n14715 & ~n14729;
  assign n14731 = n14691 & n14730;
  assign n14732 = ~n14682 & n14731;
  assign n14733 = n14677 & n14732;
  assign n14734 = ~n14667 & n14733;
  assign n14735 = n14734 ^ n12521;
  assign n14736 = n14735 ^ x615;
  assign n14737 = ~n14602 & n14736;
  assign n14738 = n14427 ^ n13461;
  assign n14739 = ~n14147 & ~n14738;
  assign n14740 = n13461 & n14430;
  assign n14741 = ~n14739 & ~n14740;
  assign n14742 = n13461 & n13825;
  assign n14743 = n14742 ^ n13825;
  assign n14744 = n14743 ^ n14742;
  assign n14745 = n14742 ^ n14738;
  assign n14746 = n14745 ^ n14742;
  assign n14747 = ~n14744 & n14746;
  assign n14748 = n14747 ^ n14742;
  assign n14749 = n14147 & n14748;
  assign n14750 = n14749 ^ n14742;
  assign n14751 = n14741 & ~n14750;
  assign n14752 = n14737 & n14751;
  assign n14753 = n14602 & n14736;
  assign n14754 = ~n13461 & ~n14427;
  assign n14755 = n13825 & n14754;
  assign n14756 = n14755 ^ n14430;
  assign n14757 = ~n14147 & n14756;
  assign n14758 = n14757 ^ n14430;
  assign n14759 = ~n14750 & ~n14758;
  assign n14760 = ~n14433 & n14759;
  assign n14761 = n14753 & ~n14760;
  assign n14762 = ~n14752 & ~n14761;
  assign n14763 = ~n14602 & ~n14736;
  assign n14764 = ~n13825 & n14147;
  assign n14765 = ~n14428 & ~n14764;
  assign n14766 = n13461 & ~n14765;
  assign n14767 = ~n14755 & ~n14766;
  assign n14768 = n14763 & ~n14767;
  assign n14769 = n14602 & ~n14736;
  assign n14770 = n14147 ^ n13461;
  assign n14771 = n14770 ^ n14427;
  assign n14772 = n14738 ^ n13461;
  assign n14773 = n13825 ^ n13461;
  assign n14774 = ~n14772 & ~n14773;
  assign n14775 = n14774 ^ n13461;
  assign n14776 = ~n14771 & n14775;
  assign n14777 = n14776 ^ n13461;
  assign n14778 = n14769 & n14777;
  assign n14779 = ~n14768 & ~n14778;
  assign n14780 = n14762 & n14779;
  assign n14781 = ~n14433 & n14780;
  assign n14782 = n14781 ^ n13713;
  assign n14783 = n14782 ^ x687;
  assign n14784 = n14668 & n14697;
  assign n14785 = n14696 & ~n14705;
  assign n14786 = n14678 & ~n14785;
  assign n14787 = ~n14784 & ~n14786;
  assign n14788 = ~n14667 & n14787;
  assign n14789 = ~n14674 & ~n14688;
  assign n14790 = ~n14698 & n14789;
  assign n14791 = n14678 & ~n14790;
  assign n14792 = n14686 & ~n14703;
  assign n14793 = n14668 & ~n14792;
  assign n14794 = ~n14791 & ~n14793;
  assign n14795 = n14722 ^ n14604;
  assign n14796 = n14795 ^ n14722;
  assign n14797 = n14689 & n14699;
  assign n14798 = ~n14680 & n14797;
  assign n14799 = ~n14705 & n14798;
  assign n14800 = n14799 ^ n14722;
  assign n14801 = n14796 & n14800;
  assign n14802 = n14801 ^ n14722;
  assign n14803 = n14603 & ~n14802;
  assign n14804 = n14794 & ~n14803;
  assign n14805 = n14677 & n14804;
  assign n14806 = n14680 ^ n14668;
  assign n14807 = n14680 ^ n14678;
  assign n14808 = n14807 ^ n14678;
  assign n14809 = n14719 ^ n14678;
  assign n14810 = ~n14808 & ~n14809;
  assign n14811 = n14810 ^ n14678;
  assign n14812 = n14806 & n14811;
  assign n14813 = n14812 ^ n14668;
  assign n14814 = n14805 & ~n14813;
  assign n14815 = n14788 & n14814;
  assign n14816 = ~n14704 & n14815;
  assign n14817 = n14816 ^ n10735;
  assign n14818 = n14817 ^ x603;
  assign n14819 = n14263 ^ x574;
  assign n14820 = n14517 ^ x579;
  assign n14821 = n14819 & n14820;
  assign n14822 = n13037 & n13190;
  assign n14823 = ~n13185 & n13838;
  assign n14824 = n13221 & n14823;
  assign n14825 = ~n13216 & n14824;
  assign n14826 = n13192 & ~n14825;
  assign n14827 = ~n14822 & ~n14826;
  assign n14828 = ~n13187 & n13217;
  assign n14829 = n13205 & ~n14828;
  assign n14830 = ~n13648 & n13854;
  assign n14831 = n13061 & ~n14830;
  assign n14832 = ~n14829 & ~n14831;
  assign n14833 = ~n13193 & n13850;
  assign n14834 = n13177 & ~n14833;
  assign n14835 = ~n13170 & ~n13205;
  assign n14836 = n13171 & n13177;
  assign n14837 = n13202 & ~n14836;
  assign n14838 = ~n13179 & n14837;
  assign n14839 = ~n13193 & n14838;
  assign n14840 = ~n14835 & ~n14839;
  assign n14841 = n13640 & n14840;
  assign n14842 = ~n14834 & ~n14841;
  assign n14843 = n14832 & n14842;
  assign n14844 = n14827 & n14843;
  assign n14845 = n13197 & n14844;
  assign n14846 = n13183 & n14845;
  assign n14847 = n14846 ^ n11149;
  assign n14848 = n14847 ^ x576;
  assign n14849 = n14216 ^ x575;
  assign n14850 = n14848 & n14849;
  assign n14851 = n14456 ^ x578;
  assign n14852 = n12908 & ~n12927;
  assign n14853 = n12958 & n12961;
  assign n14854 = ~n14852 & ~n14853;
  assign n14855 = ~n12975 & n13672;
  assign n14856 = n12933 & ~n14855;
  assign n14857 = n12980 & n13659;
  assign n14858 = ~n12947 & n14857;
  assign n14859 = ~n12931 & n14858;
  assign n14860 = n12944 & ~n14859;
  assign n14861 = ~n14856 & ~n14860;
  assign n14862 = ~n12961 & ~n12983;
  assign n14863 = ~n12975 & n14326;
  assign n14864 = ~n14862 & ~n14863;
  assign n14865 = ~n12953 & ~n14864;
  assign n14866 = ~n12971 & n14865;
  assign n14867 = ~n12973 & ~n14866;
  assign n14868 = n14861 & ~n14867;
  assign n14869 = n14854 & n14868;
  assign n14870 = ~n13658 & n14869;
  assign n14871 = ~n13693 & n14870;
  assign n14872 = n13663 & n14871;
  assign n14873 = ~n13675 & n14872;
  assign n14874 = ~n12940 & n14873;
  assign n14875 = n12937 & n14874;
  assign n14876 = n14875 ^ n10950;
  assign n14877 = n14876 ^ x577;
  assign n14878 = n14851 & ~n14877;
  assign n14879 = n14850 & n14878;
  assign n14880 = n14821 & n14879;
  assign n14881 = ~n14819 & ~n14820;
  assign n14882 = ~n14848 & n14849;
  assign n14883 = ~n14851 & ~n14877;
  assign n14884 = n14882 & n14883;
  assign n14885 = n14881 & n14884;
  assign n14886 = n14848 & ~n14849;
  assign n14887 = n14878 & n14886;
  assign n14888 = ~n14819 & n14820;
  assign n14889 = n14819 & ~n14820;
  assign n14890 = ~n14888 & ~n14889;
  assign n14891 = n14887 & ~n14890;
  assign n14892 = ~n14885 & ~n14891;
  assign n14893 = ~n14880 & n14892;
  assign n14894 = n14851 & n14877;
  assign n14895 = ~n14848 & ~n14849;
  assign n14896 = n14894 & n14895;
  assign n14897 = n14883 & n14895;
  assign n14898 = ~n14896 & ~n14897;
  assign n14899 = n14881 & ~n14898;
  assign n14900 = n14850 & n14883;
  assign n14901 = n14900 ^ n14820;
  assign n14902 = n14901 ^ n14900;
  assign n14903 = n14900 ^ n14884;
  assign n14904 = n14902 & n14903;
  assign n14905 = n14904 ^ n14900;
  assign n14906 = n14819 & n14905;
  assign n14907 = ~n14899 & ~n14906;
  assign n14908 = n14878 & n14882;
  assign n14909 = n14889 & n14908;
  assign n14910 = n14886 & n14894;
  assign n14911 = n14821 & n14910;
  assign n14912 = ~n14909 & ~n14911;
  assign n14913 = n14883 & n14886;
  assign n14914 = n14888 & n14913;
  assign n14915 = ~n14851 & n14877;
  assign n14916 = n14850 & n14915;
  assign n14917 = n14882 & n14894;
  assign n14918 = ~n14916 & ~n14917;
  assign n14919 = ~n14910 & n14918;
  assign n14920 = ~n14879 & n14919;
  assign n14921 = ~n14900 & n14920;
  assign n14922 = n14881 & ~n14921;
  assign n14923 = n14886 & n14915;
  assign n14924 = n14820 & n14923;
  assign n14925 = ~n14890 & n14916;
  assign n14926 = ~n14924 & ~n14925;
  assign n14927 = n14882 & n14915;
  assign n14928 = n14850 & n14894;
  assign n14929 = ~n14927 & ~n14928;
  assign n14930 = ~n14888 & n14929;
  assign n14931 = ~n14890 & ~n14930;
  assign n14932 = ~n14908 & ~n14928;
  assign n14933 = ~n14884 & n14932;
  assign n14934 = ~n14889 & n14933;
  assign n14935 = n14931 & ~n14934;
  assign n14936 = n14898 & ~n14927;
  assign n14937 = ~n14900 & n14936;
  assign n14938 = n14821 & ~n14937;
  assign n14939 = ~n14935 & ~n14938;
  assign n14940 = n14926 & n14939;
  assign n14941 = ~n14922 & n14940;
  assign n14942 = ~n14914 & n14941;
  assign n14943 = n14878 & n14895;
  assign n14944 = n14943 ^ n14889;
  assign n14945 = n14943 ^ n14888;
  assign n14946 = n14945 ^ n14888;
  assign n14947 = n14895 & n14915;
  assign n14948 = n14947 ^ n14888;
  assign n14949 = ~n14946 & ~n14948;
  assign n14950 = n14949 ^ n14888;
  assign n14951 = n14944 & n14950;
  assign n14952 = n14951 ^ n14889;
  assign n14953 = n14942 & ~n14952;
  assign n14954 = n14912 & n14953;
  assign n14955 = n14907 & n14954;
  assign n14956 = n14893 & n14955;
  assign n14957 = n14956 ^ n11228;
  assign n14958 = n14957 ^ x598;
  assign n14959 = n14818 & ~n14958;
  assign n14960 = ~n13398 & ~n13434;
  assign n14961 = ~n13402 & ~n13451;
  assign n14962 = ~n14960 & ~n14961;
  assign n14963 = ~n13412 & ~n13424;
  assign n14964 = n14963 ^ n12598;
  assign n14965 = n14964 ^ n14963;
  assign n14966 = n14963 ^ n13420;
  assign n14967 = n14965 & n14966;
  assign n14968 = n14967 ^ n14963;
  assign n14969 = ~n13448 & ~n14968;
  assign n14970 = ~n14962 & ~n14969;
  assign n14971 = n13414 & n13448;
  assign n14972 = ~n13387 & ~n13401;
  assign n14973 = n13434 & ~n14972;
  assign n14974 = ~n13411 & ~n14973;
  assign n14975 = ~n13385 & ~n13424;
  assign n14976 = n13393 & ~n14975;
  assign n14977 = ~n13402 & n14963;
  assign n14978 = ~n13389 & n14977;
  assign n14979 = n12599 & ~n14978;
  assign n14980 = ~n14976 & ~n14979;
  assign n14981 = ~n13406 & n14960;
  assign n14982 = ~n13410 & ~n13425;
  assign n14983 = n13434 & ~n14982;
  assign n14984 = ~n13395 & ~n13419;
  assign n14985 = ~n13385 & n14984;
  assign n14986 = ~n13404 & n14985;
  assign n14987 = n13398 & ~n14986;
  assign n14988 = ~n14983 & ~n14987;
  assign n14989 = ~n14981 & n14988;
  assign n14990 = n14980 & n14989;
  assign n14991 = ~n13397 & n14990;
  assign n14992 = n14974 & n14991;
  assign n14993 = ~n14971 & n14992;
  assign n14994 = n14970 & n14993;
  assign n14995 = ~n13413 & n14994;
  assign n14996 = n14995 ^ n12017;
  assign n14997 = n14996 ^ x600;
  assign n14998 = ~n14358 & ~n14374;
  assign n14999 = n14382 & ~n14998;
  assign n15000 = ~n14380 & ~n14383;
  assign n15001 = n14353 & ~n15000;
  assign n15002 = n14218 & n14400;
  assign n15003 = n14367 ^ n14217;
  assign n15004 = n15003 ^ n14367;
  assign n15005 = n14371 ^ n14367;
  assign n15006 = n15004 & n15005;
  assign n15007 = n15006 ^ n14367;
  assign n15008 = n14373 & n15007;
  assign n15009 = ~n15002 & ~n15008;
  assign n15010 = ~n14365 & n14396;
  assign n15011 = n14218 & ~n15010;
  assign n15012 = n14351 & n14355;
  assign n15013 = n14353 & n14394;
  assign n15014 = n14218 & n14367;
  assign n15015 = n14355 & ~n14389;
  assign n15016 = ~n15014 & ~n15015;
  assign n15017 = ~n15013 & n15016;
  assign n15018 = ~n15012 & n15017;
  assign n15019 = ~n14365 & ~n14387;
  assign n15020 = n14353 & ~n15019;
  assign n15021 = ~n14358 & ~n14383;
  assign n15022 = ~n14371 & n15021;
  assign n15023 = n14218 & ~n15022;
  assign n15024 = ~n15020 & ~n15023;
  assign n15025 = n14355 & ~n14396;
  assign n15026 = ~n14376 & ~n14388;
  assign n15027 = ~n14390 & n15026;
  assign n15028 = ~n14394 & n15027;
  assign n15029 = n14382 & ~n15028;
  assign n15030 = ~n15025 & ~n15029;
  assign n15031 = n15024 & n15030;
  assign n15032 = n14360 & n15031;
  assign n15033 = n15018 & n15032;
  assign n15034 = ~n15011 & n15033;
  assign n15035 = ~n14362 & ~n14376;
  assign n15036 = n15035 ^ n14380;
  assign n15037 = n15036 ^ n14380;
  assign n15038 = n14380 ^ n14217;
  assign n15039 = n15038 ^ n14380;
  assign n15040 = ~n15037 & ~n15039;
  assign n15041 = n15040 ^ n14380;
  assign n15042 = ~n14373 & n15041;
  assign n15043 = n15042 ^ n14380;
  assign n15044 = n15034 & ~n15043;
  assign n15045 = n15009 & n15044;
  assign n15046 = ~n15001 & n15045;
  assign n15047 = ~n14999 & n15046;
  assign n15048 = n15047 ^ n11469;
  assign n15049 = n15048 ^ x602;
  assign n15050 = ~n14997 & n15049;
  assign n15051 = n13751 & n13767;
  assign n15052 = n13777 & ~n15051;
  assign n15053 = n13769 & n13773;
  assign n15054 = n13700 & n13753;
  assign n15055 = n13760 & n15054;
  assign n15056 = ~n15053 & ~n15055;
  assign n15057 = ~n13701 & ~n13806;
  assign n15058 = n13769 & ~n15057;
  assign n15059 = n13760 & n13767;
  assign n15060 = n13751 & n13764;
  assign n15061 = ~n15059 & ~n15060;
  assign n15062 = ~n13794 & ~n13806;
  assign n15063 = ~n13790 & n15062;
  assign n15064 = n13751 & ~n15063;
  assign n15065 = ~n13758 & ~n13807;
  assign n15066 = n13751 & ~n15065;
  assign n15067 = n13753 & n13757;
  assign n15068 = ~n13795 & ~n13802;
  assign n15069 = ~n15067 & n15068;
  assign n15070 = ~n13807 & n15069;
  assign n15071 = n13765 & ~n15070;
  assign n15072 = ~n13755 & ~n13795;
  assign n15073 = ~n13791 & ~n15072;
  assign n15074 = ~n15071 & ~n15073;
  assign n15075 = ~n15066 & n15074;
  assign n15077 = n13757 & n13793;
  assign n15078 = ~n15054 & ~n15077;
  assign n15076 = n13803 & ~n13806;
  assign n15079 = n15078 ^ n15076;
  assign n15080 = n15079 ^ n15078;
  assign n15081 = n15078 ^ n13714;
  assign n15082 = n15081 ^ n15078;
  assign n15083 = ~n15080 & ~n15082;
  assign n15084 = n15083 ^ n15078;
  assign n15085 = ~n13750 & ~n15084;
  assign n15086 = n15085 ^ n15078;
  assign n15087 = n15075 & n15086;
  assign n15088 = ~n15064 & n15087;
  assign n15089 = n15061 & n15088;
  assign n15090 = ~n15058 & n15089;
  assign n15091 = n15056 & n15090;
  assign n15092 = n13772 & n15091;
  assign n15093 = n15052 & n15092;
  assign n15094 = n15093 ^ n11785;
  assign n15095 = n15094 ^ x599;
  assign n15096 = n14519 & n14556;
  assign n15097 = n14545 & n15096;
  assign n15098 = ~n14557 & ~n14571;
  assign n15099 = ~n14569 & n15098;
  assign n15100 = n14579 & ~n15099;
  assign n15101 = n14460 & n14585;
  assign n15102 = ~n14460 & ~n14569;
  assign n15103 = n15098 & n15102;
  assign n15104 = ~n14584 & n15103;
  assign n15105 = n14542 & n14568;
  assign n15106 = ~n14570 & ~n14584;
  assign n15107 = ~n15105 & n15106;
  assign n15108 = ~n14545 & n15107;
  assign n15109 = ~n15104 & ~n15108;
  assign n15110 = n14457 & n15109;
  assign n15111 = n14581 & ~n15096;
  assign n15112 = ~n14558 & n15111;
  assign n15113 = n14579 & ~n15112;
  assign n15114 = ~n14585 & n15107;
  assign n15115 = n14459 & ~n15114;
  assign n15116 = ~n15113 & ~n15115;
  assign n15117 = ~n15110 & n15116;
  assign n15118 = ~n15101 & n15117;
  assign n15119 = ~n15100 & n15118;
  assign n15120 = ~n15097 & n15119;
  assign n15121 = n14566 ^ n14561;
  assign n15122 = n15121 ^ n14561;
  assign n15123 = n14561 ^ n14458;
  assign n15124 = n15123 ^ n14561;
  assign n15125 = ~n15122 & n15124;
  assign n15126 = n15125 ^ n14561;
  assign n15127 = ~n14457 & ~n15126;
  assign n15128 = n15127 ^ n14561;
  assign n15129 = n15120 & n15128;
  assign n15130 = ~n14544 & n15129;
  assign n15131 = n14567 ^ n14460;
  assign n15132 = n14567 ^ n14459;
  assign n15133 = n15132 ^ n14459;
  assign n15134 = n14548 ^ n14459;
  assign n15135 = ~n15133 & ~n15134;
  assign n15136 = n15135 ^ n14459;
  assign n15137 = n15131 & n15136;
  assign n15138 = n15137 ^ n14460;
  assign n15139 = n15130 & ~n15138;
  assign n15140 = n15139 ^ n11634;
  assign n15141 = n15140 ^ x601;
  assign n15142 = n15095 & ~n15141;
  assign n15143 = n15050 & n15142;
  assign n15144 = n14959 & n15143;
  assign n15145 = ~n15095 & n15141;
  assign n15146 = n14997 & ~n15049;
  assign n15147 = n15145 & n15146;
  assign n15148 = n14959 & n15147;
  assign n15149 = n14818 & n14958;
  assign n15150 = n15142 & n15146;
  assign n15151 = n15149 & n15150;
  assign n15152 = ~n14818 & n14958;
  assign n15153 = n15143 & n15152;
  assign n15154 = ~n15151 & ~n15153;
  assign n15155 = ~n15148 & n15154;
  assign n15156 = ~n14997 & ~n15049;
  assign n15157 = ~n15095 & ~n15141;
  assign n15158 = n15156 & n15157;
  assign n15159 = n14997 & n15049;
  assign n15160 = n15157 & n15159;
  assign n15161 = ~n15158 & ~n15160;
  assign n15162 = n14959 & ~n15161;
  assign n15164 = ~n14818 & ~n14958;
  assign n15163 = n15142 & n15159;
  assign n15165 = n15164 ^ n15163;
  assign n15166 = n15163 ^ n15152;
  assign n15167 = n15166 ^ n15152;
  assign n15168 = n15095 & n15141;
  assign n15169 = n15156 & n15168;
  assign n15170 = n15169 ^ n15152;
  assign n15171 = ~n15167 & ~n15170;
  assign n15172 = n15171 ^ n15152;
  assign n15173 = n15165 & n15172;
  assign n15174 = n15173 ^ n15164;
  assign n15175 = ~n15162 & ~n15174;
  assign n15176 = n15145 & n15159;
  assign n15177 = n14958 & n15176;
  assign n15178 = n15050 & n15168;
  assign n15179 = n15146 & n15168;
  assign n15180 = ~n15178 & ~n15179;
  assign n15181 = ~n15163 & ~n15169;
  assign n15182 = n15180 & n15181;
  assign n15183 = n14959 & ~n15182;
  assign n15184 = n15145 & n15156;
  assign n15185 = n15050 & n15157;
  assign n15186 = ~n15147 & ~n15185;
  assign n15187 = ~n15184 & n15186;
  assign n15188 = ~n15160 & n15187;
  assign n15189 = ~n14958 & n15188;
  assign n15190 = n15050 & n15145;
  assign n15191 = n15146 & n15157;
  assign n15192 = ~n15190 & ~n15191;
  assign n15193 = n14958 ^ n14818;
  assign n15194 = ~n15184 & ~n15185;
  assign n15195 = ~n15164 & n15194;
  assign n15196 = ~n15193 & ~n15195;
  assign n15197 = n15192 & ~n15196;
  assign n15198 = ~n15189 & ~n15197;
  assign n15199 = ~n15183 & ~n15198;
  assign n15200 = ~n15177 & n15199;
  assign n15203 = n15159 & n15168;
  assign n15204 = n15142 & n15156;
  assign n15205 = ~n15203 & ~n15204;
  assign n15201 = ~n15158 & ~n15179;
  assign n15202 = ~n15150 & n15201;
  assign n15206 = n15205 ^ n15202;
  assign n15207 = n15206 ^ n15205;
  assign n15208 = n15205 ^ n14958;
  assign n15209 = n15208 ^ n15205;
  assign n15210 = ~n15207 & n15209;
  assign n15211 = n15210 ^ n15205;
  assign n15212 = n15193 & ~n15211;
  assign n15213 = n15212 ^ n15205;
  assign n15214 = n15200 & n15213;
  assign n15215 = n15175 & n15214;
  assign n15216 = n15155 & n15215;
  assign n15217 = ~n15144 & n15216;
  assign n15218 = n15217 ^ n13749;
  assign n15219 = n15218 ^ x682;
  assign n15220 = ~n14783 & ~n15219;
  assign n15221 = n13385 & n13393;
  assign n15222 = n12599 & ~n14961;
  assign n15223 = ~n15221 & ~n15222;
  assign n15224 = n13393 & n13410;
  assign n15225 = ~n13406 & n13434;
  assign n15226 = ~n15224 & ~n15225;
  assign n15227 = n13385 & n13434;
  assign n15228 = ~n13401 & n13420;
  assign n15229 = ~n13389 & n15228;
  assign n15230 = ~n13405 & n15229;
  assign n15231 = n13398 & ~n15230;
  assign n15232 = ~n15227 & ~n15231;
  assign n15233 = n13390 & ~n13401;
  assign n15234 = ~n13404 & n15233;
  assign n15235 = n13393 & ~n15234;
  assign n15236 = n14960 ^ n13395;
  assign n15237 = n15236 ^ n13395;
  assign n15238 = n13425 ^ n13395;
  assign n15239 = n15237 & n15238;
  assign n15240 = n15239 ^ n13395;
  assign n15241 = ~n15235 & ~n15240;
  assign n15242 = n15232 & n15241;
  assign n15243 = n15226 & n15242;
  assign n15244 = ~n14969 & n15243;
  assign n15245 = n14974 & n15244;
  assign n15246 = ~n13392 & n15245;
  assign n15247 = ~n14971 & n15246;
  assign n15248 = n15223 & n15247;
  assign n15249 = n15248 ^ n13036;
  assign n15250 = n15249 ^ x628;
  assign n15251 = n14889 & ~n14918;
  assign n15252 = ~n14890 & n14897;
  assign n15253 = n14893 & ~n15252;
  assign n15254 = ~n14890 & n14923;
  assign n15255 = n14889 & n14943;
  assign n15256 = n14888 & n14896;
  assign n15257 = ~n15255 & ~n15256;
  assign n15258 = ~n15254 & n15257;
  assign n15259 = n14889 & n14896;
  assign n15260 = n14849 ^ n14848;
  assign n15261 = n14877 ^ n14851;
  assign n15262 = n15261 ^ n14849;
  assign n15263 = n15260 & ~n15262;
  assign n15264 = ~n14917 & ~n15263;
  assign n15265 = ~n14947 & n15264;
  assign n15266 = n14821 & ~n15265;
  assign n15267 = ~n15259 & ~n15266;
  assign n15268 = ~n14879 & n14930;
  assign n15269 = n15268 ^ n14881;
  assign n15270 = ~n14913 & ~n14943;
  assign n15271 = n15270 ^ n15268;
  assign n15272 = n15271 ^ n15270;
  assign n15273 = ~n14908 & ~n14927;
  assign n15274 = ~n14916 & n15273;
  assign n15275 = ~n14900 & n15274;
  assign n15276 = n14888 & ~n15275;
  assign n15277 = n15276 ^ n15270;
  assign n15278 = ~n15272 & n15277;
  assign n15279 = n15278 ^ n15270;
  assign n15280 = ~n15269 & n15279;
  assign n15281 = n15280 ^ n14881;
  assign n15282 = n15267 & ~n15281;
  assign n15283 = n14907 & n15282;
  assign n15284 = n15258 & n15283;
  assign n15285 = n15253 & n15284;
  assign n15286 = ~n15251 & n15285;
  assign n15287 = n15286 ^ n13059;
  assign n15288 = n15287 ^ x633;
  assign n15289 = n15250 & n15288;
  assign n15290 = n13230 ^ x562;
  assign n15291 = n14348 ^ x567;
  assign n15292 = n15290 & n15291;
  assign n15293 = n12092 ^ x563;
  assign n15294 = n14183 ^ x566;
  assign n15295 = n13955 & ~n13970;
  assign n15296 = n13999 & n14013;
  assign n15297 = ~n13953 & ~n13959;
  assign n15298 = ~n14017 & ~n15297;
  assign n15299 = ~n13996 & n14526;
  assign n15300 = ~n13977 & n15299;
  assign n15301 = n13894 & ~n15300;
  assign n15302 = ~n15298 & ~n15301;
  assign n15303 = ~n13892 & n13975;
  assign n15304 = n13970 & n14203;
  assign n15305 = n13963 & ~n15304;
  assign n15306 = ~n13966 & ~n14005;
  assign n15307 = n13999 & ~n15306;
  assign n15308 = ~n13983 & n14009;
  assign n15309 = ~n14000 & n15308;
  assign n15310 = n13955 & ~n15309;
  assign n15311 = ~n15307 & ~n15310;
  assign n15312 = ~n15305 & n15311;
  assign n15313 = ~n15303 & n15312;
  assign n15314 = n15302 & n15313;
  assign n15315 = ~n14186 & n15314;
  assign n15316 = ~n15296 & n15315;
  assign n15317 = ~n15295 & n15316;
  assign n15318 = n13956 ^ n13892;
  assign n15319 = n15318 ^ n13956;
  assign n15320 = n14000 ^ n13956;
  assign n15321 = n15320 ^ n13956;
  assign n15322 = ~n15319 & n15321;
  assign n15323 = n15322 ^ n13956;
  assign n15324 = ~n13893 & n15323;
  assign n15325 = n15324 ^ n13956;
  assign n15326 = n15317 & ~n15325;
  assign n15327 = n13995 & n15326;
  assign n15328 = n15327 ^ n12237;
  assign n15329 = n15328 ^ x565;
  assign n15330 = n15294 & n15329;
  assign n15331 = n15293 & n15330;
  assign n15332 = ~n12567 & ~n12581;
  assign n15333 = ~n12532 & n15332;
  assign n15334 = n12175 & ~n15333;
  assign n15335 = n14475 & ~n14491;
  assign n15336 = ~n12562 & n15335;
  assign n15337 = n12530 & ~n15336;
  assign n15338 = ~n15334 & ~n15337;
  assign n15339 = n12570 & n14483;
  assign n15340 = ~n12547 & n15339;
  assign n15341 = n12526 & ~n15340;
  assign n15343 = ~n12564 & n12576;
  assign n15342 = ~n12549 & n12578;
  assign n15344 = n15343 ^ n15342;
  assign n15345 = n15343 ^ n12542;
  assign n15346 = n15343 & n15345;
  assign n15347 = n15346 ^ n15343;
  assign n15348 = n15344 & n15347;
  assign n15349 = n15348 ^ n15346;
  assign n15350 = n15349 ^ n15343;
  assign n15351 = n15350 ^ n12542;
  assign n15352 = ~n15341 & n15351;
  assign n15353 = n15352 ^ n15341;
  assign n15354 = n15338 & ~n15353;
  assign n15355 = ~n14607 & n15354;
  assign n15356 = n12540 & n15355;
  assign n15357 = n15356 ^ n12201;
  assign n15358 = n15357 ^ x564;
  assign n15359 = ~n15294 & n15358;
  assign n15360 = ~n15293 & n15359;
  assign n15361 = n15329 & n15360;
  assign n15362 = ~n15331 & ~n15361;
  assign n15363 = ~n15293 & ~n15358;
  assign n15364 = n15363 ^ n15329;
  assign n15365 = n15293 & ~n15294;
  assign n15366 = n15365 ^ n15363;
  assign n15367 = n15366 ^ n15365;
  assign n15368 = n15365 ^ n15294;
  assign n15369 = n15367 & ~n15368;
  assign n15370 = n15369 ^ n15365;
  assign n15371 = ~n15364 & ~n15370;
  assign n15372 = n15371 ^ n15329;
  assign n15373 = n15362 & n15372;
  assign n15374 = n15292 & ~n15373;
  assign n15375 = ~n15290 & ~n15291;
  assign n15376 = n15358 ^ n15294;
  assign n15377 = ~n15329 & ~n15376;
  assign n15378 = ~n15293 & n15377;
  assign n15379 = n15358 ^ n15293;
  assign n15380 = n15294 & ~n15329;
  assign n15381 = ~n15379 & n15380;
  assign n15382 = ~n15294 & ~n15358;
  assign n15383 = n15293 & n15382;
  assign n15384 = n15293 & ~n15358;
  assign n15385 = ~n15360 & ~n15384;
  assign n15386 = n15329 & ~n15385;
  assign n15387 = ~n15383 & ~n15386;
  assign n15388 = ~n15381 & n15387;
  assign n15389 = ~n15378 & n15388;
  assign n15390 = n15375 & ~n15389;
  assign n15391 = ~n15374 & ~n15390;
  assign n15392 = n15291 ^ n15290;
  assign n15393 = ~n15329 & n15376;
  assign n15394 = n15293 & n15393;
  assign n15395 = n15330 ^ n15293;
  assign n15396 = n15395 ^ n15330;
  assign n15397 = n15330 ^ n15329;
  assign n15398 = n15397 ^ n15330;
  assign n15399 = ~n15396 & n15398;
  assign n15400 = n15399 ^ n15330;
  assign n15401 = ~n15358 & n15400;
  assign n15402 = n15401 ^ n15330;
  assign n15403 = ~n15394 & ~n15402;
  assign n15404 = ~n15378 & n15403;
  assign n15405 = n15404 ^ n15291;
  assign n15406 = n15405 ^ n15404;
  assign n15407 = n15294 & ~n15379;
  assign n15408 = ~n15294 & ~n15329;
  assign n15409 = n15408 ^ n15293;
  assign n15410 = n15409 ^ n15408;
  assign n15411 = n15329 & ~n15382;
  assign n15412 = n15411 ^ n15408;
  assign n15413 = n15410 & n15412;
  assign n15414 = n15413 ^ n15408;
  assign n15415 = ~n15407 & ~n15414;
  assign n15416 = n15415 ^ n15404;
  assign n15417 = n15406 & ~n15416;
  assign n15418 = n15417 ^ n15404;
  assign n15419 = n15392 & ~n15418;
  assign n15420 = n15391 & ~n15419;
  assign n15421 = n15420 ^ n13072;
  assign n15422 = n15421 ^ x630;
  assign n15423 = n14355 & n14394;
  assign n15424 = n14382 & ~n15035;
  assign n15425 = ~n15423 & ~n15424;
  assign n15426 = n14373 & n14400;
  assign n15427 = n14377 & n14407;
  assign n15428 = n14353 & ~n15427;
  assign n15429 = ~n15426 & ~n15428;
  assign n15430 = ~n14184 & ~n15010;
  assign n15431 = ~n14374 & n15021;
  assign n15432 = n14355 & ~n15431;
  assign n15433 = n14402 & n15035;
  assign n15434 = ~n14383 & n15433;
  assign n15435 = n14218 & ~n15434;
  assign n15436 = ~n15432 & ~n15435;
  assign n15437 = ~n15430 & n15436;
  assign n15438 = n15429 & n15437;
  assign n15439 = n15425 & n15438;
  assign n15440 = ~n14999 & n15439;
  assign n15441 = n15018 & n15440;
  assign n15442 = ~n14352 & n15441;
  assign n15443 = n15442 ^ n13130;
  assign n15444 = n15443 ^ x629;
  assign n15445 = n15422 & ~n15444;
  assign n15446 = n14099 & n14108;
  assign n15447 = ~n14092 & ~n14123;
  assign n15448 = n14089 & ~n15447;
  assign n15449 = ~n15446 & ~n15448;
  assign n15450 = n14080 & n14116;
  assign n15451 = ~n14047 & n14114;
  assign n15452 = n14097 & ~n15451;
  assign n15453 = ~n14048 & n14089;
  assign n15454 = n14094 & n14108;
  assign n15455 = n14081 & n14103;
  assign n15456 = ~n15454 & ~n15455;
  assign n15457 = ~n15453 & n15456;
  assign n15458 = n14043 & n14083;
  assign n15459 = ~n14110 & ~n15458;
  assign n15460 = ~n14122 & ~n15459;
  assign n15461 = ~n14087 & ~n14094;
  assign n15462 = ~n14123 & n15461;
  assign n15463 = n14081 & ~n15462;
  assign n15464 = ~n15460 & ~n15463;
  assign n15465 = ~n14107 & ~n14124;
  assign n15466 = n14103 & n14108;
  assign n15467 = n15465 & ~n15466;
  assign n15468 = n15467 ^ n14049;
  assign n15469 = n15468 ^ n15467;
  assign n15470 = n13891 & n14046;
  assign n15471 = ~n14113 & ~n15470;
  assign n15472 = n15471 ^ n15467;
  assign n15473 = n15472 ^ n15467;
  assign n15474 = n15469 & ~n15473;
  assign n15475 = n15474 ^ n15467;
  assign n15476 = ~n14080 & ~n15475;
  assign n15477 = n15476 ^ n15467;
  assign n15478 = n15464 & n15477;
  assign n15479 = ~n14101 & n15478;
  assign n15480 = n15457 & n15479;
  assign n15481 = ~n15452 & n15480;
  assign n15482 = ~n15450 & n15481;
  assign n15483 = n15449 & n15482;
  assign n15484 = n14091 & n15483;
  assign n15485 = n15484 ^ n13168;
  assign n15486 = n15485 ^ x632;
  assign n15487 = n13760 & ~n15069;
  assign n15488 = ~n13773 & ~n15054;
  assign n15489 = n13751 & ~n15488;
  assign n15490 = ~n15487 & ~n15489;
  assign n15491 = n13765 & ~n15068;
  assign n15492 = n13760 & ~n13808;
  assign n15493 = ~n13755 & n15488;
  assign n15494 = n15493 ^ n13796;
  assign n15495 = n15493 ^ n13714;
  assign n15496 = n15495 ^ n15493;
  assign n15497 = n15494 & n15496;
  assign n15498 = n15497 ^ n15493;
  assign n15499 = n13750 & ~n15498;
  assign n15500 = ~n15492 & ~n15499;
  assign n15501 = ~n15491 & n15500;
  assign n15502 = n15077 ^ n13803;
  assign n15503 = n15502 ^ n13803;
  assign n15504 = n13803 ^ n13714;
  assign n15505 = n15504 ^ n13803;
  assign n15506 = n15503 & n15505;
  assign n15507 = n15506 ^ n13803;
  assign n15508 = ~n13750 & ~n15507;
  assign n15509 = n15508 ^ n13803;
  assign n15510 = n15501 & n15509;
  assign n15511 = ~n15064 & n15510;
  assign n15512 = n15061 & n15511;
  assign n15513 = ~n15058 & n15512;
  assign n15514 = n13762 & n15513;
  assign n15515 = n15490 & n15514;
  assign n15516 = n13771 & n15515;
  assign n15517 = n15516 ^ n13099;
  assign n15518 = n15517 ^ x631;
  assign n15519 = ~n15486 & ~n15518;
  assign n15520 = n15445 & n15519;
  assign n15521 = n15289 & n15520;
  assign n15522 = n15422 & n15444;
  assign n15523 = ~n15486 & n15518;
  assign n15524 = n15522 & n15523;
  assign n15525 = n15486 & ~n15518;
  assign n15526 = n15522 & n15525;
  assign n15527 = ~n15524 & ~n15526;
  assign n15528 = n15289 & ~n15527;
  assign n15529 = ~n15250 & n15288;
  assign n15530 = ~n15422 & n15444;
  assign n15531 = n15525 & n15530;
  assign n15532 = n15519 & n15522;
  assign n15533 = ~n15531 & ~n15532;
  assign n15534 = n15529 & ~n15533;
  assign n15535 = ~n15528 & ~n15534;
  assign n15536 = ~n15521 & n15535;
  assign n15537 = n15486 & n15518;
  assign n15538 = ~n15422 & ~n15444;
  assign n15539 = n15537 & n15538;
  assign n15540 = n15529 & n15539;
  assign n15541 = n15519 & n15538;
  assign n15542 = n15289 & n15541;
  assign n15543 = ~n15540 & ~n15542;
  assign n15544 = n15445 & n15537;
  assign n15545 = n15445 & n15525;
  assign n15546 = ~n15544 & ~n15545;
  assign n15547 = n15289 & ~n15546;
  assign n15548 = n15525 & n15538;
  assign n15549 = ~n15520 & ~n15548;
  assign n15550 = n15529 & ~n15549;
  assign n15551 = ~n15547 & ~n15550;
  assign n15552 = ~n15250 & ~n15288;
  assign n15553 = n15486 ^ n15422;
  assign n15554 = n15553 ^ n15444;
  assign n15555 = n15554 ^ n15486;
  assign n15556 = n15555 ^ n15444;
  assign n15557 = n15556 ^ n15518;
  assign n15558 = n15486 ^ n15444;
  assign n15559 = n15518 ^ n15486;
  assign n15560 = n15559 ^ n15486;
  assign n15561 = n15558 & ~n15560;
  assign n15562 = n15561 ^ n15486;
  assign n15563 = ~n15557 & n15562;
  assign n15564 = n15563 ^ n15554;
  assign n15565 = n15552 & ~n15564;
  assign n15566 = n15250 & ~n15288;
  assign n15567 = n15445 & n15523;
  assign n15568 = ~n15548 & ~n15567;
  assign n15569 = ~n15541 & ~n15545;
  assign n15570 = ~n15532 & n15569;
  assign n15571 = n15568 & n15570;
  assign n15572 = ~n15526 & n15571;
  assign n15573 = n15566 & ~n15572;
  assign n15575 = n15523 & n15530;
  assign n15574 = ~n15529 & ~n15566;
  assign n15576 = n15575 ^ n15574;
  assign n15577 = n15522 & n15537;
  assign n15578 = n15577 ^ n15574;
  assign n15579 = n15578 ^ n15577;
  assign n15580 = n15577 ^ n15289;
  assign n15581 = n15579 & ~n15580;
  assign n15582 = n15581 ^ n15577;
  assign n15583 = ~n15576 & n15582;
  assign n15584 = n15583 ^ n15575;
  assign n15585 = ~n15573 & ~n15584;
  assign n15586 = ~n15565 & n15585;
  assign n15587 = n15551 & n15586;
  assign n15588 = n15567 ^ n15250;
  assign n15589 = n15588 ^ n15567;
  assign n15590 = n15567 ^ n15531;
  assign n15591 = n15589 & n15590;
  assign n15592 = n15591 ^ n15567;
  assign n15593 = n15288 & n15592;
  assign n15594 = n15587 & ~n15593;
  assign n15595 = n15543 & n15594;
  assign n15596 = n15536 & n15595;
  assign n15597 = n15596 ^ n13655;
  assign n15598 = n15597 ^ x686;
  assign n15599 = n14146 ^ x609;
  assign n15600 = n15048 ^ x604;
  assign n15601 = ~n15599 & n15600;
  assign n15602 = n15379 ^ n15293;
  assign n15603 = n15294 ^ n15293;
  assign n15604 = n15603 ^ n15358;
  assign n15605 = n15604 ^ n15293;
  assign n15606 = n15605 ^ n15293;
  assign n15607 = n15602 & n15606;
  assign n15608 = n15607 ^ n15293;
  assign n15609 = ~n15329 & n15608;
  assign n15610 = n15609 ^ n15604;
  assign n15611 = n15375 & ~n15610;
  assign n15612 = n15290 & ~n15291;
  assign n15613 = n15376 ^ n15329;
  assign n15614 = n15613 ^ n15293;
  assign n15615 = n15614 ^ n15358;
  assign n15616 = n15615 ^ n15329;
  assign n15617 = n15358 ^ n15329;
  assign n15618 = n15379 ^ n15358;
  assign n15619 = ~n15617 & n15618;
  assign n15620 = n15619 ^ n15358;
  assign n15621 = ~n15616 & n15620;
  assign n15622 = n15621 ^ n15613;
  assign n15623 = n15612 & n15622;
  assign n15624 = ~n15611 & ~n15623;
  assign n15625 = n15380 & n15384;
  assign n15626 = ~n15294 & n15379;
  assign n15627 = ~n15293 & n15330;
  assign n15628 = ~n15329 & n15359;
  assign n15629 = ~n15627 & ~n15628;
  assign n15630 = ~n15626 & n15629;
  assign n15631 = ~n15625 & n15630;
  assign n15632 = n15292 & ~n15631;
  assign n15633 = ~n15290 & n15291;
  assign n15634 = n15293 & n15380;
  assign n15635 = ~n15363 & ~n15365;
  assign n15636 = n15329 & ~n15635;
  assign n15637 = ~n15634 & ~n15636;
  assign n15638 = ~n15378 & n15637;
  assign n15639 = n15633 & ~n15638;
  assign n15640 = ~n15632 & ~n15639;
  assign n15641 = n15624 & n15640;
  assign n15642 = n15641 ^ n13476;
  assign n15643 = n15642 ^ x606;
  assign n15644 = n14601 ^ x608;
  assign n15645 = ~n15643 & ~n15644;
  assign n15646 = n14817 ^ x605;
  assign n15647 = n14889 & n14910;
  assign n15648 = n14821 & ~n15273;
  assign n15649 = ~n15647 & ~n15648;
  assign n15650 = ~n14900 & ~n14923;
  assign n15651 = n14881 & ~n15650;
  assign n15652 = n14884 & n14889;
  assign n15653 = ~n14890 & n14947;
  assign n15654 = ~n15652 & ~n15653;
  assign n15655 = ~n14900 & ~n14928;
  assign n15656 = ~n14897 & n15655;
  assign n15657 = ~n14913 & n15656;
  assign n15658 = n14821 & ~n15657;
  assign n15659 = ~n14917 & n14930;
  assign n15660 = ~n14884 & n15655;
  assign n15661 = ~n14879 & n15660;
  assign n15662 = n14888 & ~n15661;
  assign n15663 = ~n14881 & ~n15662;
  assign n15664 = ~n15659 & ~n15663;
  assign n15665 = ~n15658 & ~n15664;
  assign n15666 = n15654 & n15665;
  assign n15667 = n14887 ^ n14881;
  assign n15668 = n14898 ^ n14820;
  assign n15669 = n14887 ^ n14820;
  assign n15670 = n15669 ^ n14820;
  assign n15671 = n15668 & ~n15670;
  assign n15672 = n15671 ^ n14820;
  assign n15673 = n15667 & n15672;
  assign n15674 = n15673 ^ n14881;
  assign n15675 = n15666 & ~n15674;
  assign n15676 = n14912 & n15675;
  assign n15677 = ~n15651 & n15676;
  assign n15678 = n15258 & n15677;
  assign n15679 = n15649 & n15678;
  assign n15680 = ~n15251 & n15679;
  assign n15681 = n15680 ^ n13518;
  assign n15682 = n15681 ^ x607;
  assign n15683 = ~n15646 & n15682;
  assign n15684 = n15645 & n15683;
  assign n15685 = n15601 & n15684;
  assign n15686 = n15599 & n15600;
  assign n15687 = n15646 & ~n15682;
  assign n15688 = n15645 & n15687;
  assign n15689 = n15686 & n15688;
  assign n15690 = n15643 & n15644;
  assign n15691 = n15687 & n15690;
  assign n15692 = n15686 & n15691;
  assign n15693 = ~n15689 & ~n15692;
  assign n15694 = ~n15599 & ~n15600;
  assign n15695 = n15646 & n15682;
  assign n15696 = n15645 & n15695;
  assign n15697 = ~n15643 & n15644;
  assign n15698 = n15687 & n15697;
  assign n15699 = ~n15696 & ~n15698;
  assign n15700 = ~n15691 & n15699;
  assign n15701 = n15694 & ~n15700;
  assign n15702 = n15600 ^ n15599;
  assign n15703 = n15690 & n15695;
  assign n15704 = ~n15702 & n15703;
  assign n15705 = n15643 & ~n15644;
  assign n15706 = n15683 & n15705;
  assign n15707 = n15686 & n15706;
  assign n15708 = ~n15704 & ~n15707;
  assign n15709 = n15599 & ~n15600;
  assign n15710 = n15644 ^ n15643;
  assign n15711 = n15710 ^ n15682;
  assign n15712 = n15646 & n15711;
  assign n15713 = n15709 & n15712;
  assign n15714 = n15695 & n15697;
  assign n15715 = n15687 & n15705;
  assign n15716 = ~n15714 & ~n15715;
  assign n15717 = ~n15698 & n15716;
  assign n15718 = n15683 & n15697;
  assign n15719 = ~n15646 & ~n15682;
  assign n15720 = n15645 & n15719;
  assign n15721 = ~n15718 & ~n15720;
  assign n15722 = n15683 & n15690;
  assign n15723 = n15705 & n15719;
  assign n15724 = ~n15722 & ~n15723;
  assign n15725 = n15721 & n15724;
  assign n15726 = n15717 & n15725;
  assign n15727 = n15601 & ~n15726;
  assign n15728 = ~n15713 & ~n15727;
  assign n15729 = n15690 & n15719;
  assign n15730 = ~n15684 & ~n15729;
  assign n15731 = n15721 & n15730;
  assign n15732 = n15731 ^ n15600;
  assign n15733 = n15732 ^ n15731;
  assign n15734 = n15697 & n15719;
  assign n15735 = ~n15684 & ~n15722;
  assign n15736 = ~n15688 & n15735;
  assign n15737 = ~n15734 & n15736;
  assign n15738 = n15737 ^ n15731;
  assign n15739 = n15738 ^ n15731;
  assign n15740 = ~n15733 & ~n15739;
  assign n15741 = n15740 ^ n15731;
  assign n15742 = ~n15599 & ~n15741;
  assign n15743 = n15742 ^ n15731;
  assign n15744 = n15728 & n15743;
  assign n15745 = n15708 & n15744;
  assign n15746 = ~n15701 & n15745;
  assign n15747 = n15693 & n15746;
  assign n15748 = ~n15685 & n15747;
  assign n15749 = n15748 ^ n13592;
  assign n15750 = n15749 ^ x684;
  assign n15751 = ~n15598 & n15750;
  assign n15752 = n15375 & ~n15415;
  assign n15753 = n15373 & n15612;
  assign n15754 = ~n15752 & ~n15753;
  assign n15755 = n15292 & ~n15404;
  assign n15756 = ~n15389 & n15633;
  assign n15757 = ~n15755 & ~n15756;
  assign n15758 = n15754 & n15757;
  assign n15759 = n15758 ^ n12294;
  assign n15760 = n15759 ^ x622;
  assign n15761 = n15443 ^ x627;
  assign n15762 = ~n15760 & ~n15761;
  assign n15763 = n15249 ^ x626;
  assign n15764 = ~n14693 & ~n14705;
  assign n15765 = n14605 & ~n15764;
  assign n15766 = n14678 & n14697;
  assign n15767 = ~n14666 & ~n14670;
  assign n15768 = n14668 & ~n15767;
  assign n15769 = ~n15766 & ~n15768;
  assign n15770 = n14605 & n14697;
  assign n15771 = n14668 & ~n14700;
  assign n15772 = ~n15770 & ~n15771;
  assign n15773 = n14664 ^ n14627;
  assign n15774 = n15773 ^ n14627;
  assign n15775 = n14661 ^ n14627;
  assign n15776 = n15775 ^ n14627;
  assign n15777 = n15774 & ~n15776;
  assign n15778 = n15777 ^ n14627;
  assign n15779 = n14663 & ~n15778;
  assign n15780 = n14672 & n15779;
  assign n15781 = ~n14680 & ~n14719;
  assign n15782 = n14672 & ~n15781;
  assign n15783 = ~n14687 & ~n15782;
  assign n15784 = n14789 & n15783;
  assign n15785 = n15784 ^ n14604;
  assign n15786 = n15785 ^ n15784;
  assign n15787 = ~n14695 & ~n14718;
  assign n15788 = ~n14704 & n15787;
  assign n15789 = ~n14685 & n15788;
  assign n15790 = ~n14674 & n15789;
  assign n15791 = ~n14670 & n15790;
  assign n15792 = n15791 ^ n15784;
  assign n15793 = n15792 ^ n15784;
  assign n15794 = ~n15786 & ~n15793;
  assign n15795 = n15794 ^ n15784;
  assign n15796 = ~n14603 & ~n15795;
  assign n15797 = n15796 ^ n15784;
  assign n15798 = ~n15780 & n15797;
  assign n15799 = n15772 & n15798;
  assign n15800 = n15769 & n15799;
  assign n15801 = ~n15765 & n15800;
  assign n15802 = ~n14813 & n15801;
  assign n15803 = ~n14667 & n15802;
  assign n15804 = n15803 ^ n13309;
  assign n15805 = n15804 ^ x625;
  assign n15806 = n15763 & ~n15805;
  assign n15807 = ~n13758 & ~n13775;
  assign n15808 = n13765 & ~n15807;
  assign n15809 = ~n13790 & ~n15067;
  assign n15810 = n13750 & ~n15809;
  assign n15811 = ~n15808 & ~n15810;
  assign n15812 = n15062 & n15068;
  assign n15813 = n13751 & ~n15812;
  assign n15814 = ~n13794 & ~n13802;
  assign n15815 = ~n13807 & n15814;
  assign n15816 = ~n13769 & n15815;
  assign n15817 = n15065 & ~n15077;
  assign n15818 = ~n13765 & n15817;
  assign n15819 = ~n15816 & ~n15818;
  assign n15820 = n13750 & n15819;
  assign n15821 = ~n15813 & ~n15820;
  assign n15822 = n15811 & n15821;
  assign n15823 = n13760 ^ n13701;
  assign n15824 = n13769 ^ n13760;
  assign n15825 = n15824 ^ n13769;
  assign n15826 = ~n13755 & ~n15077;
  assign n15827 = n15826 ^ n13769;
  assign n15828 = n15825 & n15827;
  assign n15829 = n15828 ^ n13769;
  assign n15830 = n15823 & ~n15829;
  assign n15831 = n15830 ^ n13701;
  assign n15832 = n15822 & ~n15831;
  assign n15833 = n15056 & n15832;
  assign n15834 = n15052 & n15833;
  assign n15835 = n15490 & n15834;
  assign n15836 = n13771 & n15835;
  assign n15837 = n15836 ^ n12173;
  assign n15838 = n15837 ^ x623;
  assign n15839 = n14460 & ~n14581;
  assign n15840 = ~n14558 & ~n14560;
  assign n15841 = n14459 & ~n15840;
  assign n15842 = ~n15839 & ~n15841;
  assign n15843 = n14459 & n14547;
  assign n15844 = ~n14550 & ~n15096;
  assign n15845 = ~n14548 & n15844;
  assign n15846 = ~n14558 & n15845;
  assign n15847 = n14545 & ~n15846;
  assign n15848 = ~n14459 & n15845;
  assign n15849 = ~n14579 & n15106;
  assign n15850 = ~n14457 & ~n15849;
  assign n15851 = ~n14557 & ~n15850;
  assign n15852 = ~n15848 & ~n15851;
  assign n15853 = n14543 ^ n14457;
  assign n15854 = n15853 ^ n14543;
  assign n15855 = n15102 & ~n15105;
  assign n15856 = ~n14545 & ~n14584;
  assign n15857 = ~n15855 & ~n15856;
  assign n15858 = ~n14567 & ~n15857;
  assign n15859 = ~n14557 & n15858;
  assign n15860 = n15859 ^ n14543;
  assign n15861 = n15854 & ~n15860;
  assign n15862 = n15861 ^ n14543;
  assign n15863 = ~n15852 & ~n15862;
  assign n15864 = ~n15847 & n15863;
  assign n15865 = ~n15843 & n15864;
  assign n15866 = ~n14543 & ~n14560;
  assign n15867 = n15866 ^ n14457;
  assign n15868 = n15867 ^ n15866;
  assign n15869 = n14573 & ~n14584;
  assign n15870 = n15869 ^ n15866;
  assign n15871 = ~n15868 & n15870;
  assign n15872 = n15871 ^ n15866;
  assign n15873 = ~n14458 & ~n15872;
  assign n15874 = n15865 & ~n15873;
  assign n15875 = n15842 & n15874;
  assign n15876 = ~n15101 & n15875;
  assign n15877 = n15876 ^ n13276;
  assign n15878 = n15877 ^ x624;
  assign n15879 = ~n15838 & n15878;
  assign n15880 = n15806 & n15879;
  assign n15881 = n15762 & n15880;
  assign n15882 = n15760 & ~n15761;
  assign n15883 = n15763 & n15805;
  assign n15884 = n15879 & n15883;
  assign n15885 = ~n15763 & ~n15805;
  assign n15886 = n15879 & n15885;
  assign n15887 = ~n15884 & ~n15886;
  assign n15888 = n15882 & ~n15887;
  assign n15889 = ~n15881 & ~n15888;
  assign n15890 = ~n15760 & n15761;
  assign n15891 = n15838 & ~n15878;
  assign n15892 = n15806 & n15891;
  assign n15893 = n15890 & n15892;
  assign n15894 = ~n15838 & ~n15878;
  assign n15895 = n15885 & n15894;
  assign n15896 = n15882 & n15895;
  assign n15897 = ~n15893 & ~n15896;
  assign n15898 = n15760 & n15761;
  assign n15899 = ~n15762 & ~n15898;
  assign n15900 = n15806 & n15894;
  assign n15901 = ~n15886 & ~n15900;
  assign n15902 = ~n15899 & ~n15901;
  assign n15903 = n15897 & ~n15902;
  assign n15904 = ~n15763 & n15805;
  assign n15905 = n15879 & n15904;
  assign n15906 = n15838 & n15878;
  assign n15907 = n15806 & n15906;
  assign n15908 = n15904 & n15906;
  assign n15909 = ~n15907 & ~n15908;
  assign n15910 = ~n15905 & n15909;
  assign n15911 = n15890 & ~n15910;
  assign n15912 = n15898 & n15907;
  assign n15913 = n15885 & n15906;
  assign n15914 = ~n15892 & ~n15913;
  assign n15915 = n15882 & ~n15914;
  assign n15916 = ~n15912 & ~n15915;
  assign n15917 = n15894 & n15904;
  assign n15918 = ~n15899 & n15917;
  assign n15919 = n15884 & n15898;
  assign n15920 = n15883 & n15894;
  assign n15921 = ~n15895 & ~n15920;
  assign n15922 = n15890 & ~n15921;
  assign n15923 = ~n15919 & ~n15922;
  assign n15924 = ~n15918 & n15923;
  assign n15925 = n15760 & n15908;
  assign n15926 = n15891 & n15904;
  assign n15927 = n15898 & n15926;
  assign n15928 = ~n15925 & ~n15927;
  assign n15929 = n15885 & n15891;
  assign n15930 = ~n15899 & n15929;
  assign n15931 = n15883 & n15906;
  assign n15932 = ~n15913 & ~n15931;
  assign n15933 = n15890 & ~n15932;
  assign n15934 = ~n15930 & ~n15933;
  assign n15935 = n15883 & n15891;
  assign n15936 = ~n15880 & ~n15935;
  assign n15937 = n15882 & ~n15936;
  assign n15938 = ~n15926 & ~n15931;
  assign n15939 = ~n15884 & n15938;
  assign n15940 = n15762 & ~n15939;
  assign n15941 = ~n15937 & ~n15940;
  assign n15942 = n15934 & n15941;
  assign n15943 = n15928 & n15942;
  assign n15944 = n15924 & n15943;
  assign n15945 = n15916 & n15944;
  assign n15946 = ~n15911 & n15945;
  assign n15947 = n15903 & n15946;
  assign n15948 = n15889 & n15947;
  assign n15949 = n15948 ^ n13635;
  assign n15950 = n15949 ^ x683;
  assign n15951 = n15094 ^ x597;
  assign n15952 = n14457 & n15105;
  assign n15953 = ~n14585 & n15098;
  assign n15954 = ~n14560 & n15953;
  assign n15955 = n14545 & ~n15954;
  assign n15956 = ~n15952 & ~n15955;
  assign n15957 = n14576 & n14579;
  assign n15958 = ~n14558 & ~n14569;
  assign n15959 = n14460 & ~n15958;
  assign n15960 = n14573 & n14581;
  assign n15961 = n14459 & ~n15960;
  assign n15962 = ~n15959 & ~n15961;
  assign n15963 = ~n15957 & n15962;
  assign n15964 = n15956 & n15963;
  assign n15965 = ~n14554 & n15964;
  assign n15966 = ~n15138 & n15965;
  assign n15967 = n15842 & n15966;
  assign n15968 = ~n15101 & n15967;
  assign n15969 = n15968 ^ n12925;
  assign n15970 = n15969 ^ x592;
  assign n15971 = ~n15951 & ~n15970;
  assign n15972 = n14116 & ~n14122;
  assign n15973 = ~n14047 & ~n15470;
  assign n15974 = ~n14085 & n15973;
  assign n15975 = ~n14110 & n15974;
  assign n15976 = n14108 & ~n15975;
  assign n15977 = ~n14092 & ~n15458;
  assign n15978 = ~n14116 & n15977;
  assign n15979 = ~n14044 & n15978;
  assign n15980 = n14097 & ~n15979;
  assign n15981 = ~n14099 & ~n14130;
  assign n15982 = n14081 & ~n15981;
  assign n15983 = ~n15980 & ~n15982;
  assign n15984 = ~n15976 & n15983;
  assign n15985 = ~n15972 & n15984;
  assign n15986 = n14123 ^ n14089;
  assign n15987 = ~n14094 & ~n15458;
  assign n15988 = n15987 ^ n14080;
  assign n15989 = n14089 ^ n14080;
  assign n15990 = n15989 ^ n14080;
  assign n15991 = n15988 & n15990;
  assign n15992 = n15991 ^ n14080;
  assign n15993 = n15986 & ~n15992;
  assign n15994 = n15993 ^ n14123;
  assign n15995 = n15985 & ~n15994;
  assign n15996 = n14112 & n15995;
  assign n15997 = n14106 & n15996;
  assign n15998 = n14096 & n15997;
  assign n15999 = n15457 & n15998;
  assign n16000 = n15999 ^ n12844;
  assign n16001 = n16000 ^ x594;
  assign n16002 = n14957 ^ x596;
  assign n16003 = ~n16001 & n16002;
  assign n16004 = n15612 & ~n15630;
  assign n16005 = n15610 & n15633;
  assign n16006 = ~n16004 & ~n16005;
  assign n16007 = n15622 ^ n15291;
  assign n16008 = n16007 ^ n15622;
  assign n16009 = n15638 ^ n15622;
  assign n16010 = ~n16008 & n16009;
  assign n16011 = n16010 ^ n15622;
  assign n16012 = ~n15392 & ~n16011;
  assign n16013 = n16006 & ~n16012;
  assign n16014 = ~n15625 & n16013;
  assign n16015 = n16014 ^ n12903;
  assign n16016 = n16015 ^ x593;
  assign n16017 = n14373 & n14383;
  assign n16018 = ~n14390 & ~n14400;
  assign n16019 = ~n14374 & n16018;
  assign n16020 = n14353 & ~n16019;
  assign n16021 = n14355 & ~n14391;
  assign n16022 = ~n14387 & n14397;
  assign n16023 = n14382 & ~n16022;
  assign n16024 = ~n14358 & n15026;
  assign n16025 = ~n14380 & n16024;
  assign n16026 = n14218 & ~n16025;
  assign n16027 = ~n16023 & ~n16026;
  assign n16028 = ~n16021 & n16027;
  assign n16029 = ~n16020 & n16028;
  assign n16030 = ~n16017 & n16029;
  assign n16031 = ~n14354 & n16030;
  assign n16032 = n14370 & n16031;
  assign n16033 = n15009 & n16032;
  assign n16034 = ~n15001 & n16033;
  assign n16035 = n15425 & n16034;
  assign n16036 = n15017 & n16035;
  assign n16037 = ~n14352 & n16036;
  assign n16038 = n16037 ^ n12876;
  assign n16039 = n16038 ^ x595;
  assign n16040 = ~n16016 & n16039;
  assign n16041 = n16003 & n16040;
  assign n16042 = n15971 & n16041;
  assign n16043 = ~n15951 & n15970;
  assign n16044 = ~n16016 & ~n16039;
  assign n16045 = n16003 & n16044;
  assign n16046 = n16043 & n16045;
  assign n16047 = ~n16042 & ~n16046;
  assign n16048 = n15951 & ~n15970;
  assign n16049 = n16001 & n16002;
  assign n16050 = n16016 & ~n16039;
  assign n16051 = n16049 & n16050;
  assign n16052 = n16048 & n16051;
  assign n16053 = n15951 & n15970;
  assign n16054 = ~n16002 & n16050;
  assign n16055 = ~n16001 & n16054;
  assign n16056 = n16053 & n16055;
  assign n16057 = ~n16052 & ~n16056;
  assign n16058 = n16047 & n16057;
  assign n16059 = n16016 & n16039;
  assign n16060 = ~n16002 & n16059;
  assign n16061 = ~n16001 & n16060;
  assign n16062 = n16053 & n16061;
  assign n16063 = n15971 & n16055;
  assign n16064 = ~n16062 & ~n16063;
  assign n16065 = n16043 & n16060;
  assign n16066 = n15971 & n16051;
  assign n16067 = ~n16065 & ~n16066;
  assign n16068 = ~n16002 & n16040;
  assign n16069 = ~n16001 & n16068;
  assign n16070 = n15971 & n16069;
  assign n16071 = n16001 & n16060;
  assign n16072 = n16003 & n16059;
  assign n16073 = n16001 & n16054;
  assign n16074 = ~n16072 & ~n16073;
  assign n16075 = ~n16071 & n16074;
  assign n16076 = n16048 & ~n16075;
  assign n16077 = ~n16070 & ~n16076;
  assign n16078 = ~n15971 & ~n16053;
  assign n16079 = n16001 & n16068;
  assign n16080 = n16044 & n16049;
  assign n16081 = ~n16079 & ~n16080;
  assign n16082 = ~n16078 & ~n16081;
  assign n16083 = ~n16002 & n16044;
  assign n16084 = n16001 & n16083;
  assign n16085 = n16040 & n16049;
  assign n16086 = ~n16055 & ~n16085;
  assign n16087 = n16074 & n16086;
  assign n16088 = ~n16084 & n16087;
  assign n16089 = n16043 & ~n16088;
  assign n16090 = ~n16082 & ~n16089;
  assign n16091 = ~n16001 & n16083;
  assign n16092 = ~n16085 & ~n16091;
  assign n16093 = n16053 & ~n16092;
  assign n16094 = ~n16045 & ~n16069;
  assign n16095 = ~n16079 & ~n16085;
  assign n16096 = n16094 & n16095;
  assign n16097 = n16048 & ~n16096;
  assign n16098 = n16049 & n16059;
  assign n16099 = n16003 & n16050;
  assign n16100 = ~n16098 & ~n16099;
  assign n16101 = ~n15971 & n16100;
  assign n16102 = ~n16073 & ~n16098;
  assign n16103 = ~n16053 & n16102;
  assign n16104 = ~n16101 & ~n16103;
  assign n16105 = ~n16078 & n16104;
  assign n16106 = ~n16097 & ~n16105;
  assign n16107 = ~n16093 & n16106;
  assign n16108 = n16090 & n16107;
  assign n16109 = n16077 & n16108;
  assign n16110 = n16067 & n16109;
  assign n16111 = n16064 & n16110;
  assign n16112 = n16058 & n16111;
  assign n16113 = n16112 ^ n13698;
  assign n16114 = n16113 ^ x685;
  assign n16115 = ~n15950 & ~n16114;
  assign n16116 = n15751 & n16115;
  assign n16117 = n15598 & ~n15750;
  assign n16118 = n16115 & n16117;
  assign n16119 = ~n16116 & ~n16118;
  assign n16120 = n15220 & ~n16119;
  assign n16121 = ~n14783 & n15219;
  assign n16122 = n16118 & n16121;
  assign n16123 = ~n15598 & ~n15750;
  assign n16124 = n16115 & n16123;
  assign n16125 = n15219 & n16124;
  assign n16126 = ~n16122 & ~n16125;
  assign n16127 = n14783 & ~n15219;
  assign n16128 = n15950 & n16114;
  assign n16129 = n16117 & n16128;
  assign n16130 = n16127 & n16129;
  assign n16131 = n15598 & n15750;
  assign n16132 = n16115 & n16131;
  assign n16133 = n14783 & n15219;
  assign n16134 = ~n15220 & ~n16133;
  assign n16135 = n16132 & ~n16134;
  assign n16136 = ~n16130 & ~n16135;
  assign n16137 = n16126 & n16136;
  assign n16138 = ~n15950 & n16114;
  assign n16139 = n15751 & n16138;
  assign n16140 = n15220 & n16139;
  assign n16141 = n16117 & n16138;
  assign n16142 = n16123 & n16138;
  assign n16143 = ~n16141 & ~n16142;
  assign n16144 = n16133 & ~n16143;
  assign n16145 = n16123 & n16128;
  assign n16146 = n15220 & n16145;
  assign n16147 = n15950 & ~n16114;
  assign n16148 = n15751 & n16147;
  assign n16149 = n16133 & n16148;
  assign n16150 = ~n16146 & ~n16149;
  assign n16151 = n16119 & ~n16132;
  assign n16152 = ~n16139 & n16151;
  assign n16153 = n16127 & ~n16152;
  assign n16154 = n16131 & n16147;
  assign n16155 = n16117 & n16147;
  assign n16156 = ~n16148 & ~n16155;
  assign n16157 = ~n16145 & n16156;
  assign n16158 = ~n16154 & n16157;
  assign n16159 = n16121 & ~n16158;
  assign n16160 = n16128 & n16131;
  assign n16161 = n16123 & n16147;
  assign n16162 = ~n16129 & ~n16161;
  assign n16163 = ~n16133 & n16162;
  assign n16164 = n15751 & n16128;
  assign n16165 = ~n16161 & ~n16164;
  assign n16166 = ~n15220 & n16165;
  assign n16167 = ~n16163 & ~n16166;
  assign n16168 = ~n16160 & ~n16167;
  assign n16169 = ~n16134 & ~n16168;
  assign n16170 = ~n16159 & ~n16169;
  assign n16171 = ~n16153 & n16170;
  assign n16172 = n16150 & n16171;
  assign n16173 = ~n16144 & n16172;
  assign n16174 = ~n16140 & n16173;
  assign n16175 = n16137 & n16174;
  assign n16176 = ~n16120 & n16175;
  assign n16177 = n15219 ^ n14783;
  assign n16178 = n16131 & n16138;
  assign n16179 = ~n16139 & ~n16178;
  assign n16180 = n16179 ^ n15219;
  assign n16181 = n16180 ^ n16179;
  assign n16182 = ~n16145 & ~n16160;
  assign n16183 = ~n16154 & n16182;
  assign n16184 = n16183 ^ n16179;
  assign n16185 = ~n16181 & n16184;
  assign n16186 = n16185 ^ n16179;
  assign n16187 = n16177 & ~n16186;
  assign n16188 = n16176 & ~n16187;
  assign n16189 = n16188 ^ n13824;
  assign n16190 = n16189 ^ x709;
  assign n16191 = n15143 & ~n15193;
  assign n16192 = ~n15150 & n15181;
  assign n16193 = n15149 & ~n16192;
  assign n16194 = ~n16191 & ~n16193;
  assign n16195 = n15164 & n15179;
  assign n16196 = n15180 & ~n15204;
  assign n16197 = n15152 & ~n16196;
  assign n16198 = ~n16195 & ~n16197;
  assign n16199 = ~n15184 & ~n15190;
  assign n16200 = n14959 & ~n16199;
  assign n16201 = n14959 & n15203;
  assign n16202 = n15152 & ~n15161;
  assign n16203 = ~n16201 & ~n16202;
  assign n16204 = ~n15144 & n16203;
  assign n16205 = ~n15176 & ~n15184;
  assign n16206 = n15152 & ~n16205;
  assign n16207 = ~n15147 & n15192;
  assign n16208 = n15149 & ~n16207;
  assign n16209 = ~n16206 & ~n16208;
  assign n16210 = n15176 & ~n15193;
  assign n16211 = ~n15150 & ~n15169;
  assign n16212 = n14959 & ~n16211;
  assign n16213 = n15186 & ~n15191;
  assign n16214 = n15164 & ~n16213;
  assign n16215 = ~n16212 & ~n16214;
  assign n16216 = ~n16210 & n16215;
  assign n16217 = n16209 & n16216;
  assign n16218 = n16204 & n16217;
  assign n16219 = ~n16200 & n16218;
  assign n16220 = n16198 & n16219;
  assign n16221 = n16194 & n16220;
  assign n16222 = n15175 & n16221;
  assign n16223 = n16222 ^ n12092;
  assign n16224 = n16223 ^ x657;
  assign n16225 = n13460 ^ x616;
  assign n16226 = n15837 ^ x621;
  assign n16227 = n16225 & ~n16226;
  assign n16228 = n14099 & ~n14122;
  assign n16229 = ~n14103 & ~n14123;
  assign n16230 = n14108 & ~n16229;
  assign n16231 = ~n16228 & ~n16230;
  assign n16232 = n14081 & ~n15465;
  assign n16233 = ~n14124 & n15461;
  assign n16234 = ~n14085 & n16233;
  assign n16235 = n14097 & ~n16234;
  assign n16236 = ~n15470 & n15978;
  assign n16237 = n14089 & ~n16236;
  assign n16238 = n14114 & ~n15470;
  assign n16239 = ~n14116 & n16238;
  assign n16240 = n14108 & ~n16239;
  assign n16241 = ~n16237 & ~n16240;
  assign n16242 = ~n14110 & n14131;
  assign n16243 = n14081 & ~n16242;
  assign n16244 = ~n14087 & n16229;
  assign n16245 = ~n14099 & n16244;
  assign n16246 = n14089 & ~n16245;
  assign n16247 = ~n14044 & n16238;
  assign n16248 = n14097 & ~n16247;
  assign n16249 = ~n16246 & ~n16248;
  assign n16250 = ~n16243 & n16249;
  assign n16251 = n16241 & n16250;
  assign n16252 = ~n16235 & n16251;
  assign n16253 = ~n16232 & n16252;
  assign n16254 = n16231 & n16253;
  assign n16255 = n15456 & n16254;
  assign n16256 = n16255 ^ n12417;
  assign n16257 = n16256 ^ x618;
  assign n16258 = n14820 & n14947;
  assign n16259 = ~n14879 & n15273;
  assign n16260 = n14889 & ~n16259;
  assign n16261 = ~n14887 & n14898;
  assign n16262 = ~n14916 & n16261;
  assign n16263 = n14821 & ~n16262;
  assign n16264 = ~n16260 & ~n16263;
  assign n16265 = ~n16258 & n16264;
  assign n16266 = n14918 & n15655;
  assign n16267 = ~n14943 & n16266;
  assign n16268 = n16267 ^ n14820;
  assign n16269 = n16268 ^ n16267;
  assign n16270 = ~n14896 & ~n15263;
  assign n16271 = n16270 ^ n16267;
  assign n16272 = ~n16269 & n16271;
  assign n16273 = n16272 ^ n16267;
  assign n16274 = ~n14819 & ~n16273;
  assign n16275 = n16265 & ~n16274;
  assign n16276 = ~n15651 & n16275;
  assign n16277 = n15649 & n16276;
  assign n16278 = n15253 & n16277;
  assign n16279 = ~n15251 & n16278;
  assign n16280 = n16279 ^ n12469;
  assign n16281 = n16280 ^ x619;
  assign n16282 = n15759 ^ x620;
  assign n16283 = n14735 ^ x617;
  assign n16284 = n16282 & ~n16283;
  assign n16285 = ~n16281 & n16284;
  assign n16286 = n16257 & n16285;
  assign n16287 = n16227 & n16286;
  assign n16288 = n16225 & n16226;
  assign n16289 = ~n16257 & n16281;
  assign n16290 = n16282 & n16283;
  assign n16291 = n16289 & n16290;
  assign n16292 = n16288 & n16291;
  assign n16293 = ~n16225 & n16226;
  assign n16294 = n16257 & n16281;
  assign n16295 = ~n16282 & ~n16283;
  assign n16296 = n16294 & n16295;
  assign n16297 = n16293 & n16296;
  assign n16298 = ~n16225 & ~n16226;
  assign n16299 = n16257 & ~n16281;
  assign n16300 = ~n16282 & n16283;
  assign n16301 = n16299 & n16300;
  assign n16302 = ~n16291 & ~n16301;
  assign n16303 = n16298 & ~n16302;
  assign n16304 = ~n16297 & ~n16303;
  assign n16305 = ~n16292 & n16304;
  assign n16306 = n16284 & n16289;
  assign n16307 = ~n16257 & ~n16281;
  assign n16308 = n16295 & n16307;
  assign n16309 = ~n16306 & ~n16308;
  assign n16310 = n16293 & ~n16309;
  assign n16311 = n16300 & n16307;
  assign n16312 = n16227 & n16311;
  assign n16313 = n16284 & n16294;
  assign n16314 = n16288 & n16313;
  assign n16315 = ~n16312 & ~n16314;
  assign n16316 = n16290 & n16299;
  assign n16317 = n16294 & n16300;
  assign n16318 = n16289 & n16300;
  assign n16319 = ~n16291 & ~n16318;
  assign n16320 = ~n16257 & n16285;
  assign n16321 = n16319 & ~n16320;
  assign n16322 = ~n16317 & n16321;
  assign n16323 = ~n16316 & n16322;
  assign n16324 = n16293 & ~n16323;
  assign n16325 = n16290 & n16294;
  assign n16326 = ~n16318 & ~n16325;
  assign n16327 = n16295 & n16299;
  assign n16328 = ~n16313 & ~n16327;
  assign n16329 = ~n16306 & n16328;
  assign n16330 = n16326 & n16329;
  assign n16331 = n16227 & ~n16330;
  assign n16332 = ~n16296 & ~n16311;
  assign n16333 = n16298 & ~n16332;
  assign n16334 = n16289 & n16295;
  assign n16335 = ~n16308 & ~n16334;
  assign n16336 = n16288 & ~n16335;
  assign n16337 = ~n16333 & ~n16336;
  assign n16338 = ~n16285 & n16337;
  assign n16339 = ~n16301 & n16338;
  assign n16340 = n16288 & ~n16339;
  assign n16341 = ~n16331 & ~n16340;
  assign n16342 = ~n16324 & n16341;
  assign n16345 = n16290 & n16307;
  assign n16343 = ~n16317 & n16338;
  assign n16344 = ~n16325 & n16343;
  assign n16346 = n16345 ^ n16344;
  assign n16347 = n16346 ^ n16345;
  assign n16348 = n16345 ^ n16226;
  assign n16349 = n16348 ^ n16345;
  assign n16350 = ~n16347 & ~n16349;
  assign n16351 = n16350 ^ n16345;
  assign n16352 = ~n16225 & n16351;
  assign n16353 = n16352 ^ n16345;
  assign n16354 = n16342 & ~n16353;
  assign n16355 = n16315 & n16354;
  assign n16356 = ~n16310 & n16355;
  assign n16357 = n16305 & n16356;
  assign n16358 = ~n16287 & n16357;
  assign n16359 = n16358 ^ n12597;
  assign n16360 = n16359 ^ x652;
  assign n16361 = ~n16224 & ~n16360;
  assign n16362 = n15523 & n15538;
  assign n16363 = ~n15526 & ~n16362;
  assign n16364 = n15552 & ~n16363;
  assign n16365 = n15289 & ~n15568;
  assign n16366 = ~n16364 & ~n16365;
  assign n16367 = ~n15564 & n15566;
  assign n16368 = ~n15575 & ~n15577;
  assign n16369 = n15519 & n15530;
  assign n16370 = ~n15545 & ~n16369;
  assign n16371 = n15568 & n16370;
  assign n16372 = n16368 & n16371;
  assign n16373 = n15552 & ~n16372;
  assign n16374 = ~n16367 & ~n16373;
  assign n16375 = ~n15539 & ~n15575;
  assign n16376 = ~n16369 & n16375;
  assign n16377 = n15289 & ~n16376;
  assign n16378 = n15546 & ~n16362;
  assign n16379 = ~n15524 & n16378;
  assign n16380 = n15568 & n16379;
  assign n16381 = n15529 & ~n16380;
  assign n16382 = ~n16377 & ~n16381;
  assign n16383 = n16374 & n16382;
  assign n16384 = n15536 & n16383;
  assign n16385 = n16366 & n16384;
  assign n16386 = n16385 ^ n13230;
  assign n16387 = n16386 ^ x656;
  assign n16388 = n15890 & ~n15901;
  assign n16389 = n15882 & n15917;
  assign n16390 = ~n15920 & n15938;
  assign n16391 = n15762 & ~n16390;
  assign n16392 = ~n16389 & ~n16391;
  assign n16393 = ~n16388 & n16392;
  assign n16394 = n15909 ^ n15900;
  assign n16395 = n16394 ^ n15900;
  assign n16396 = n15900 ^ n15761;
  assign n16397 = n16396 ^ n15900;
  assign n16398 = ~n16395 & n16397;
  assign n16399 = n16398 ^ n15900;
  assign n16400 = ~n15760 & n16399;
  assign n16401 = n16400 ^ n15900;
  assign n16402 = n15905 ^ n15898;
  assign n16403 = n15905 ^ n15762;
  assign n16404 = n16403 ^ n15762;
  assign n16405 = n15914 ^ n15762;
  assign n16406 = ~n16404 & n16405;
  assign n16407 = n16406 ^ n15762;
  assign n16408 = n16402 & n16407;
  assign n16409 = n16408 ^ n15898;
  assign n16410 = ~n16401 & ~n16409;
  assign n16411 = ~n15908 & ~n15931;
  assign n16412 = n15882 & ~n16411;
  assign n16413 = ~n15907 & ~n15913;
  assign n16414 = n16413 ^ n15762;
  assign n16415 = n16414 ^ n16413;
  assign n16416 = ~n15929 & ~n15935;
  assign n16417 = n16416 ^ n16413;
  assign n16418 = ~n16415 & n16417;
  assign n16419 = n16418 ^ n16413;
  assign n16420 = ~n16412 & n16419;
  assign n16421 = n16410 & n16420;
  assign n16422 = n15924 & n16421;
  assign n16423 = n16393 & n16422;
  assign n16424 = n15889 & n16423;
  assign n16425 = n16424 ^ n13382;
  assign n16426 = n16425 ^ x655;
  assign n16427 = ~n16387 & n16426;
  assign n16428 = n14760 & n14769;
  assign n16429 = n14602 ^ n14433;
  assign n16430 = n16429 ^ n14433;
  assign n16431 = n14751 ^ n14433;
  assign n16432 = n16431 ^ n14433;
  assign n16433 = ~n16430 & ~n16432;
  assign n16434 = n16433 ^ n14433;
  assign n16435 = ~n14736 & n16434;
  assign n16436 = n16435 ^ n14433;
  assign n16437 = ~n16428 & ~n16436;
  assign n16438 = n14737 & ~n14767;
  assign n16439 = n14753 & n14777;
  assign n16440 = ~n16438 & ~n16439;
  assign n16441 = n16437 & n16440;
  assign n16442 = n16441 ^ n12805;
  assign n16443 = n16442 ^ x654;
  assign n16444 = n16051 & n16053;
  assign n16445 = n16048 & n16091;
  assign n16446 = ~n16444 & ~n16445;
  assign n16447 = n16048 & n16080;
  assign n16448 = n16064 & ~n16447;
  assign n16449 = ~n16078 & n16084;
  assign n16450 = ~n16041 & n16095;
  assign n16451 = n16053 & ~n16450;
  assign n16452 = ~n16449 & ~n16451;
  assign n16453 = n16043 & n16072;
  assign n16454 = ~n16041 & ~n16069;
  assign n16455 = ~n16099 & n16454;
  assign n16456 = ~n16085 & n16455;
  assign n16457 = n16048 & ~n16456;
  assign n16458 = n16081 & n16102;
  assign n16459 = ~n16091 & n16458;
  assign n16460 = n16043 & ~n16459;
  assign n16461 = ~n16061 & n16102;
  assign n16462 = ~n16045 & n16461;
  assign n16463 = n15971 & ~n16462;
  assign n16464 = ~n16460 & ~n16463;
  assign n16465 = ~n16457 & n16464;
  assign n16466 = ~n16453 & n16465;
  assign n16467 = n16452 & n16466;
  assign n16468 = n16448 & n16467;
  assign n16469 = ~n16071 & n16468;
  assign n16470 = n16446 & n16469;
  assign n16471 = n16058 & n16470;
  assign n16472 = n16471 ^ n13003;
  assign n16473 = n16472 ^ x653;
  assign n16474 = ~n16443 & ~n16473;
  assign n16475 = n16427 & n16474;
  assign n16476 = n16361 & n16475;
  assign n16477 = ~n16224 & n16360;
  assign n16478 = n16224 & ~n16360;
  assign n16479 = ~n16477 & ~n16478;
  assign n16480 = n16387 & n16426;
  assign n16481 = n16474 & n16480;
  assign n16482 = ~n16387 & ~n16426;
  assign n16483 = n16474 & n16482;
  assign n16484 = ~n16481 & ~n16483;
  assign n16485 = n16479 & ~n16484;
  assign n16486 = n16387 & ~n16426;
  assign n16487 = n16443 & ~n16473;
  assign n16488 = n16486 & n16487;
  assign n16489 = n16482 & n16487;
  assign n16490 = n16427 & n16487;
  assign n16491 = n16474 & n16486;
  assign n16492 = ~n16490 & ~n16491;
  assign n16493 = ~n16489 & n16492;
  assign n16494 = ~n16488 & n16493;
  assign n16495 = n16477 & ~n16494;
  assign n16496 = ~n16485 & ~n16495;
  assign n16497 = n16443 & n16473;
  assign n16498 = n16427 & n16497;
  assign n16499 = ~n16443 & n16473;
  assign n16500 = ~n16387 & n16499;
  assign n16501 = n16480 & n16497;
  assign n16502 = ~n16500 & ~n16501;
  assign n16503 = ~n16498 & n16502;
  assign n16504 = n16478 & ~n16503;
  assign n16505 = n16224 & n16360;
  assign n16506 = n16482 & n16497;
  assign n16507 = ~n16490 & ~n16506;
  assign n16508 = n16505 & ~n16507;
  assign n16509 = ~n16504 & ~n16508;
  assign n16510 = n16480 & n16487;
  assign n16511 = n16361 & n16510;
  assign n16512 = n16486 & n16499;
  assign n16513 = n16361 & n16512;
  assign n16514 = n16486 & n16497;
  assign n16515 = n16361 & n16514;
  assign n16516 = ~n16513 & ~n16515;
  assign n16517 = ~n16498 & ~n16501;
  assign n16518 = n16361 & ~n16517;
  assign n16519 = n16480 & n16499;
  assign n16520 = ~n16498 & ~n16519;
  assign n16521 = ~n16512 & n16520;
  assign n16522 = ~n16514 & n16521;
  assign n16523 = n16505 & ~n16522;
  assign n16524 = ~n16518 & ~n16523;
  assign n16525 = n16502 & ~n16519;
  assign n16526 = n16477 & ~n16525;
  assign n16527 = ~n16475 & ~n16488;
  assign n16528 = ~n16489 & n16527;
  assign n16529 = ~n16491 & n16528;
  assign n16530 = n16478 & ~n16529;
  assign n16531 = ~n16526 & ~n16530;
  assign n16532 = n16524 & n16531;
  assign n16533 = n16516 & n16532;
  assign n16534 = ~n16511 & n16533;
  assign n16535 = n16509 & n16534;
  assign n16536 = n16496 & n16535;
  assign n16537 = ~n16476 & n16536;
  assign n16538 = n16537 ^ n13460;
  assign n16539 = n16538 ^ x710;
  assign n16540 = n15143 & n15149;
  assign n16541 = n14958 & ~n15180;
  assign n16542 = ~n16540 & ~n16541;
  assign n16543 = n15152 & n15169;
  assign n16544 = ~n15203 & n16192;
  assign n16545 = n15164 & ~n16544;
  assign n16546 = ~n16543 & ~n16545;
  assign n16547 = ~n15160 & n16205;
  assign n16548 = n14959 & ~n16547;
  assign n16549 = ~n15193 & ~n16205;
  assign n16550 = n15152 & n15157;
  assign n16551 = ~n15150 & ~n15204;
  assign n16552 = ~n15178 & n16551;
  assign n16553 = n14959 & ~n16552;
  assign n16554 = ~n16550 & ~n16553;
  assign n16555 = ~n16549 & n16554;
  assign n16556 = n15186 ^ n14958;
  assign n16557 = n16556 ^ n15186;
  assign n16558 = n15192 ^ n15186;
  assign n16559 = ~n16557 & n16558;
  assign n16560 = n16559 ^ n15186;
  assign n16561 = ~n15193 & ~n16560;
  assign n16562 = n16555 & ~n16561;
  assign n16563 = ~n15144 & n16562;
  assign n16564 = ~n16548 & n16563;
  assign n16565 = n16546 & n16564;
  assign n16566 = n16542 & n16565;
  assign n16567 = n15155 & n16566;
  assign n16568 = n16567 ^ n14316;
  assign n16569 = n16568 ^ x666;
  assign n16570 = n15882 & n15920;
  assign n16571 = n15890 & n15926;
  assign n16572 = ~n16570 & ~n16571;
  assign n16573 = n15884 & n15899;
  assign n16574 = n15938 & n16416;
  assign n16575 = n15898 & ~n16574;
  assign n16576 = ~n16573 & ~n16575;
  assign n16577 = ~n15892 & n15909;
  assign n16578 = n15762 & ~n16577;
  assign n16579 = ~n15880 & ~n15905;
  assign n16580 = n15898 & ~n16579;
  assign n16581 = n15909 & ~n15913;
  assign n16582 = ~n15929 & n16581;
  assign n16583 = n15882 & ~n16582;
  assign n16584 = ~n16580 & ~n16583;
  assign n16585 = ~n16578 & n16584;
  assign n16586 = n16576 & n16585;
  assign n16587 = n16572 & n16586;
  assign n16588 = n16393 & n16587;
  assign n16589 = ~n15911 & n16588;
  assign n16590 = n15903 & n16589;
  assign n16591 = n16590 ^ n14288;
  assign n16592 = n16591 ^ x667;
  assign n16593 = ~n16569 & ~n16592;
  assign n16594 = n14427 ^ n14147;
  assign n16595 = ~n13461 & n16594;
  assign n16596 = ~n14750 & ~n16595;
  assign n16597 = n14763 & ~n16596;
  assign n16598 = n14771 ^ n13461;
  assign n16599 = n16598 ^ n13461;
  assign n16600 = ~n14772 & ~n16599;
  assign n16601 = n16600 ^ n13461;
  assign n16602 = ~n13825 & ~n16601;
  assign n16603 = n16602 ^ n14771;
  assign n16604 = n14753 & ~n16603;
  assign n16605 = ~n16597 & ~n16604;
  assign n16606 = ~n13461 & ~n14765;
  assign n16607 = n14742 ^ n14147;
  assign n16608 = n16607 ^ n14742;
  assign n16609 = n14427 ^ n13825;
  assign n16610 = n14754 & ~n16609;
  assign n16611 = n16610 ^ n16609;
  assign n16612 = n16611 ^ n14742;
  assign n16613 = ~n16608 & ~n16612;
  assign n16614 = n16613 ^ n14742;
  assign n16615 = ~n16606 & ~n16614;
  assign n16616 = n14769 & n16615;
  assign n16617 = n13825 & ~n14738;
  assign n16618 = n14427 & n14764;
  assign n16619 = ~n16617 & ~n16618;
  assign n16620 = ~n14147 & ~n16611;
  assign n16621 = n16619 & ~n16620;
  assign n16622 = n14737 & ~n16621;
  assign n16623 = ~n16616 & ~n16622;
  assign n16624 = n16605 & n16623;
  assign n16625 = n16624 ^ n14263;
  assign n16626 = n16625 ^ x668;
  assign n16627 = n15971 & n16071;
  assign n16628 = n16053 & n16073;
  assign n16629 = ~n16627 & ~n16628;
  assign n16630 = n16450 & n16461;
  assign n16631 = ~n16051 & n16630;
  assign n16632 = n16043 & ~n16631;
  assign n16633 = n15970 ^ n15951;
  assign n16635 = ~n16084 & n16095;
  assign n16634 = n16081 & n16454;
  assign n16636 = n16635 ^ n16634;
  assign n16637 = n16635 ^ n15970;
  assign n16638 = n16637 ^ n16635;
  assign n16639 = n16636 & n16638;
  assign n16640 = n16639 ^ n16635;
  assign n16641 = ~n16633 & ~n16640;
  assign n16642 = ~n16632 & ~n16641;
  assign n16643 = ~n16078 & n16099;
  assign n16644 = n16075 & n16086;
  assign n16645 = ~n16098 & n16644;
  assign n16646 = n16048 & ~n16645;
  assign n16647 = ~n16643 & ~n16646;
  assign n16648 = n16642 & n16647;
  assign n16649 = n16629 & n16648;
  assign n16650 = ~n16066 & n16649;
  assign n16651 = n16448 & n16650;
  assign n16652 = n16047 & n16651;
  assign n16653 = n16446 & n16652;
  assign n16654 = n16653 ^ n14348;
  assign n16655 = n16654 ^ x665;
  assign n16656 = ~n16626 & ~n16655;
  assign n16657 = n16593 & n16656;
  assign n16658 = n16015 ^ x639;
  assign n16659 = n15485 ^ x634;
  assign n16660 = n16658 & ~n16659;
  assign n16661 = n13406 & n14985;
  assign n16662 = n12599 & ~n16661;
  assign n16663 = n13390 & ~n13414;
  assign n16664 = ~n13405 & n16663;
  assign n16665 = n13398 & ~n16664;
  assign n16666 = ~n16662 & ~n16665;
  assign n16667 = n13434 & ~n14963;
  assign n16668 = n13393 & ~n15230;
  assign n16669 = ~n16667 & ~n16668;
  assign n16670 = n16666 & n16669;
  assign n16671 = n15226 & n16670;
  assign n16672 = n15223 & n16671;
  assign n16673 = n14970 & n16672;
  assign n16674 = ~n13413 & n16673;
  assign n16675 = ~n13411 & n16674;
  assign n16676 = n16675 ^ n13919;
  assign n16677 = n16676 ^ x636;
  assign n16678 = n15287 ^ x635;
  assign n16679 = ~n16677 & n16678;
  assign n16680 = n14678 & ~n14686;
  assign n16681 = n14789 & n15788;
  assign n16682 = ~n14705 & n16681;
  assign n16683 = n14672 & ~n16682;
  assign n16684 = ~n16680 & ~n16683;
  assign n16685 = n14668 & ~n15790;
  assign n16686 = ~n14670 & ~n14698;
  assign n16687 = n14603 & ~n16686;
  assign n16688 = ~n14703 & n14720;
  assign n16689 = n14605 & ~n16688;
  assign n16690 = ~n16687 & ~n16689;
  assign n16691 = ~n16685 & n16690;
  assign n16692 = n16684 & n16691;
  assign n16693 = n15769 & n16692;
  assign n16694 = ~n15765 & n16693;
  assign n16695 = ~n14682 & n16694;
  assign n16696 = n14788 & n16695;
  assign n16697 = n16696 ^ n13949;
  assign n16698 = n16697 ^ x637;
  assign n16699 = n15969 ^ x638;
  assign n16700 = n16698 & ~n16699;
  assign n16701 = n16679 & n16700;
  assign n16702 = n16698 & n16699;
  assign n16703 = n16677 & n16678;
  assign n16704 = n16702 & n16703;
  assign n16705 = ~n16701 & ~n16704;
  assign n16706 = n16660 & ~n16705;
  assign n16707 = n16658 & n16659;
  assign n16708 = ~n16698 & n16699;
  assign n16709 = n16677 & ~n16678;
  assign n16710 = n16708 & n16709;
  assign n16711 = ~n16698 & ~n16699;
  assign n16712 = ~n16677 & ~n16678;
  assign n16713 = n16711 & n16712;
  assign n16714 = ~n16710 & ~n16713;
  assign n16715 = n16707 & ~n16714;
  assign n16716 = ~n16706 & ~n16715;
  assign n16717 = n16703 & n16708;
  assign n16718 = n16703 & n16711;
  assign n16719 = ~n16717 & ~n16718;
  assign n16720 = n16660 & ~n16719;
  assign n16721 = ~n16658 & n16659;
  assign n16722 = n16700 & n16709;
  assign n16723 = ~n16710 & ~n16722;
  assign n16724 = n16702 & n16709;
  assign n16725 = n16700 & n16712;
  assign n16726 = ~n16724 & ~n16725;
  assign n16727 = n16723 & n16726;
  assign n16728 = n16721 & ~n16727;
  assign n16729 = n16701 & n16721;
  assign n16730 = n16679 & n16708;
  assign n16731 = n16730 ^ n16707;
  assign n16732 = n16730 ^ n16721;
  assign n16733 = n16732 ^ n16721;
  assign n16734 = n16722 ^ n16721;
  assign n16735 = ~n16733 & ~n16734;
  assign n16736 = n16735 ^ n16721;
  assign n16737 = n16731 & n16736;
  assign n16738 = n16737 ^ n16707;
  assign n16740 = ~n16658 & ~n16659;
  assign n16739 = n16679 & n16711;
  assign n16741 = n16740 ^ n16739;
  assign n16742 = n16659 ^ n16658;
  assign n16743 = n16742 ^ n16717;
  assign n16744 = n16742 ^ n16739;
  assign n16745 = n16744 ^ n16742;
  assign n16746 = ~n16743 & ~n16745;
  assign n16747 = n16746 ^ n16742;
  assign n16748 = n16741 & n16747;
  assign n16749 = n16748 ^ n16740;
  assign n16750 = ~n16738 & ~n16749;
  assign n16751 = ~n16707 & ~n16740;
  assign n16752 = n16700 & n16703;
  assign n16753 = n16679 & n16702;
  assign n16754 = ~n16752 & ~n16753;
  assign n16755 = ~n16751 & ~n16754;
  assign n16756 = n16702 & n16712;
  assign n16757 = ~n16724 & ~n16756;
  assign n16758 = n16660 & ~n16757;
  assign n16759 = ~n16755 & ~n16758;
  assign n16760 = n16750 & n16759;
  assign n16761 = n16704 ^ n16659;
  assign n16762 = n16761 ^ n16704;
  assign n16763 = n16709 & n16711;
  assign n16764 = n16763 ^ n16704;
  assign n16765 = ~n16762 & n16764;
  assign n16766 = n16765 ^ n16704;
  assign n16767 = n16742 & n16766;
  assign n16768 = n16760 & ~n16767;
  assign n16769 = ~n16729 & n16768;
  assign n16770 = ~n16728 & n16769;
  assign n16771 = ~n16720 & n16770;
  assign n16772 = ~n16725 & ~n16763;
  assign n16773 = n16772 ^ n16740;
  assign n16774 = n16772 ^ n16707;
  assign n16775 = n16774 ^ n16707;
  assign n16776 = n16708 & n16712;
  assign n16777 = ~n16756 & ~n16776;
  assign n16778 = n16777 ^ n16707;
  assign n16779 = n16775 & n16778;
  assign n16780 = n16779 ^ n16707;
  assign n16781 = ~n16773 & n16780;
  assign n16782 = n16781 ^ n16740;
  assign n16783 = n16771 & ~n16782;
  assign n16784 = n16716 & n16783;
  assign n16785 = n16784 ^ n14216;
  assign n16786 = n16785 ^ x669;
  assign n16787 = n15601 & n15720;
  assign n16788 = ~n15706 & ~n15722;
  assign n16789 = n15694 & ~n16788;
  assign n16790 = ~n16787 & ~n16789;
  assign n16791 = ~n15703 & ~n15715;
  assign n16792 = n15601 & ~n16791;
  assign n16793 = n15694 & n15714;
  assign n16794 = ~n15702 & n15723;
  assign n16795 = ~n16793 & ~n16794;
  assign n16796 = ~n15729 & ~n15734;
  assign n16797 = ~n15706 & n16796;
  assign n16798 = n15709 & ~n16797;
  assign n16799 = n15694 & n15718;
  assign n16800 = n15601 & ~n16796;
  assign n16801 = ~n16799 & ~n16800;
  assign n16802 = n15695 & n15705;
  assign n16803 = ~n15714 & ~n16802;
  assign n16804 = n15702 & ~n16803;
  assign n16805 = ~n15696 & ~n15715;
  assign n16806 = ~n15720 & n16805;
  assign n16807 = n16806 ^ n15600;
  assign n16808 = n16807 ^ n16806;
  assign n16809 = ~n15696 & ~n15703;
  assign n16810 = n15736 & n16809;
  assign n16811 = ~n15698 & n16810;
  assign n16812 = n16811 ^ n16806;
  assign n16813 = n16808 & n16812;
  assign n16814 = n16813 ^ n16806;
  assign n16815 = n15599 & ~n16814;
  assign n16816 = ~n16804 & ~n16815;
  assign n16817 = n16801 & n16816;
  assign n16818 = ~n16798 & n16817;
  assign n16819 = n16795 & n16818;
  assign n16820 = ~n16792 & n16819;
  assign n16821 = ~n15701 & n16820;
  assign n16822 = n16790 & n16821;
  assign n16823 = ~n15692 & n16822;
  assign n16824 = ~n15685 & n16823;
  assign n16825 = n16824 ^ n14183;
  assign n16826 = n16825 ^ x664;
  assign n16827 = ~n16786 & ~n16826;
  assign n16828 = n16657 & n16827;
  assign n16829 = n16786 & ~n16826;
  assign n16830 = n16626 & ~n16655;
  assign n16831 = n16569 & n16830;
  assign n16832 = n16592 & n16831;
  assign n16833 = n16829 & n16832;
  assign n16834 = ~n16828 & ~n16833;
  assign n16835 = n16626 & n16655;
  assign n16836 = n16593 & n16835;
  assign n16837 = n16829 & n16836;
  assign n16838 = ~n16569 & n16830;
  assign n16839 = n16786 & n16826;
  assign n16840 = ~n16827 & ~n16839;
  assign n16841 = n16838 & ~n16840;
  assign n16842 = n16592 & n16841;
  assign n16843 = ~n16837 & ~n16842;
  assign n16844 = n16569 & n16592;
  assign n16845 = ~n16626 & n16655;
  assign n16846 = n16844 & n16845;
  assign n16847 = ~n16569 & n16592;
  assign n16848 = n16835 & n16847;
  assign n16849 = ~n16846 & ~n16848;
  assign n16850 = n16829 & ~n16849;
  assign n16851 = ~n16786 & n16826;
  assign n16852 = ~n16592 & n16838;
  assign n16853 = n16569 & ~n16592;
  assign n16854 = n16656 & n16853;
  assign n16855 = ~n16832 & ~n16854;
  assign n16856 = ~n16852 & n16855;
  assign n16857 = ~n16836 & n16856;
  assign n16858 = n16851 & ~n16857;
  assign n16859 = n16656 & n16847;
  assign n16860 = ~n16854 & ~n16859;
  assign n16861 = ~n16829 & ~n16839;
  assign n16862 = ~n16860 & ~n16861;
  assign n16863 = ~n16831 & ~n16838;
  assign n16864 = n16829 & ~n16863;
  assign n16865 = ~n16592 & n16864;
  assign n16866 = ~n16862 & ~n16865;
  assign n16867 = n16845 & n16847;
  assign n16868 = ~n16848 & ~n16867;
  assign n16869 = n16835 & n16853;
  assign n16870 = ~n16846 & ~n16869;
  assign n16871 = n16868 & n16870;
  assign n16872 = n16851 & ~n16871;
  assign n16873 = n16593 & n16845;
  assign n16874 = n16835 & n16844;
  assign n16875 = n16845 & n16853;
  assign n16876 = ~n16874 & ~n16875;
  assign n16877 = ~n16836 & n16876;
  assign n16878 = ~n16827 & n16877;
  assign n16879 = ~n16867 & ~n16874;
  assign n16880 = ~n16869 & n16879;
  assign n16881 = ~n16839 & n16880;
  assign n16882 = ~n16878 & ~n16881;
  assign n16883 = ~n16873 & ~n16882;
  assign n16884 = ~n16840 & ~n16883;
  assign n16885 = ~n16872 & ~n16884;
  assign n16886 = n16656 & n16844;
  assign n16887 = n16886 ^ n16827;
  assign n16888 = ~n16592 & n16831;
  assign n16889 = n16888 ^ n16839;
  assign n16890 = n16839 ^ n16827;
  assign n16891 = n16890 ^ n16839;
  assign n16892 = ~n16889 & n16891;
  assign n16893 = n16892 ^ n16839;
  assign n16894 = n16887 & ~n16893;
  assign n16895 = n16894 ^ n16886;
  assign n16896 = n16885 & ~n16895;
  assign n16897 = n16866 & n16896;
  assign n16898 = ~n16858 & n16897;
  assign n16899 = ~n16850 & n16898;
  assign n16900 = n16843 & n16899;
  assign n16901 = n16834 & n16900;
  assign n16902 = n16901 ^ n14426;
  assign n16903 = n16902 ^ x708;
  assign n16904 = ~n16539 & ~n16903;
  assign n16905 = ~n16190 & n16904;
  assign n16906 = n15529 & n15575;
  assign n16907 = n15524 & n15566;
  assign n16908 = ~n16906 & ~n16907;
  assign n16909 = ~n15544 & n15549;
  assign n16910 = n15552 & ~n16909;
  assign n16911 = n15530 & n15537;
  assign n16912 = ~n15532 & ~n16911;
  assign n16913 = n16368 & n16912;
  assign n16914 = n15552 & ~n16913;
  assign n16915 = ~n16362 & ~n16369;
  assign n16916 = ~n15524 & ~n16911;
  assign n16917 = n16909 & n16916;
  assign n16918 = n16915 & n16917;
  assign n16919 = n15289 & ~n16918;
  assign n16920 = ~n16914 & ~n16919;
  assign n16923 = ~n15526 & ~n15531;
  assign n16921 = n15569 & ~n16362;
  assign n16922 = ~n15539 & n16921;
  assign n16924 = n16923 ^ n16922;
  assign n16925 = n16923 ^ n15574;
  assign n16926 = n16923 & ~n16925;
  assign n16927 = n16926 ^ n16923;
  assign n16928 = n16924 & n16927;
  assign n16929 = n16928 ^ n16926;
  assign n16930 = n16929 ^ n16923;
  assign n16931 = n16930 ^ n15574;
  assign n16932 = n16920 & ~n16931;
  assign n16933 = n16932 ^ n16920;
  assign n16934 = ~n16910 & n16933;
  assign n16935 = n16908 & n16934;
  assign n16936 = ~n15593 & n16935;
  assign n16937 = n16369 ^ n15567;
  assign n16938 = ~n15589 & n16937;
  assign n16939 = n16938 ^ n15567;
  assign n16940 = ~n15288 & n16939;
  assign n16941 = n16936 & ~n16940;
  assign n16942 = n16941 ^ n13863;
  assign n16943 = n16942 ^ x649;
  assign n16944 = n16359 ^ x650;
  assign n16945 = n16943 & n16944;
  assign n16946 = n16721 & n16730;
  assign n16947 = ~n16705 & n16740;
  assign n16948 = ~n16946 & ~n16947;
  assign n16949 = n16707 & ~n16754;
  assign n16950 = ~n16763 & ~n16776;
  assign n16951 = n16757 & n16950;
  assign n16952 = n16740 & ~n16951;
  assign n16953 = ~n16719 & ~n16751;
  assign n16954 = ~n16756 & n16950;
  assign n16955 = n16707 & ~n16954;
  assign n16956 = ~n16717 & ~n16739;
  assign n16957 = ~n16725 & ~n16752;
  assign n16958 = n16757 & n16957;
  assign n16959 = n16956 & n16958;
  assign n16960 = n16721 & ~n16959;
  assign n16961 = ~n16955 & ~n16960;
  assign n16962 = ~n16953 & n16961;
  assign n16963 = ~n16707 & ~n16721;
  assign n16964 = n16713 & ~n16963;
  assign n16965 = n16699 ^ n16677;
  assign n16966 = n16965 ^ n16678;
  assign n16967 = n16966 ^ n16678;
  assign n16968 = n16967 ^ n16966;
  assign n16969 = n16966 ^ n16699;
  assign n16970 = ~n16968 & n16969;
  assign n16971 = n16970 ^ n16966;
  assign n16972 = n16698 & ~n16971;
  assign n16973 = n16972 ^ n16966;
  assign n16974 = n16660 & ~n16973;
  assign n16975 = ~n16964 & ~n16974;
  assign n16976 = n16962 & n16975;
  assign n16977 = ~n16952 & n16976;
  assign n16978 = ~n16949 & n16977;
  assign n16979 = ~n16706 & n16978;
  assign n16980 = n16948 & n16979;
  assign n16981 = n16980 ^ n14040;
  assign n16982 = n16981 ^ x647;
  assign n16983 = ~n15723 & n16809;
  assign n16984 = ~n15734 & n16983;
  assign n16985 = n15709 & ~n16984;
  assign n16986 = ~n16792 & ~n16985;
  assign n16987 = n15601 & n15698;
  assign n16988 = n15688 & n15694;
  assign n16989 = ~n16987 & ~n16988;
  assign n16990 = n15599 & n15720;
  assign n16991 = n15686 & n15722;
  assign n16992 = ~n15706 & ~n15729;
  assign n16993 = ~n15688 & n16992;
  assign n16994 = n15601 & ~n16993;
  assign n16995 = ~n16991 & ~n16994;
  assign n16996 = ~n15691 & ~n16802;
  assign n16997 = n15709 & ~n16996;
  assign n16998 = n15718 ^ n15702;
  assign n16999 = n16998 ^ n15718;
  assign n17000 = n15717 & n15730;
  assign n17001 = n17000 ^ n15718;
  assign n17002 = ~n16999 & ~n17001;
  assign n17003 = n17002 ^ n15718;
  assign n17004 = ~n16997 & ~n17003;
  assign n17005 = n16995 & n17004;
  assign n17006 = ~n16990 & n17005;
  assign n17007 = n16989 & n17006;
  assign n17008 = n16790 & n17007;
  assign n17009 = n16986 & n17008;
  assign n17010 = ~n15692 & n17009;
  assign n17011 = n17010 ^ n13889;
  assign n17012 = n17011 ^ x648;
  assign n17013 = ~n16982 & ~n17012;
  assign n17014 = n16945 & n17013;
  assign n17015 = n16472 ^ x651;
  assign n17016 = n15898 & n15913;
  assign n17017 = n15887 & ~n15917;
  assign n17018 = ~n15920 & n17017;
  assign n17019 = n15890 & ~n17018;
  assign n17020 = ~n17016 & ~n17019;
  assign n17021 = ~n15926 & ~n15935;
  assign n17022 = ~n15899 & ~n17021;
  assign n17032 = ~n15908 & n15914;
  assign n17033 = n15890 & ~n17032;
  assign n17034 = ~n16570 & ~n17033;
  assign n17035 = ~n15929 & n17034;
  assign n17023 = ~n15929 & n16579;
  assign n17024 = ~n15898 & n17023;
  assign n17025 = ~n15905 & ~n15929;
  assign n17026 = n15762 & ~n17025;
  assign n17027 = ~n15895 & ~n17026;
  assign n17028 = ~n15880 & n17027;
  assign n17029 = ~n15917 & n17028;
  assign n17030 = ~n17024 & ~n17029;
  assign n17031 = ~n15900 & ~n17030;
  assign n17036 = n17035 ^ n17031;
  assign n17037 = ~n15899 & n17036;
  assign n17038 = n17037 ^ n17035;
  assign n17039 = ~n15888 & n17038;
  assign n17040 = ~n17022 & n17039;
  assign n17041 = n17020 & n17040;
  assign n17042 = n15909 ^ n15760;
  assign n17043 = n17042 ^ n15909;
  assign n17044 = n15938 ^ n15909;
  assign n17045 = n17043 & n17044;
  assign n17046 = n17045 ^ n15909;
  assign n17047 = ~n15761 & ~n17046;
  assign n17048 = n17041 & ~n17047;
  assign n17049 = n15916 & n17048;
  assign n17050 = n17049 ^ n14079;
  assign n17051 = n17050 ^ x646;
  assign n17052 = n17015 & n17051;
  assign n17053 = n17014 & n17052;
  assign n17054 = ~n16982 & n17012;
  assign n17055 = ~n16943 & n16944;
  assign n17056 = n17054 & n17055;
  assign n17057 = ~n17015 & n17051;
  assign n17058 = n17056 & n17057;
  assign n17059 = ~n17053 & ~n17058;
  assign n17060 = n16982 & n17012;
  assign n17061 = n16945 & n17060;
  assign n17062 = n17015 & ~n17051;
  assign n17063 = n17061 & n17062;
  assign n17064 = n17013 & n17055;
  assign n17065 = ~n17015 & ~n17051;
  assign n17066 = n17064 & n17065;
  assign n17067 = ~n17063 & ~n17066;
  assign n17068 = n17059 & n17067;
  assign n17069 = ~n16943 & ~n16944;
  assign n17070 = n17013 & n17069;
  assign n17071 = n17062 & n17070;
  assign n17072 = n17060 & n17069;
  assign n17073 = n17052 & n17072;
  assign n17074 = n17056 & n17062;
  assign n17075 = ~n17073 & ~n17074;
  assign n17076 = ~n17071 & n17075;
  assign n17077 = n16945 & n17054;
  assign n17078 = ~n17070 & ~n17077;
  assign n17079 = n17057 & ~n17078;
  assign n17080 = n16982 & ~n17012;
  assign n17081 = n17055 & n17080;
  assign n17082 = n17052 & n17081;
  assign n17083 = n16943 & ~n16944;
  assign n17084 = n17080 & n17083;
  assign n17085 = ~n17072 & ~n17081;
  assign n17086 = ~n17084 & n17085;
  assign n17087 = n17062 & ~n17086;
  assign n17088 = ~n17082 & ~n17087;
  assign n17089 = n17060 & n17083;
  assign n17090 = ~n17081 & ~n17089;
  assign n17091 = n17065 & ~n17090;
  assign n17092 = n17013 & n17083;
  assign n17093 = n17069 & n17080;
  assign n17094 = ~n17092 & ~n17093;
  assign n17095 = n17055 & n17060;
  assign n17096 = n16945 & n17080;
  assign n17097 = ~n17089 & ~n17096;
  assign n17098 = ~n17095 & n17097;
  assign n17099 = n17094 & n17098;
  assign n17100 = n17057 & ~n17099;
  assign n17101 = n17051 ^ n17015;
  assign n17108 = ~n17014 & ~n17092;
  assign n17102 = ~n17084 & ~n17095;
  assign n17103 = n17054 & n17083;
  assign n17104 = n17054 & n17069;
  assign n17105 = ~n17077 & ~n17104;
  assign n17106 = ~n17103 & n17105;
  assign n17107 = n17102 & n17106;
  assign n17109 = n17108 ^ n17107;
  assign n17110 = n17109 ^ n17107;
  assign n17111 = n17107 ^ n17051;
  assign n17112 = n17111 ^ n17107;
  assign n17113 = ~n17110 & ~n17112;
  assign n17114 = n17113 ^ n17107;
  assign n17115 = n17101 & ~n17114;
  assign n17116 = n17115 ^ n17107;
  assign n17117 = ~n17100 & n17116;
  assign n17118 = ~n17091 & n17117;
  assign n17119 = n17088 & n17118;
  assign n17120 = ~n17079 & n17119;
  assign n17121 = n17076 & n17120;
  assign n17122 = n17068 & n17121;
  assign n17123 = n17122 ^ n14146;
  assign n17124 = n17123 ^ x707;
  assign n17129 = n16539 ^ n16190;
  assign n17125 = ~n16539 & n16903;
  assign n17126 = n16190 & n17125;
  assign n17127 = n16539 & ~n16903;
  assign n17128 = ~n17126 & ~n17127;
  assign n17130 = n17129 ^ n17128;
  assign n17131 = ~n17124 & n17130;
  assign n17132 = n17131 ^ n17129;
  assign n17133 = ~n16905 & n17132;
  assign n17134 = n15949 ^ x681;
  assign n17135 = n15702 & n15706;
  assign n17136 = ~n15688 & n15730;
  assign n17137 = n15709 & ~n17136;
  assign n17138 = n15686 & ~n15725;
  assign n17139 = n15724 & n16796;
  assign n17140 = ~n15691 & n17139;
  assign n17141 = n15694 & ~n17140;
  assign n17142 = ~n17138 & ~n17141;
  assign n17143 = ~n17137 & n17142;
  assign n17144 = ~n17135 & n17143;
  assign n17145 = ~n15696 & ~n15734;
  assign n17146 = ~n15722 & n17145;
  assign n17147 = n17146 ^ n16803;
  assign n17148 = n17147 ^ n16803;
  assign n17149 = n16803 ^ n15600;
  assign n17150 = n17149 ^ n16803;
  assign n17151 = ~n17148 & n17150;
  assign n17152 = n17151 ^ n16803;
  assign n17153 = n15702 & ~n17152;
  assign n17154 = n17153 ^ n16803;
  assign n17155 = n17144 & n17154;
  assign n17156 = n16989 & n17155;
  assign n17157 = n16986 & n17156;
  assign n17158 = n15693 & n17157;
  assign n17159 = ~n15685 & n17158;
  assign n17160 = n17159 ^ n14456;
  assign n17161 = n17160 ^ x676;
  assign n17162 = n17134 & ~n17161;
  assign n17163 = n14763 & ~n16621;
  assign n17164 = n14753 & ~n16615;
  assign n17165 = ~n17163 & ~n17164;
  assign n17166 = n14736 ^ n14602;
  assign n17167 = n16596 ^ n14736;
  assign n17168 = n17167 ^ n16596;
  assign n17169 = n16603 ^ n16596;
  assign n17170 = ~n17168 & ~n17169;
  assign n17171 = n17170 ^ n16596;
  assign n17172 = n17166 & n17171;
  assign n17173 = n17165 & ~n17172;
  assign n17174 = n17173 ^ n14469;
  assign n17175 = n17174 ^ x678;
  assign n17176 = ~n16726 & n16740;
  assign n17177 = n16721 & ~n16951;
  assign n17178 = ~n17176 & ~n17177;
  assign n17179 = ~n16722 & ~n16776;
  assign n17180 = ~n16751 & ~n17179;
  assign n17181 = n16721 & ~n16956;
  assign n17182 = ~n16704 & ~n16718;
  assign n17183 = ~n16756 & n17182;
  assign n17184 = n16714 & n17183;
  assign n17185 = n16754 & n17184;
  assign n17186 = n16660 & ~n17185;
  assign n17188 = ~n16753 & n17182;
  assign n17187 = ~n16730 & n16956;
  assign n17189 = n17188 ^ n17187;
  assign n17190 = n17187 ^ n16659;
  assign n17191 = n16742 & ~n17190;
  assign n17192 = n17191 ^ n16659;
  assign n17193 = n17189 & ~n17192;
  assign n17194 = n17193 ^ n17188;
  assign n17195 = ~n16701 & n17194;
  assign n17196 = ~n16751 & ~n17195;
  assign n17197 = ~n17186 & ~n17196;
  assign n17198 = ~n17181 & n17197;
  assign n17199 = ~n16767 & n17198;
  assign n17200 = ~n16729 & n17199;
  assign n17201 = ~n17180 & n17200;
  assign n17202 = n17178 & n17201;
  assign n17203 = ~n16715 & n17202;
  assign n17204 = n17203 ^ n14539;
  assign n17205 = n17204 ^ x679;
  assign n17206 = n17175 & n17205;
  assign n17207 = n16288 & n16334;
  assign n17208 = n16227 & ~n16319;
  assign n17209 = ~n17207 & ~n17208;
  assign n17210 = n16293 & n16316;
  assign n17211 = n16298 & n16306;
  assign n17212 = n16227 & n16334;
  assign n17213 = ~n17211 & ~n17212;
  assign n17214 = ~n17210 & n17213;
  assign n17215 = n16227 & n16308;
  assign n17216 = ~n16320 & ~n16334;
  assign n17217 = n16298 & ~n17216;
  assign n17218 = ~n17215 & ~n17217;
  assign n17219 = n16298 & n16311;
  assign n17220 = ~n16317 & ~n16345;
  assign n17221 = ~n16313 & n17220;
  assign n17222 = n16227 & ~n17221;
  assign n17223 = ~n17219 & ~n17222;
  assign n17224 = ~n16311 & n17220;
  assign n17225 = n16329 & n17224;
  assign n17226 = n16293 & ~n17225;
  assign n17227 = ~n16316 & ~n16345;
  assign n17228 = ~n16301 & ~n16325;
  assign n17229 = n17227 & n17228;
  assign n17230 = n16298 & ~n17229;
  assign n17231 = n16323 & n16328;
  assign n17232 = n16288 & ~n17231;
  assign n17233 = ~n17230 & ~n17232;
  assign n17234 = ~n17226 & n17233;
  assign n17235 = n17223 & n17234;
  assign n17236 = ~n16297 & n17235;
  assign n17237 = n17218 & n17236;
  assign n17238 = n17214 & n17237;
  assign n17239 = n17209 & n17238;
  assign n17240 = ~n16287 & n17239;
  assign n17241 = n17240 ^ n14517;
  assign n17242 = n17241 ^ x677;
  assign n17243 = n15218 ^ x680;
  assign n17244 = ~n17242 & ~n17243;
  assign n17245 = n17206 & n17244;
  assign n17246 = n17162 & n17245;
  assign n17247 = ~n17175 & n17205;
  assign n17248 = n17244 & n17247;
  assign n17249 = ~n17242 & n17243;
  assign n17250 = n17175 & ~n17205;
  assign n17251 = n17249 & n17250;
  assign n17252 = ~n17248 & ~n17251;
  assign n17253 = n17162 & ~n17252;
  assign n17254 = ~n17246 & ~n17253;
  assign n17255 = ~n17175 & ~n17205;
  assign n17256 = n17249 & n17255;
  assign n17257 = n17162 & n17256;
  assign n17258 = n17134 & n17161;
  assign n17259 = n17242 & ~n17243;
  assign n17260 = n17206 & n17259;
  assign n17261 = n17247 & n17259;
  assign n17262 = n17242 & n17243;
  assign n17263 = n17250 & n17262;
  assign n17264 = ~n17261 & ~n17263;
  assign n17265 = ~n17260 & n17264;
  assign n17266 = n17258 & ~n17265;
  assign n17267 = ~n17257 & ~n17266;
  assign n17268 = n17161 ^ n17134;
  assign n17269 = n17255 & n17259;
  assign n17270 = ~n17268 & n17269;
  assign n17271 = ~n17134 & n17161;
  assign n17272 = n17247 & n17249;
  assign n17273 = n17244 & n17250;
  assign n17274 = ~n17272 & ~n17273;
  assign n17275 = n17206 & n17249;
  assign n17276 = n17255 & n17262;
  assign n17277 = ~n17275 & ~n17276;
  assign n17278 = ~n17245 & ~n17256;
  assign n17279 = n17264 & n17278;
  assign n17280 = n17277 & n17279;
  assign n17281 = n17274 & n17280;
  assign n17282 = n17271 & n17281;
  assign n17283 = n17250 & n17259;
  assign n17284 = n17277 & ~n17283;
  assign n17285 = ~n17260 & n17284;
  assign n17286 = n17162 & ~n17285;
  assign n17287 = ~n17282 & ~n17286;
  assign n17288 = n17274 & n17278;
  assign n17289 = n17258 & ~n17288;
  assign n17290 = ~n17134 & ~n17161;
  assign n17291 = n17206 & n17262;
  assign n17292 = n17252 & ~n17291;
  assign n17293 = n17279 & n17292;
  assign n17294 = n17290 & ~n17293;
  assign n17295 = ~n17289 & ~n17294;
  assign n17296 = n17287 & n17295;
  assign n17297 = ~n17270 & n17296;
  assign n17298 = n17267 & n17297;
  assign n17299 = n17254 & n17298;
  assign n17300 = n17299 ^ n14601;
  assign n17301 = n17300 ^ x706;
  assign n17302 = n15597 ^ x640;
  assign n17303 = n16981 ^ x645;
  assign n17304 = ~n17302 & n17303;
  assign n17305 = n16293 & n16311;
  assign n17306 = n16227 & n16296;
  assign n17307 = ~n17305 & ~n17306;
  assign n17308 = ~n16287 & n17307;
  assign n17309 = ~n16301 & ~n16318;
  assign n17310 = n16293 & ~n17309;
  assign n17311 = ~n16296 & ~n16327;
  assign n17312 = ~n16345 & n17311;
  assign n17313 = n16298 & ~n17312;
  assign n17314 = ~n17310 & ~n17313;
  assign n17315 = n16227 & n16306;
  assign n17316 = ~n16308 & n16329;
  assign n17317 = n16288 & ~n17316;
  assign n17318 = n16298 & ~n16326;
  assign n17319 = ~n16291 & n17227;
  assign n17320 = ~n16311 & n17319;
  assign n17321 = n16227 & ~n17320;
  assign n17322 = ~n17318 & ~n17321;
  assign n17323 = ~n16325 & n17220;
  assign n17324 = n17323 ^ n16225;
  assign n17325 = n17324 ^ n17323;
  assign n17326 = ~n16285 & ~n16313;
  assign n17327 = n17326 ^ n17323;
  assign n17328 = ~n17325 & n17327;
  assign n17329 = n17328 ^ n17323;
  assign n17330 = n16226 & ~n17329;
  assign n17331 = n17322 & ~n17330;
  assign n17332 = n16305 & n17331;
  assign n17333 = ~n17317 & n17332;
  assign n17334 = ~n17315 & n17333;
  assign n17335 = n17314 & n17334;
  assign n17336 = n17214 & n17335;
  assign n17337 = n17308 & n17336;
  assign n17338 = n17337 ^ n14626;
  assign n17339 = n17338 ^ x643;
  assign n17340 = n15152 & n15176;
  assign n17341 = n14958 & n15147;
  assign n17342 = ~n17340 & ~n17341;
  assign n17343 = ~n15158 & ~n15190;
  assign n17344 = n15149 & ~n17343;
  assign n17345 = n14959 & ~n15181;
  assign n17346 = ~n17344 & ~n17345;
  assign n17347 = n17342 & n17346;
  assign n17348 = n15185 & ~n15193;
  assign n17349 = ~n15204 & n16205;
  assign n17350 = n15164 & ~n17349;
  assign n17351 = ~n15178 & ~n15203;
  assign n17352 = n15149 & ~n17351;
  assign n17353 = ~n15150 & n15180;
  assign n17354 = n15164 & ~n17353;
  assign n17355 = ~n17352 & ~n17354;
  assign n17356 = n15163 & ~n15193;
  assign n17357 = ~n15169 & n16551;
  assign n17358 = n15152 & ~n17357;
  assign n17359 = n15187 & ~n15204;
  assign n17360 = n14959 & ~n17359;
  assign n17361 = ~n17358 & ~n17360;
  assign n17362 = ~n17356 & n17361;
  assign n17363 = n17355 & n17362;
  assign n17364 = n15154 & n17363;
  assign n17365 = ~n17350 & n17364;
  assign n17366 = ~n17348 & n17365;
  assign n17367 = n17347 & n17366;
  assign n17368 = n16204 & n17367;
  assign n17369 = n17368 ^ n14660;
  assign n17370 = n17369 ^ x642;
  assign n17371 = n17339 & n17370;
  assign n17372 = n14782 ^ x641;
  assign n17373 = n17050 ^ x644;
  assign n17374 = ~n17372 & n17373;
  assign n17375 = n17371 & n17374;
  assign n17376 = n17304 & n17375;
  assign n17377 = ~n17302 & ~n17303;
  assign n17378 = ~n17339 & ~n17370;
  assign n17379 = n17372 & ~n17373;
  assign n17380 = n17378 & n17379;
  assign n17381 = n17377 & n17380;
  assign n17382 = ~n17376 & ~n17381;
  assign n17383 = n17302 & n17303;
  assign n17384 = n17339 & ~n17370;
  assign n17385 = n17379 & n17384;
  assign n17386 = n17383 & n17385;
  assign n17387 = ~n17339 & n17370;
  assign n17388 = n17374 & n17387;
  assign n17389 = ~n17372 & ~n17373;
  assign n17390 = n17378 & n17389;
  assign n17391 = ~n17388 & ~n17390;
  assign n17392 = n17304 & ~n17391;
  assign n17393 = ~n17386 & ~n17392;
  assign n17394 = n17302 & ~n17303;
  assign n17395 = n17379 & n17387;
  assign n17396 = ~n17385 & ~n17395;
  assign n17397 = n17394 & ~n17396;
  assign n17398 = n17372 & n17373;
  assign n17399 = n17371 & n17398;
  assign n17400 = n17394 & n17399;
  assign n17401 = n17383 & n17395;
  assign n17402 = ~n17400 & ~n17401;
  assign n17403 = n17371 & n17379;
  assign n17404 = n17377 & n17403;
  assign n17405 = n17304 & n17380;
  assign n17406 = n17383 & n17388;
  assign n17407 = n17387 & n17398;
  assign n17408 = ~n17304 & n17407;
  assign n17409 = n17374 & n17378;
  assign n17410 = n17374 & n17384;
  assign n17411 = n17371 & n17389;
  assign n17412 = ~n17375 & ~n17411;
  assign n17413 = ~n17410 & n17412;
  assign n17414 = ~n17409 & n17413;
  assign n17415 = n17394 & ~n17414;
  assign n17416 = ~n17408 & ~n17415;
  assign n17417 = ~n17395 & ~n17399;
  assign n17418 = n17384 & n17398;
  assign n17419 = ~n17403 & ~n17418;
  assign n17420 = n17417 & n17419;
  assign n17421 = n17304 & ~n17420;
  assign n17422 = ~n17377 & ~n17383;
  assign n17423 = n17378 & n17398;
  assign n17424 = n17384 & n17389;
  assign n17425 = ~n17410 & ~n17424;
  assign n17426 = ~n17411 & n17425;
  assign n17427 = ~n17377 & n17426;
  assign n17428 = n17387 & n17389;
  assign n17429 = ~n17410 & ~n17428;
  assign n17430 = n17412 & n17429;
  assign n17431 = ~n17383 & n17430;
  assign n17432 = ~n17427 & ~n17431;
  assign n17433 = ~n17423 & ~n17432;
  assign n17434 = ~n17422 & ~n17433;
  assign n17435 = ~n17421 & ~n17434;
  assign n17436 = n17416 & n17435;
  assign n17437 = ~n17406 & n17436;
  assign n17438 = ~n17405 & n17437;
  assign n17439 = ~n17404 & n17438;
  assign n17440 = n17402 & n17439;
  assign n17441 = ~n17397 & n17440;
  assign n17442 = n17393 & n17441;
  assign n17443 = n17382 & n17442;
  assign n17444 = n17443 ^ n14735;
  assign n17445 = n17444 ^ x711;
  assign n17446 = n17301 & ~n17445;
  assign n17447 = n17133 & n17446;
  assign n17448 = ~n17301 & n17445;
  assign n17449 = ~n16190 & n16903;
  assign n17450 = n16539 & n17449;
  assign n17451 = n16190 & ~n16903;
  assign n17452 = n17451 ^ n17124;
  assign n17453 = n17452 ^ n17451;
  assign n17454 = n17125 ^ n16903;
  assign n17455 = n16190 & ~n17454;
  assign n17456 = n17455 ^ n16903;
  assign n17457 = n17456 ^ n17451;
  assign n17458 = ~n17453 & ~n17457;
  assign n17459 = n17458 ^ n17451;
  assign n17460 = ~n16905 & ~n17459;
  assign n17461 = ~n17450 & n17460;
  assign n17462 = n17448 & ~n17461;
  assign n17463 = ~n17447 & ~n17462;
  assign n17464 = ~n17301 & ~n17445;
  assign n17465 = n16903 ^ n16190;
  assign n17466 = n17129 ^ n16539;
  assign n17467 = n17124 ^ n16903;
  assign n17468 = n17467 ^ n16539;
  assign n17469 = n17468 ^ n16539;
  assign n17470 = n17466 & n17469;
  assign n17471 = n17470 ^ n16539;
  assign n17472 = n17465 & ~n17471;
  assign n17473 = n17472 ^ n17467;
  assign n17474 = n17464 & ~n17473;
  assign n17475 = n17301 & n17445;
  assign n17476 = ~n16190 & n17124;
  assign n17477 = n17127 & n17476;
  assign n17479 = n16190 & n16539;
  assign n17478 = ~n16539 & n17449;
  assign n17480 = n17479 ^ n17478;
  assign n17481 = n17124 & n17480;
  assign n17482 = n17481 ^ n17479;
  assign n17483 = ~n17477 & ~n17482;
  assign n17484 = n16903 & n17479;
  assign n17485 = ~n17450 & ~n17451;
  assign n17486 = ~n16904 & n17485;
  assign n17487 = ~n17124 & ~n17486;
  assign n17488 = ~n17484 & ~n17487;
  assign n17489 = n17483 & n17488;
  assign n17490 = n17475 & ~n17489;
  assign n17491 = ~n17474 & ~n17490;
  assign n17492 = n17463 & n17491;
  assign n17493 = n17492 ^ n16625;
  assign n17494 = n17493 ^ x764;
  assign n17495 = n16223 ^ x659;
  assign n17496 = n16328 & n17220;
  assign n17497 = n16298 & ~n17496;
  assign n17498 = ~n16286 & n16326;
  assign n17499 = ~n16327 & n17498;
  assign n17500 = n16293 & ~n17499;
  assign n17501 = ~n17497 & ~n17500;
  assign n17502 = n16227 & ~n17228;
  assign n17503 = n16282 ^ n16257;
  assign n17504 = n17503 ^ n16281;
  assign n17505 = n17504 ^ n16257;
  assign n17506 = n17505 ^ n16281;
  assign n17507 = n17506 ^ n16283;
  assign n17508 = n16283 ^ n16257;
  assign n17509 = n17508 ^ n16257;
  assign n17510 = n16281 ^ n16257;
  assign n17511 = n17510 ^ n16257;
  assign n17512 = ~n17509 & n17511;
  assign n17513 = n17512 ^ n16257;
  assign n17514 = ~n17507 & ~n17513;
  assign n17515 = n17514 ^ n17504;
  assign n17516 = n16288 & ~n17515;
  assign n17517 = ~n17502 & ~n17516;
  assign n17518 = n17501 & n17517;
  assign n17519 = n16315 & n17518;
  assign n17520 = ~n16310 & n17519;
  assign n17521 = n17218 & n17520;
  assign n17522 = n17308 & n17521;
  assign n17523 = n17209 & n17522;
  assign n17524 = n16304 & n17523;
  assign n17525 = n17524 ^ n15357;
  assign n17526 = n17525 ^ x660;
  assign n17527 = n17495 & n17526;
  assign n17528 = n16660 & n16717;
  assign n17529 = n16723 & n16950;
  assign n17530 = ~n16753 & n17529;
  assign n17531 = ~n16659 & ~n17530;
  assign n17532 = ~n17528 & ~n17531;
  assign n17533 = n16739 & ~n16751;
  assign n17534 = n16957 & n17183;
  assign n17535 = n16707 & ~n17534;
  assign n17536 = ~n16713 & ~n16724;
  assign n17537 = ~n16722 & n17536;
  assign n17538 = n16719 & n17537;
  assign n17539 = ~n16776 & n17538;
  assign n17540 = n16721 & ~n17539;
  assign n17541 = ~n17535 & ~n17540;
  assign n17542 = ~n17533 & n17541;
  assign n17543 = n17532 & n17542;
  assign n17544 = n16716 & n17543;
  assign n17545 = n16948 & n17544;
  assign n17546 = ~n16729 & n17545;
  assign n17547 = n17546 ^ n15328;
  assign n17548 = n17547 ^ x661;
  assign n17549 = n16825 ^ x662;
  assign n17550 = n17548 & ~n17549;
  assign n17551 = n17527 & n17550;
  assign n17552 = ~n17495 & n17526;
  assign n17553 = ~n17548 & ~n17549;
  assign n17554 = n17552 & n17553;
  assign n17555 = ~n17551 & ~n17554;
  assign n17556 = n16386 ^ x658;
  assign n17557 = n16654 ^ x663;
  assign n17558 = n17556 & ~n17557;
  assign n17559 = n17526 ^ n17495;
  assign n17560 = n17559 ^ n17549;
  assign n17561 = n17549 ^ n17548;
  assign n17562 = n17548 ^ n17526;
  assign n17563 = n17562 ^ n17548;
  assign n17564 = ~n17561 & n17563;
  assign n17565 = n17564 ^ n17548;
  assign n17566 = ~n17560 & ~n17565;
  assign n17567 = n17566 ^ n17549;
  assign n17568 = n17558 & n17567;
  assign n17569 = n17556 & n17557;
  assign n17570 = n17527 & n17548;
  assign n17571 = n17495 & ~n17526;
  assign n17572 = ~n17548 & n17571;
  assign n17573 = n17549 & n17572;
  assign n17574 = ~n17570 & ~n17573;
  assign n17575 = n17548 & n17549;
  assign n17576 = ~n17495 & n17575;
  assign n17577 = ~n17495 & ~n17526;
  assign n17578 = n17550 & n17577;
  assign n17579 = n17527 & n17553;
  assign n17580 = ~n17578 & ~n17579;
  assign n17581 = ~n17576 & n17580;
  assign n17582 = n17574 & n17581;
  assign n17583 = ~n17554 & n17582;
  assign n17584 = n17569 & ~n17583;
  assign n17585 = ~n17568 & ~n17584;
  assign n17586 = ~n17552 & ~n17572;
  assign n17587 = n17549 & ~n17586;
  assign n17588 = n17550 & n17571;
  assign n17589 = n17527 & n17549;
  assign n17590 = ~n17548 & n17589;
  assign n17591 = ~n17588 & ~n17590;
  assign n17592 = ~n17587 & n17591;
  assign n17593 = ~n17578 & n17592;
  assign n17594 = n17593 ^ n17557;
  assign n17595 = n17594 ^ n17593;
  assign n17596 = n17527 & n17575;
  assign n17597 = n17553 & n17577;
  assign n17598 = ~n17596 & ~n17597;
  assign n17599 = n17581 & n17598;
  assign n17600 = ~n17587 & n17599;
  assign n17601 = n17600 ^ n17593;
  assign n17602 = n17595 & ~n17601;
  assign n17603 = n17602 ^ n17593;
  assign n17604 = ~n17556 & ~n17603;
  assign n17605 = n17585 & ~n17604;
  assign n17606 = n17555 & n17605;
  assign n17607 = n17606 ^ n16015;
  assign n17608 = n17607 ^ x689;
  assign n17609 = n17062 & n17081;
  assign n17610 = ~n17079 & ~n17609;
  assign n17611 = ~n17064 & ~n17103;
  assign n17612 = ~n17070 & n17611;
  assign n17613 = n17052 & ~n17612;
  assign n17614 = n17057 & n17103;
  assign n17615 = ~n17613 & ~n17614;
  assign n17616 = n17062 & ~n17102;
  assign n17617 = ~n17077 & ~n17092;
  assign n17618 = ~n17093 & n17617;
  assign n17619 = n17065 & ~n17618;
  assign n17620 = n17052 & n17096;
  assign n17621 = n17065 & n17072;
  assign n17622 = ~n17620 & ~n17621;
  assign n17623 = ~n17072 & ~n17095;
  assign n17624 = ~n17061 & n17623;
  assign n17625 = n17052 & ~n17624;
  assign n17626 = n17094 & n17611;
  assign n17627 = n17062 & ~n17626;
  assign n17628 = ~n17625 & ~n17627;
  assign n17629 = n17098 ^ n17051;
  assign n17630 = n17629 ^ n17098;
  assign n17631 = n17086 & ~n17093;
  assign n17632 = n17631 ^ n17098;
  assign n17633 = n17630 & n17632;
  assign n17634 = n17633 ^ n17098;
  assign n17635 = ~n17015 & ~n17634;
  assign n17636 = n17628 & ~n17635;
  assign n17637 = n17622 & n17636;
  assign n17638 = ~n17619 & n17637;
  assign n17639 = ~n17616 & n17638;
  assign n17640 = n17615 & n17639;
  assign n17641 = n17610 & n17640;
  assign n17642 = n17068 & n17641;
  assign n17643 = n17642 ^ n16000;
  assign n17644 = n17643 ^ x690;
  assign n17645 = n17608 & n17644;
  assign n17646 = n16625 ^ x670;
  assign n17647 = n17241 ^ x675;
  assign n17648 = ~n17646 & ~n17647;
  assign n17649 = ~n15544 & n16912;
  assign n17650 = n15289 & ~n17649;
  assign n17651 = n15546 & n16915;
  assign n17652 = ~n15531 & n17651;
  assign n17653 = n16368 & n17652;
  assign n17654 = n15566 & ~n17653;
  assign n17655 = ~n17650 & ~n17654;
  assign n17656 = n15549 & n16916;
  assign n17657 = ~n15539 & n17656;
  assign n17658 = n15552 & ~n17657;
  assign n17659 = ~n15577 & n16915;
  assign n17660 = ~n15544 & n17659;
  assign n17661 = ~n15526 & n17660;
  assign n17662 = n15529 & ~n17661;
  assign n17663 = ~n17658 & ~n17662;
  assign n17664 = n17655 & n17663;
  assign n17665 = ~n16940 & n17664;
  assign n17666 = n15535 & n17665;
  assign n17667 = n15543 & n17666;
  assign n17668 = n16366 & n17667;
  assign n17669 = n17668 ^ n14847;
  assign n17670 = n17669 ^ x672;
  assign n17671 = n17160 ^ x674;
  assign n17672 = n17670 & ~n17671;
  assign n17673 = n16785 ^ x671;
  assign n17674 = n15971 & ~n16075;
  assign n17675 = ~n16079 & ~n16098;
  assign n17676 = n16053 & ~n17675;
  assign n17677 = ~n16053 & ~n16085;
  assign n17678 = ~n15971 & ~n16080;
  assign n17679 = ~n16084 & n17678;
  assign n17680 = ~n17677 & ~n17679;
  assign n17681 = n16094 & ~n17680;
  assign n17682 = ~n16078 & ~n17681;
  assign n17683 = ~n17676 & ~n17682;
  assign n17684 = ~n17674 & n17683;
  assign n17685 = ~n16083 & n16100;
  assign n17686 = ~n16041 & n17685;
  assign n17687 = n17686 ^ n15970;
  assign n17688 = n17687 ^ n17686;
  assign n17689 = n17686 ^ n16630;
  assign n17690 = ~n17688 & n17689;
  assign n17691 = n17690 ^ n17686;
  assign n17692 = n16633 & ~n17691;
  assign n17693 = n17684 & ~n17692;
  assign n17694 = n16067 & n17693;
  assign n17695 = n16446 & n17694;
  assign n17696 = n16058 & n17695;
  assign n17697 = n17696 ^ n14876;
  assign n17698 = n17697 ^ x673;
  assign n17699 = ~n17673 & ~n17698;
  assign n17700 = n17672 & n17699;
  assign n17701 = n17648 & n17700;
  assign n17702 = ~n17646 & n17647;
  assign n17703 = ~n17673 & n17698;
  assign n17704 = ~n17670 & ~n17671;
  assign n17705 = n17703 & n17704;
  assign n17706 = ~n17670 & n17671;
  assign n17707 = n17699 & n17706;
  assign n17708 = ~n17705 & ~n17707;
  assign n17709 = n17702 & ~n17708;
  assign n17710 = ~n17701 & ~n17709;
  assign n17711 = n17699 & n17704;
  assign n17712 = n17702 & n17711;
  assign n17713 = n17646 & n17647;
  assign n17714 = n17672 & n17673;
  assign n17715 = n17673 & ~n17698;
  assign n17716 = n17706 & n17715;
  assign n17717 = ~n17714 & ~n17716;
  assign n17718 = n17713 & ~n17717;
  assign n17719 = ~n17712 & ~n17718;
  assign n17720 = n17647 ^ n17646;
  assign n17721 = n17670 & n17671;
  assign n17722 = n17699 & n17721;
  assign n17723 = n17720 & n17722;
  assign n17724 = n17704 & n17715;
  assign n17725 = n17646 & n17724;
  assign n17726 = ~n17723 & ~n17725;
  assign n17727 = n17646 & ~n17647;
  assign n17728 = n17672 & n17703;
  assign n17729 = ~n17707 & ~n17728;
  assign n17730 = n17727 & ~n17729;
  assign n17731 = n17671 ^ n17670;
  assign n17732 = n17673 & n17698;
  assign n17733 = ~n17731 & n17732;
  assign n17734 = n17703 & n17706;
  assign n17735 = n17703 & n17721;
  assign n17736 = n17672 & n17715;
  assign n17737 = ~n17716 & ~n17736;
  assign n17738 = ~n17735 & n17737;
  assign n17739 = ~n17734 & n17738;
  assign n17740 = ~n17733 & n17739;
  assign n17741 = ~n17724 & n17740;
  assign n17742 = n17648 & ~n17741;
  assign n17743 = n17698 ^ n17670;
  assign n17744 = n17743 ^ n17698;
  assign n17745 = n17698 ^ n17671;
  assign n17746 = n17745 ^ n17698;
  assign n17747 = n17744 & ~n17746;
  assign n17748 = n17747 ^ n17698;
  assign n17749 = ~n17673 & n17748;
  assign n17750 = n17713 & n17749;
  assign n17751 = n17706 & n17732;
  assign n17752 = n17704 & n17732;
  assign n17753 = n17672 & n17732;
  assign n17754 = n17715 & n17721;
  assign n17755 = ~n17753 & ~n17754;
  assign n17756 = ~n17752 & n17755;
  assign n17757 = ~n17751 & n17756;
  assign n17758 = n17727 & ~n17757;
  assign n17759 = ~n17670 & n17732;
  assign n17760 = ~n17672 & ~n17721;
  assign n17761 = n17715 & ~n17760;
  assign n17762 = ~n17759 & ~n17761;
  assign n17763 = n17702 & ~n17762;
  assign n17764 = ~n17758 & ~n17763;
  assign n17765 = ~n17750 & n17764;
  assign n17766 = ~n17742 & n17765;
  assign n17767 = ~n17730 & n17766;
  assign n17768 = n17726 & n17767;
  assign n17769 = n17719 & n17768;
  assign n17770 = n17710 & n17769;
  assign n17771 = n17770 ^ n14957;
  assign n17772 = n17771 ^ x692;
  assign n17773 = n16839 & ~n16879;
  assign n17774 = n16851 & n16873;
  assign n17775 = n16827 & ~n16870;
  assign n17776 = ~n17774 & ~n17775;
  assign n17777 = ~n17773 & n17776;
  assign n17778 = n16839 & n16873;
  assign n17779 = n16836 & n16851;
  assign n17780 = ~n17778 & ~n17779;
  assign n17781 = n16839 & n16846;
  assign n17782 = ~n16657 & n16855;
  assign n17783 = ~n16886 & n17782;
  assign n17784 = n16829 & ~n17783;
  assign n17785 = ~n16839 & ~n16851;
  assign n17786 = n16859 & ~n17785;
  assign n17787 = ~n16886 & ~n16888;
  assign n17788 = ~n16852 & n17787;
  assign n17789 = n16839 & ~n17788;
  assign n17790 = ~n16848 & ~n16875;
  assign n17791 = ~n16869 & n17790;
  assign n17792 = ~n16836 & n17791;
  assign n17793 = n16829 & ~n17792;
  assign n17794 = ~n16859 & ~n16873;
  assign n17795 = ~n16831 & n17794;
  assign n17796 = n16827 & ~n17795;
  assign n17797 = ~n17793 & ~n17796;
  assign n17798 = ~n17789 & n17797;
  assign n17799 = ~n17786 & n17798;
  assign n17800 = n16827 & ~n16868;
  assign n17801 = n16592 & n16838;
  assign n17802 = n16855 & ~n17801;
  assign n17803 = ~n16867 & n17802;
  assign n17804 = ~n16875 & n17803;
  assign n17805 = n16851 & ~n17804;
  assign n17806 = ~n17800 & ~n17805;
  assign n17807 = n17799 & n17806;
  assign n17808 = ~n17784 & n17807;
  assign n17809 = ~n17781 & n17808;
  assign n17810 = n17780 & n17809;
  assign n17811 = n17777 & n17810;
  assign n17812 = n17811 ^ n16038;
  assign n17813 = n17812 ^ x691;
  assign n17814 = ~n17772 & n17813;
  assign n17815 = n17645 & n17814;
  assign n17816 = ~n17283 & ~n17291;
  assign n17817 = ~n17276 & n17816;
  assign n17818 = n17162 & ~n17817;
  assign n17819 = n17244 & n17255;
  assign n17820 = ~n17251 & ~n17819;
  assign n17821 = n17271 & ~n17820;
  assign n17822 = ~n17273 & ~n17275;
  assign n17823 = n17258 & ~n17822;
  assign n17824 = ~n17821 & ~n17823;
  assign n17825 = ~n17276 & n17820;
  assign n17826 = n17258 & ~n17825;
  assign n17827 = ~n17261 & n17274;
  assign n17828 = n17162 & ~n17827;
  assign n17829 = ~n17826 & ~n17828;
  assign n17830 = n17281 & n17290;
  assign n17831 = n17279 & n17816;
  assign n17832 = n17271 & ~n17831;
  assign n17833 = ~n17830 & ~n17832;
  assign n17834 = n17829 & n17833;
  assign n17835 = ~n17246 & n17834;
  assign n17836 = n17824 & n17835;
  assign n17837 = n17267 & n17836;
  assign n17838 = ~n17818 & n17837;
  assign n17839 = n17838 ^ n15969;
  assign n17840 = n17839 ^ x688;
  assign n17841 = n16129 & n16133;
  assign n17842 = ~n16124 & ~n16132;
  assign n17843 = n16127 & ~n17842;
  assign n17844 = ~n17841 & ~n17843;
  assign n17845 = n15219 & n16164;
  assign n17846 = ~n16134 & n16154;
  assign n17847 = ~n17845 & ~n17846;
  assign n17848 = ~n16154 & ~n16161;
  assign n17849 = ~n16155 & n17848;
  assign n17850 = n16121 & ~n17849;
  assign n17851 = n16127 & ~n16179;
  assign n17852 = n16121 & n16142;
  assign n17853 = ~n16120 & ~n17852;
  assign n17854 = ~n16148 & ~n16160;
  assign n17855 = n15220 & ~n17854;
  assign n17856 = n16156 & n16182;
  assign n17857 = n16127 & ~n17856;
  assign n17858 = ~n17855 & ~n17857;
  assign n17859 = ~n16141 & ~n16178;
  assign n17860 = ~n16124 & n17859;
  assign n17861 = n16121 & ~n17860;
  assign n17862 = n16119 & ~n16124;
  assign n17863 = ~n16141 & n17862;
  assign n17864 = n17863 ^ n17859;
  assign n17865 = n17859 ^ n15219;
  assign n17866 = n17865 ^ n17859;
  assign n17867 = n17864 & n17866;
  assign n17868 = n17867 ^ n17859;
  assign n17869 = ~n16177 & ~n17868;
  assign n17870 = ~n17861 & ~n17869;
  assign n17871 = n17858 & n17870;
  assign n17872 = n17853 & n17871;
  assign n17873 = ~n17851 & n17872;
  assign n17874 = ~n17850 & n17873;
  assign n17875 = n17847 & n17874;
  assign n17876 = n17844 & n17875;
  assign n17877 = n16150 & n17876;
  assign n17878 = n17877 ^ n15094;
  assign n17879 = n17878 ^ x693;
  assign n17880 = n17840 & ~n17879;
  assign n17881 = n17815 & n17880;
  assign n17882 = ~n17840 & n17879;
  assign n17883 = n17815 & n17882;
  assign n17884 = n17840 & n17879;
  assign n17885 = ~n17608 & n17644;
  assign n17886 = ~n17772 & ~n17813;
  assign n17887 = n17885 & n17886;
  assign n17888 = n17884 & n17887;
  assign n17889 = ~n17883 & ~n17888;
  assign n17890 = n17772 & n17813;
  assign n17891 = n17885 & n17890;
  assign n17892 = ~n17608 & ~n17644;
  assign n17893 = n17886 & n17892;
  assign n17894 = ~n17891 & ~n17893;
  assign n17895 = n17884 & ~n17894;
  assign n17896 = n17889 & ~n17895;
  assign n17897 = n17645 & n17886;
  assign n17898 = n17608 & ~n17644;
  assign n17899 = n17772 & ~n17813;
  assign n17900 = n17898 & n17899;
  assign n17901 = ~n17897 & ~n17900;
  assign n17902 = n17882 & ~n17901;
  assign n17903 = n17645 & n17899;
  assign n17904 = n17880 & n17903;
  assign n17905 = ~n17840 & ~n17879;
  assign n17906 = n17892 & n17899;
  assign n17907 = n17905 & n17906;
  assign n17908 = ~n17904 & ~n17907;
  assign n17909 = n17814 & n17885;
  assign n17910 = n17905 & n17909;
  assign n17911 = n17884 & n17906;
  assign n17912 = ~n17910 & ~n17911;
  assign n17913 = n17814 & n17898;
  assign n17914 = n17905 & n17913;
  assign n17915 = n17814 & n17892;
  assign n17916 = ~n17891 & ~n17915;
  assign n17917 = n17885 & n17899;
  assign n17918 = ~n17913 & ~n17917;
  assign n17919 = n17916 & n17918;
  assign n17920 = ~n17903 & n17919;
  assign n17921 = n17882 & ~n17920;
  assign n17922 = n17890 & n17892;
  assign n17923 = n17645 & n17890;
  assign n17924 = n17886 & n17898;
  assign n17925 = ~n17923 & ~n17924;
  assign n17926 = ~n17922 & n17925;
  assign n17927 = ~n17906 & n17926;
  assign n17928 = n17880 & ~n17927;
  assign n17929 = n17890 & n17898;
  assign n17930 = ~n17897 & ~n17929;
  assign n17931 = ~n17923 & n17930;
  assign n17932 = n17905 & ~n17931;
  assign n17935 = ~n17887 & ~n17917;
  assign n17933 = n17925 & ~n17929;
  assign n17934 = ~n17815 & n17933;
  assign n17936 = n17935 ^ n17934;
  assign n17937 = n17936 ^ n17935;
  assign n17938 = n17935 ^ n17840;
  assign n17939 = n17938 ^ n17935;
  assign n17940 = ~n17937 & n17939;
  assign n17941 = n17940 ^ n17935;
  assign n17942 = n17879 & ~n17941;
  assign n17943 = n17942 ^ n17935;
  assign n17944 = ~n17932 & n17943;
  assign n17945 = ~n17928 & n17944;
  assign n17946 = ~n17921 & n17945;
  assign n17947 = ~n17914 & n17946;
  assign n17948 = n17912 & n17947;
  assign n17949 = n17908 & n17948;
  assign n17950 = ~n17902 & n17949;
  assign n17951 = n17896 & n17950;
  assign n17952 = ~n17881 & n17951;
  assign n17953 = n17952 ^ n16654;
  assign n17954 = n17953 ^ x761;
  assign n17955 = n17494 & n17954;
  assign n17956 = n16657 & n16839;
  assign n17957 = n16827 & n16836;
  assign n17958 = n16829 & ~n16876;
  assign n17959 = ~n17957 & ~n17958;
  assign n17960 = ~n17956 & n17959;
  assign n17961 = n16855 & n16879;
  assign n17962 = n16827 & ~n17961;
  assign n17963 = n16849 & n16860;
  assign n17964 = n17787 & n17963;
  assign n17965 = n16851 & ~n17964;
  assign n17966 = ~n16854 & ~n16886;
  assign n17967 = ~n16838 & n17966;
  assign n17968 = ~n16867 & n17967;
  assign n17969 = ~n16869 & n17968;
  assign n17970 = n16839 & ~n17969;
  assign n17971 = ~n17965 & ~n17970;
  assign n17972 = ~n17962 & n17971;
  assign n17973 = ~n16569 & n16829;
  assign n17974 = n16655 ^ n16592;
  assign n17975 = n17974 ^ n16829;
  assign n17976 = n17973 ^ n16656;
  assign n17977 = n17975 & n17976;
  assign n17978 = n17977 ^ n16656;
  assign n17979 = n17973 & n17978;
  assign n17980 = n17972 & ~n17979;
  assign n17981 = n17780 & n17980;
  assign n17982 = n17960 & n17981;
  assign n17983 = n17776 & n17982;
  assign n17984 = n16834 & n17983;
  assign n17985 = n17984 ^ n15048;
  assign n17986 = n17985 ^ x698;
  assign n17987 = n17878 ^ x695;
  assign n17988 = n17986 & ~n17987;
  assign n17989 = n17271 & n17276;
  assign n17990 = n17247 & n17262;
  assign n17991 = ~n17260 & ~n17990;
  assign n17992 = n17258 & ~n17991;
  assign n17993 = ~n17989 & ~n17992;
  assign n17994 = n17245 & n17271;
  assign n17995 = ~n17256 & ~n17273;
  assign n17996 = n17290 & ~n17995;
  assign n17997 = ~n17994 & ~n17996;
  assign n17998 = n17264 & ~n17272;
  assign n17999 = ~n17819 & n17998;
  assign n18000 = n17162 & ~n17999;
  assign n18001 = ~n17242 & n17247;
  assign n18002 = n17271 & n18001;
  assign n18003 = ~n17248 & ~n17256;
  assign n18004 = n17258 & ~n18003;
  assign n18005 = ~n17260 & ~n17263;
  assign n18006 = n17271 & ~n18005;
  assign n18007 = ~n18004 & ~n18006;
  assign n18008 = ~n17261 & ~n17275;
  assign n18009 = ~n17990 & n18008;
  assign n18010 = n17816 & n18009;
  assign n18011 = n18010 ^ n17276;
  assign n18012 = n18011 ^ n17276;
  assign n18013 = n17276 ^ n17161;
  assign n18014 = n18013 ^ n17276;
  assign n18015 = ~n18012 & ~n18014;
  assign n18016 = n18015 ^ n17276;
  assign n18017 = ~n17134 & n18016;
  assign n18018 = n18017 ^ n17276;
  assign n18019 = n18007 & ~n18018;
  assign n18020 = ~n18002 & n18019;
  assign n18021 = ~n18000 & n18020;
  assign n18022 = n17997 & n18021;
  assign n18023 = ~n17270 & n18022;
  assign n18024 = n17824 & n18023;
  assign n18025 = n17993 & n18024;
  assign n18026 = n17254 & n18025;
  assign n18027 = n18026 ^ n15140;
  assign n18028 = n18027 ^ x697;
  assign n18029 = ~n16483 & ~n16488;
  assign n18030 = n16478 & ~n18029;
  assign n18031 = n16482 & n16499;
  assign n18032 = ~n16514 & ~n18031;
  assign n18033 = n18032 ^ n16478;
  assign n18034 = n18033 ^ n18032;
  assign n18035 = n18032 ^ n16501;
  assign n18036 = n18035 ^ n18032;
  assign n18037 = ~n18034 & n18036;
  assign n18038 = n18037 ^ n18032;
  assign n18039 = ~n16477 & ~n18038;
  assign n18040 = n18039 ^ n18032;
  assign n18041 = ~n18030 & n18040;
  assign n18042 = n16361 & n16506;
  assign n18043 = ~n16489 & ~n16510;
  assign n18044 = ~n16479 & ~n18043;
  assign n18045 = ~n18042 & ~n18044;
  assign n18046 = ~n16475 & ~n16506;
  assign n18047 = ~n16519 & n18046;
  assign n18048 = ~n16491 & n18047;
  assign n18049 = n16477 & ~n18048;
  assign n18050 = n16427 & n16499;
  assign n18051 = n16521 & ~n18050;
  assign n18052 = n16478 & ~n18051;
  assign n18053 = ~n16475 & n16492;
  assign n18054 = ~n16505 & n18053;
  assign n18055 = ~n16476 & n16493;
  assign n18056 = ~n16481 & n18055;
  assign n18057 = ~n18054 & ~n18056;
  assign n18058 = n18032 & ~n18057;
  assign n18059 = n16479 & ~n18058;
  assign n18060 = ~n18052 & ~n18059;
  assign n18061 = ~n18049 & n18060;
  assign n18062 = n18045 & n18061;
  assign n18063 = n16360 ^ n16224;
  assign n18064 = n16512 ^ n16360;
  assign n18065 = n18064 ^ n16512;
  assign n18066 = n16512 ^ n16481;
  assign n18067 = ~n18065 & n18066;
  assign n18068 = n18067 ^ n16512;
  assign n18069 = ~n18063 & n18068;
  assign n18070 = n18062 & ~n18069;
  assign n18071 = n18041 & n18070;
  assign n18072 = n18071 ^ n14996;
  assign n18073 = n18072 ^ x696;
  assign n18074 = ~n18028 & n18073;
  assign n18075 = n17988 & n18074;
  assign n18076 = n17771 ^ x694;
  assign n18077 = n17383 & ~n17412;
  assign n18078 = n17303 ^ n17302;
  assign n18079 = n17407 ^ n17303;
  assign n18080 = n18079 ^ n17407;
  assign n18081 = n17409 ^ n17407;
  assign n18082 = ~n18080 & n18081;
  assign n18083 = n18082 ^ n17407;
  assign n18084 = n18078 & n18083;
  assign n18085 = ~n18077 & ~n18084;
  assign n18086 = ~n17422 & ~n17429;
  assign n18087 = n17391 & ~n17418;
  assign n18088 = n17417 & n18087;
  assign n18089 = ~n17411 & n18088;
  assign n18090 = n17394 & ~n18089;
  assign n18091 = ~n18086 & ~n18090;
  assign n18092 = ~n17380 & ~n17407;
  assign n18093 = n17383 & ~n18092;
  assign n18094 = ~n17423 & n17425;
  assign n18095 = n17304 & ~n18094;
  assign n18096 = ~n17385 & n17417;
  assign n18097 = ~n17409 & n18096;
  assign n18098 = n17377 & ~n18097;
  assign n18099 = ~n18095 & ~n18098;
  assign n18100 = ~n18093 & n18099;
  assign n18101 = n18091 & n18100;
  assign n18102 = n17382 & n18101;
  assign n18103 = n18085 & n18102;
  assign n18104 = n17393 & n18103;
  assign n18105 = ~n17403 & n18104;
  assign n18106 = n18105 ^ n14817;
  assign n18107 = n18106 ^ x699;
  assign n18108 = ~n18076 & n18107;
  assign n18109 = n18075 & n18108;
  assign n18110 = n18076 & ~n18107;
  assign n18111 = n18028 & n18073;
  assign n18112 = n17988 & n18111;
  assign n18113 = ~n17986 & ~n17987;
  assign n18114 = n18028 & ~n18073;
  assign n18115 = n18113 & n18114;
  assign n18116 = ~n18112 & ~n18115;
  assign n18117 = n18110 & ~n18116;
  assign n18118 = ~n18109 & ~n18117;
  assign n18119 = ~n18076 & ~n18107;
  assign n18120 = n18075 & n18119;
  assign n18121 = n17986 & n17987;
  assign n18122 = n18114 & n18121;
  assign n18123 = n18076 & n18107;
  assign n18124 = n18122 & n18123;
  assign n18125 = ~n17986 & n17987;
  assign n18126 = n18111 & n18125;
  assign n18127 = n18108 & n18126;
  assign n18128 = ~n18124 & ~n18127;
  assign n18129 = ~n18120 & n18128;
  assign n18130 = ~n18028 & ~n18073;
  assign n18131 = n17988 & n18130;
  assign n18132 = n18123 & n18131;
  assign n18133 = n18108 & n18122;
  assign n18134 = n18074 & n18121;
  assign n18135 = n18114 & n18125;
  assign n18136 = ~n18134 & ~n18135;
  assign n18137 = n18119 & ~n18136;
  assign n18138 = ~n18133 & ~n18137;
  assign n18139 = ~n18132 & n18138;
  assign n18140 = n18119 & n18122;
  assign n18141 = n18111 & n18121;
  assign n18142 = n18108 & n18141;
  assign n18143 = n18110 & n18134;
  assign n18144 = ~n18142 & ~n18143;
  assign n18145 = ~n18140 & n18144;
  assign n18146 = n17988 & n18114;
  assign n18147 = n18074 & n18125;
  assign n18148 = n18121 & n18130;
  assign n18149 = ~n18147 & ~n18148;
  assign n18150 = ~n18146 & n18149;
  assign n18151 = n18110 & ~n18150;
  assign n18152 = n18113 & n18130;
  assign n18153 = ~n18131 & ~n18152;
  assign n18154 = ~n18147 & n18153;
  assign n18155 = ~n18115 & n18154;
  assign n18156 = n18108 & ~n18155;
  assign n18157 = ~n18151 & ~n18156;
  assign n18158 = ~n18075 & n18149;
  assign n18159 = ~n18152 & n18158;
  assign n18160 = n18123 & ~n18159;
  assign n18166 = n18111 & n18113;
  assign n18167 = ~n18126 & ~n18166;
  assign n18161 = n18125 & n18130;
  assign n18162 = n18074 & n18113;
  assign n18163 = ~n18146 & ~n18162;
  assign n18164 = ~n18152 & n18163;
  assign n18165 = ~n18161 & n18164;
  assign n18168 = n18167 ^ n18165;
  assign n18169 = n18168 ^ n18167;
  assign n18170 = n18167 ^ n18107;
  assign n18171 = n18170 ^ n18167;
  assign n18172 = ~n18169 & ~n18171;
  assign n18173 = n18172 ^ n18167;
  assign n18174 = ~n18076 & ~n18173;
  assign n18175 = n18174 ^ n18167;
  assign n18176 = ~n18160 & n18175;
  assign n18177 = n18157 & n18176;
  assign n18178 = n18145 & n18177;
  assign n18179 = n18139 & n18178;
  assign n18180 = n18129 & n18179;
  assign n18181 = n18118 & n18180;
  assign n18182 = n18181 ^ n16568;
  assign n18183 = n18182 ^ x762;
  assign n18184 = ~n17561 & n17571;
  assign n18185 = ~n17554 & ~n18184;
  assign n18186 = n17577 ^ n17527;
  assign n18187 = ~n17548 & n18186;
  assign n18188 = n18187 ^ n17527;
  assign n18189 = n17549 & n18188;
  assign n18190 = n17548 & n17552;
  assign n18191 = ~n17579 & ~n18190;
  assign n18192 = ~n18189 & n18191;
  assign n18193 = n18185 & n18192;
  assign n18194 = n17558 & n18193;
  assign n18195 = n18188 ^ n17552;
  assign n18196 = ~n17549 & n18195;
  assign n18197 = n18196 ^ n17552;
  assign n18198 = n18185 & ~n18197;
  assign n18199 = ~n17578 & n18198;
  assign n18200 = n17569 & ~n18199;
  assign n18201 = ~n18194 & ~n18200;
  assign n18202 = ~n17556 & n17557;
  assign n18203 = ~n18189 & ~n18190;
  assign n18204 = n17591 & n18203;
  assign n18205 = n17580 & n18204;
  assign n18206 = n18202 & ~n18205;
  assign n18207 = ~n17556 & ~n17557;
  assign n18208 = n17571 ^ n17495;
  assign n18209 = ~n17575 & ~n18208;
  assign n18210 = n18209 ^ n17495;
  assign n18211 = n18191 & n18210;
  assign n18212 = ~n17554 & n18211;
  assign n18213 = n18207 & ~n18212;
  assign n18214 = ~n18206 & ~n18213;
  assign n18215 = n18201 & n18214;
  assign n18216 = n18215 ^ n15759;
  assign n18217 = n18216 ^ x718;
  assign n18218 = n16848 & ~n17785;
  assign n18219 = ~n16861 & ~n17787;
  assign n18220 = ~n18218 & ~n18219;
  assign n18221 = ~n16840 & n16875;
  assign n18222 = n16879 & n17967;
  assign n18223 = n18222 ^ n17794;
  assign n18224 = n18223 ^ n17794;
  assign n18225 = n17794 ^ n16786;
  assign n18226 = n18225 ^ n17794;
  assign n18227 = ~n18224 & ~n18226;
  assign n18228 = n18227 ^ n17794;
  assign n18229 = n16826 & ~n18228;
  assign n18230 = n18229 ^ n17794;
  assign n18231 = ~n18221 & n18230;
  assign n18232 = n18220 & n18231;
  assign n18233 = n17960 & n18232;
  assign n18234 = n16843 & n18233;
  assign n18235 = n17777 & n18234;
  assign n18236 = n16834 & n18235;
  assign n18237 = n18236 ^ n15443;
  assign n18238 = n18237 ^ x723;
  assign n18239 = ~n18217 & ~n18238;
  assign n18240 = ~n16116 & ~n16148;
  assign n18241 = n16127 & ~n18240;
  assign n18242 = n16133 & ~n17842;
  assign n18243 = ~n18241 & ~n18242;
  assign n18244 = ~n16134 & n16142;
  assign n18245 = ~n16132 & n16182;
  assign n18246 = ~n16155 & n18245;
  assign n18247 = ~n16161 & n18246;
  assign n18248 = n16121 & ~n18247;
  assign n18249 = ~n18244 & ~n18248;
  assign n18250 = n15220 & n16141;
  assign n18251 = ~n16116 & ~n16129;
  assign n18252 = n16133 & ~n18251;
  assign n18253 = ~n16161 & n17859;
  assign n18254 = n16127 & ~n18253;
  assign n18255 = ~n16139 & ~n16155;
  assign n18256 = ~n15220 & n18255;
  assign n18257 = ~n16154 & n16163;
  assign n18258 = ~n18256 & ~n18257;
  assign n18259 = ~n16164 & ~n18258;
  assign n18260 = ~n16134 & ~n18259;
  assign n18261 = ~n18254 & ~n18260;
  assign n18262 = ~n18252 & n18261;
  assign n18263 = ~n18250 & n18262;
  assign n18264 = n18249 & n18263;
  assign n18265 = n18243 & n18264;
  assign n18266 = ~n16187 & n18265;
  assign n18267 = n17853 & n18266;
  assign n18268 = n18267 ^ n15837;
  assign n18269 = n18268 ^ x719;
  assign n18270 = n16478 & ~n16492;
  assign n18271 = ~n18069 & ~n18270;
  assign n18272 = n16477 & ~n16520;
  assign n18273 = ~n16506 & ~n18050;
  assign n18274 = n16479 & ~n18273;
  assign n18275 = n16478 & ~n18046;
  assign n18276 = ~n16481 & n16527;
  assign n18277 = n16477 & ~n18276;
  assign n18278 = ~n18275 & ~n18277;
  assign n18279 = n16484 & n18043;
  assign n18280 = n16505 & ~n18279;
  assign n18281 = ~n16491 & n18029;
  assign n18282 = n16361 & ~n18281;
  assign n18283 = ~n18280 & ~n18282;
  assign n18284 = n18278 & n18283;
  assign n18285 = ~n18274 & n18284;
  assign n18286 = ~n18272 & n18285;
  assign n18287 = ~n16513 & n18286;
  assign n18288 = n16490 ^ n16360;
  assign n18289 = n18288 ^ n16490;
  assign n18290 = n16520 ^ n16490;
  assign n18291 = ~n18289 & ~n18290;
  assign n18292 = n18291 ^ n16490;
  assign n18293 = n18063 & n18292;
  assign n18294 = n18287 & ~n18293;
  assign n18295 = n18271 & n18294;
  assign n18296 = n18041 & n18295;
  assign n18297 = n18296 ^ n15249;
  assign n18298 = n18297 ^ x722;
  assign n18299 = n17258 & n17283;
  assign n18300 = n17292 & n18008;
  assign n18301 = ~n17269 & n18300;
  assign n18302 = n17271 & ~n18301;
  assign n18303 = ~n18299 & ~n18302;
  assign n18304 = ~n17269 & ~n18001;
  assign n18305 = n17991 & n18304;
  assign n18306 = ~n17263 & n18305;
  assign n18307 = n17290 & ~n18306;
  assign n18308 = n17278 & ~n17819;
  assign n18309 = n18308 ^ n18304;
  assign n18310 = n18308 ^ n17161;
  assign n18311 = n17268 ^ n17161;
  assign n18312 = n18310 & ~n18311;
  assign n18313 = n18312 ^ n17161;
  assign n18314 = n18309 & n18313;
  assign n18315 = n18314 ^ n18304;
  assign n18316 = ~n17263 & n18315;
  assign n18317 = ~n17275 & n18316;
  assign n18318 = n17134 & ~n18317;
  assign n18319 = ~n18307 & ~n18318;
  assign n18320 = n18303 & n18319;
  assign n18321 = n17997 & n18320;
  assign n18322 = ~n17818 & n18321;
  assign n18323 = n17993 & n18322;
  assign n18324 = n18323 ^ n15877;
  assign n18325 = n18324 ^ x720;
  assign n18326 = ~n18298 & n18325;
  assign n18327 = n18269 & n18326;
  assign n18328 = n17377 & ~n17425;
  assign n18329 = ~n17406 & ~n18328;
  assign n18330 = n17409 & ~n17422;
  assign n18331 = n17304 & ~n18096;
  assign n18332 = n17375 & n17377;
  assign n18333 = n17372 ^ n17339;
  assign n18334 = n18333 ^ n17370;
  assign n18335 = n18334 ^ n17373;
  assign n18336 = n17373 ^ n17370;
  assign n18337 = n18336 ^ n17370;
  assign n18338 = n17370 ^ n17339;
  assign n18339 = n18338 ^ n17370;
  assign n18340 = n18337 & n18339;
  assign n18341 = n18340 ^ n17370;
  assign n18342 = ~n18335 & ~n18341;
  assign n18343 = n17429 & ~n18342;
  assign n18344 = ~n17403 & n18343;
  assign n18345 = n17394 & ~n18344;
  assign n18346 = ~n18332 & ~n18345;
  assign n18347 = ~n17424 & ~n17428;
  assign n18348 = n17383 & ~n18347;
  assign n18349 = ~n17390 & ~n17410;
  assign n18350 = ~n17411 & n18349;
  assign n18351 = n17304 & ~n18350;
  assign n18352 = ~n18348 & ~n18351;
  assign n18355 = ~n17395 & n17419;
  assign n18356 = ~n17407 & n18355;
  assign n18353 = ~n17399 & n18092;
  assign n18354 = ~n17411 & n18353;
  assign n18357 = n18356 ^ n18354;
  assign n18358 = n18356 ^ n17303;
  assign n18359 = n18358 ^ n18356;
  assign n18360 = n18357 & n18359;
  assign n18361 = n18360 ^ n18356;
  assign n18362 = ~n18078 & ~n18361;
  assign n18363 = n18352 & ~n18362;
  assign n18364 = n18346 & n18363;
  assign n18365 = ~n17376 & n18364;
  assign n18366 = ~n18331 & n18365;
  assign n18367 = ~n18330 & n18366;
  assign n18368 = n18329 & n18367;
  assign n18369 = ~n18084 & n18368;
  assign n18370 = n18369 ^ n15804;
  assign n18371 = n18370 ^ x721;
  assign n18372 = n18327 & n18371;
  assign n18373 = ~n18325 & n18371;
  assign n18374 = n18298 & n18373;
  assign n18375 = n18269 & n18374;
  assign n18376 = ~n18372 & ~n18375;
  assign n18377 = n18239 & ~n18376;
  assign n18378 = n18298 & n18325;
  assign n18379 = ~n18269 & n18378;
  assign n18380 = ~n18371 & n18379;
  assign n18381 = n18239 & n18380;
  assign n18382 = n18217 & ~n18238;
  assign n18383 = ~n18269 & n18374;
  assign n18384 = n18382 & n18383;
  assign n18385 = ~n18217 & n18238;
  assign n18386 = ~n18298 & n18373;
  assign n18387 = n18269 & n18386;
  assign n18388 = n18298 & ~n18325;
  assign n18389 = n18269 & ~n18371;
  assign n18390 = n18388 & n18389;
  assign n18391 = ~n18387 & ~n18390;
  assign n18392 = n18385 & ~n18391;
  assign n18393 = ~n18384 & ~n18392;
  assign n18394 = ~n18269 & ~n18298;
  assign n18395 = ~n18325 & n18394;
  assign n18396 = ~n18371 & n18395;
  assign n18397 = ~n18380 & ~n18396;
  assign n18398 = n18385 & ~n18397;
  assign n18399 = n18217 & n18238;
  assign n18400 = n18269 & n18378;
  assign n18401 = n18371 & n18400;
  assign n18402 = n18326 & n18389;
  assign n18403 = ~n18401 & ~n18402;
  assign n18404 = n18399 & ~n18403;
  assign n18405 = ~n18398 & ~n18404;
  assign n18406 = n18393 & n18405;
  assign n18407 = n18372 & n18399;
  assign n18408 = n18239 & ~n18391;
  assign n18409 = ~n18407 & ~n18408;
  assign n18410 = n18373 & n18394;
  assign n18411 = n18378 & n18389;
  assign n18412 = ~n18410 & ~n18411;
  assign n18413 = n18385 & ~n18412;
  assign n18414 = n18396 & n18399;
  assign n18415 = n18325 & n18394;
  assign n18416 = ~n18371 & n18415;
  assign n18417 = n18382 & n18416;
  assign n18418 = ~n18414 & ~n18417;
  assign n18419 = n18371 & n18415;
  assign n18420 = n18382 & n18419;
  assign n18421 = ~n18269 & n18388;
  assign n18422 = ~n18371 & n18421;
  assign n18423 = ~n18410 & ~n18422;
  assign n18424 = ~n18380 & n18423;
  assign n18425 = ~n18375 & n18424;
  assign n18426 = n18399 & ~n18425;
  assign n18427 = ~n18420 & ~n18426;
  assign n18428 = n18371 & n18379;
  assign n18429 = ~n18238 & n18428;
  assign n18430 = ~n18372 & ~n18383;
  assign n18431 = n18385 & ~n18430;
  assign n18432 = ~n18396 & ~n18411;
  assign n18433 = n18432 ^ n18217;
  assign n18434 = n18433 ^ n18432;
  assign n18435 = ~n18325 & n18389;
  assign n18436 = ~n18298 & n18435;
  assign n18437 = n18391 & ~n18402;
  assign n18438 = ~n18436 & n18437;
  assign n18439 = n18438 ^ n18432;
  assign n18440 = n18434 & n18439;
  assign n18441 = n18440 ^ n18432;
  assign n18442 = ~n18238 & ~n18441;
  assign n18443 = ~n18431 & ~n18442;
  assign n18444 = ~n18429 & n18443;
  assign n18445 = n18427 & n18444;
  assign n18446 = n18418 & n18445;
  assign n18447 = ~n18413 & n18446;
  assign n18448 = n18409 & n18447;
  assign n18449 = n18406 & n18448;
  assign n18450 = ~n18381 & n18449;
  assign n18451 = ~n18377 & n18450;
  assign n18452 = n18451 ^ n16591;
  assign n18453 = n18452 ^ x763;
  assign n18454 = ~n18183 & n18453;
  assign n18455 = n17955 & n18454;
  assign n18456 = n17123 ^ x705;
  assign n18457 = n17985 ^ x700;
  assign n18458 = n18456 & ~n18457;
  assign n18459 = ~n17555 & n17557;
  assign n18460 = ~n17593 & n18202;
  assign n18461 = ~n18459 & ~n18460;
  assign n18462 = ~n17600 & n18207;
  assign n18463 = n17567 ^ n17557;
  assign n18464 = n18463 ^ n17567;
  assign n18465 = n17583 ^ n17567;
  assign n18466 = ~n18464 & n18465;
  assign n18467 = n18466 ^ n17567;
  assign n18468 = n17556 & n18467;
  assign n18469 = ~n18462 & ~n18468;
  assign n18470 = n18461 & n18469;
  assign n18471 = n18470 ^ n15642;
  assign n18472 = n18471 ^ x702;
  assign n18473 = n17300 ^ x704;
  assign n18474 = ~n18472 & n18473;
  assign n18475 = n17727 & n17733;
  assign n18476 = n17727 & n17734;
  assign n18477 = ~n17705 & ~n17735;
  assign n18478 = n17648 & ~n18477;
  assign n18479 = ~n18476 & ~n18478;
  assign n18480 = ~n17705 & ~n17722;
  assign n18481 = n17727 & ~n18480;
  assign n18482 = n17720 & n17728;
  assign n18483 = n17670 & n17732;
  assign n18484 = ~n17724 & ~n17751;
  assign n18485 = ~n18483 & n18484;
  assign n18486 = ~n17707 & n18485;
  assign n18487 = n17648 & ~n18486;
  assign n18488 = ~n18482 & ~n18487;
  assign n18489 = n17647 & ~n18484;
  assign n18490 = ~n17736 & ~n17754;
  assign n18491 = n17727 & ~n18490;
  assign n18492 = n17702 & ~n17738;
  assign n18493 = ~n17711 & ~n17734;
  assign n18494 = ~n17700 & ~n17707;
  assign n18495 = n18493 & n18494;
  assign n18496 = n17755 & n18495;
  assign n18497 = n17713 & ~n18496;
  assign n18498 = ~n18492 & ~n18497;
  assign n18499 = ~n18491 & n18498;
  assign n18500 = ~n18489 & n18499;
  assign n18501 = n18488 & n18500;
  assign n18502 = ~n18481 & n18501;
  assign n18503 = n18479 & n18502;
  assign n18504 = ~n18475 & n18503;
  assign n18505 = n17710 & n18504;
  assign n18506 = n18505 ^ n15681;
  assign n18507 = n18506 ^ x703;
  assign n18508 = n18474 & ~n18507;
  assign n18509 = n18106 ^ x701;
  assign n18510 = n18508 & ~n18509;
  assign n18511 = n18458 & n18510;
  assign n18512 = ~n18456 & ~n18457;
  assign n18513 = n18473 & n18507;
  assign n18514 = n18472 & n18513;
  assign n18515 = ~n18509 & n18514;
  assign n18516 = n18512 & n18515;
  assign n18517 = ~n18511 & ~n18516;
  assign n18518 = n18456 & n18457;
  assign n18519 = ~n18472 & n18509;
  assign n18520 = ~n18473 & n18519;
  assign n18521 = n18507 & n18520;
  assign n18522 = n18472 & ~n18507;
  assign n18523 = ~n18473 & n18522;
  assign n18524 = n18509 & n18523;
  assign n18525 = n18473 & n18522;
  assign n18526 = n18509 & n18525;
  assign n18527 = ~n18507 & n18520;
  assign n18528 = ~n18526 & ~n18527;
  assign n18529 = ~n18524 & n18528;
  assign n18530 = ~n18521 & n18529;
  assign n18531 = n18518 & ~n18530;
  assign n18532 = n18472 & ~n18473;
  assign n18533 = n18507 & n18532;
  assign n18534 = n18509 & n18533;
  assign n18535 = ~n18473 & ~n18509;
  assign n18536 = n18522 & n18535;
  assign n18537 = ~n18472 & n18535;
  assign n18538 = n18507 & n18537;
  assign n18539 = ~n18536 & ~n18538;
  assign n18540 = ~n18534 & n18539;
  assign n18541 = n18458 & ~n18540;
  assign n18542 = ~n18531 & ~n18541;
  assign n18543 = ~n18472 & n18513;
  assign n18544 = ~n18509 & n18543;
  assign n18545 = ~n18536 & ~n18544;
  assign n18546 = n18512 & ~n18545;
  assign n18547 = ~n18456 & n18457;
  assign n18548 = ~n18507 & n18537;
  assign n18549 = ~n18509 & n18525;
  assign n18550 = ~n18538 & ~n18549;
  assign n18551 = ~n18548 & n18550;
  assign n18552 = n18547 & ~n18551;
  assign n18553 = n18513 & n18519;
  assign n18554 = n18458 & n18553;
  assign n18555 = n18472 & n18535;
  assign n18556 = n18507 & n18555;
  assign n18557 = n18518 & n18556;
  assign n18558 = ~n18554 & ~n18557;
  assign n18559 = n18473 & n18519;
  assign n18560 = ~n18507 & n18559;
  assign n18561 = ~n18521 & ~n18560;
  assign n18562 = n18512 & ~n18561;
  assign n18563 = n18547 & n18553;
  assign n18564 = n18526 & n18547;
  assign n18565 = n18515 & n18518;
  assign n18566 = ~n18564 & ~n18565;
  assign n18567 = n18509 & n18514;
  assign n18568 = ~n18524 & ~n18567;
  assign n18569 = ~n18560 & n18568;
  assign n18570 = n18458 & ~n18569;
  assign n18571 = n18512 & ~n18528;
  assign n18572 = ~n18570 & ~n18571;
  assign n18573 = n18547 & ~n18568;
  assign n18574 = ~n18544 & ~n18548;
  assign n18575 = n18518 & ~n18574;
  assign n18576 = ~n18573 & ~n18575;
  assign n18577 = n18572 & n18576;
  assign n18578 = n18566 & n18577;
  assign n18579 = ~n18563 & n18578;
  assign n18580 = ~n18562 & n18579;
  assign n18581 = n18558 & n18580;
  assign n18582 = ~n18552 & n18581;
  assign n18583 = ~n18546 & n18582;
  assign n18584 = n18542 & n18583;
  assign n18585 = n18517 & n18584;
  assign n18586 = n18510 ^ n18457;
  assign n18587 = n18586 ^ n18510;
  assign n18588 = n18556 ^ n18510;
  assign n18589 = ~n18587 & n18588;
  assign n18590 = n18589 ^ n18510;
  assign n18591 = ~n18456 & n18590;
  assign n18592 = n18585 & ~n18591;
  assign n18593 = n18592 ^ n16825;
  assign n18594 = n18593 ^ x760;
  assign n18595 = n17607 ^ x735;
  assign n18596 = n17065 & ~n17102;
  assign n18597 = n17057 & ~n17090;
  assign n18598 = n17062 & n17103;
  assign n18599 = ~n18597 & ~n18598;
  assign n18600 = ~n18596 & n18599;
  assign n18601 = ~n17014 & ~n17104;
  assign n18602 = n17623 & n18601;
  assign n18603 = n17057 & ~n18602;
  assign n18604 = ~n17092 & n17611;
  assign n18605 = ~n17056 & n18604;
  assign n18606 = n17065 & ~n18605;
  assign n18607 = ~n18603 & ~n18606;
  assign n18608 = n17617 & n18601;
  assign n18609 = ~n17064 & n18608;
  assign n18610 = n17052 & ~n18609;
  assign n18611 = ~n17061 & ~n17093;
  assign n18612 = ~n17101 & ~n18611;
  assign n18613 = n17097 & n17102;
  assign n18614 = n17062 & ~n18613;
  assign n18615 = ~n18612 & ~n18614;
  assign n18616 = ~n18610 & n18615;
  assign n18617 = n18607 & n18616;
  assign n18618 = n17610 & n18617;
  assign n18619 = n17076 & n18618;
  assign n18620 = n18600 & n18619;
  assign n18621 = n18620 ^ n15485;
  assign n18622 = n18621 ^ x730;
  assign n18623 = ~n18595 & n18622;
  assign n18624 = n17839 ^ x734;
  assign n18625 = ~n16479 & ~n18032;
  assign n18626 = n16484 & ~n16501;
  assign n18627 = n16477 & ~n18626;
  assign n18628 = ~n18625 & ~n18627;
  assign n18629 = ~n16488 & n16520;
  assign n18630 = n16361 & ~n18629;
  assign n18631 = n18043 & n18048;
  assign n18632 = n16505 & ~n18631;
  assign n18633 = ~n18630 & ~n18632;
  assign n18634 = n18628 & n18633;
  assign n18635 = n18045 & n18634;
  assign n18636 = ~n18293 & n18635;
  assign n18637 = n18271 & n18636;
  assign n18638 = n16516 & n18637;
  assign n18639 = ~n16490 & n18638;
  assign n18640 = n18639 ^ n16676;
  assign n18641 = n18640 ^ x732;
  assign n18642 = ~n18624 & ~n18641;
  assign n18643 = n17727 & n17735;
  assign n18644 = n17720 & n17724;
  assign n18645 = ~n18643 & ~n18644;
  assign n18646 = n17702 & ~n17756;
  assign n18647 = ~n17716 & n18493;
  assign n18648 = ~n17728 & n18647;
  assign n18649 = n17713 & ~n18648;
  assign n18650 = n17727 & ~n18494;
  assign n18651 = n17717 & ~n17751;
  assign n18652 = n17648 & ~n18651;
  assign n18653 = n17721 & n17732;
  assign n18654 = ~n17736 & n17755;
  assign n18655 = ~n18653 & n18654;
  assign n18656 = n17713 & ~n18655;
  assign n18657 = ~n18652 & ~n18656;
  assign n18658 = n17735 ^ n17646;
  assign n18659 = ~n17711 & ~n17722;
  assign n18660 = n18659 ^ n17700;
  assign n18661 = n17700 ^ n17647;
  assign n18662 = n18661 ^ n17700;
  assign n18663 = ~n18660 & ~n18662;
  assign n18664 = n18663 ^ n17700;
  assign n18665 = n18664 ^ n17735;
  assign n18666 = n18658 & n18665;
  assign n18667 = n18666 ^ n18663;
  assign n18668 = n18667 ^ n17700;
  assign n18669 = n18668 ^ n17646;
  assign n18670 = ~n17735 & n18669;
  assign n18671 = n18670 ^ n17735;
  assign n18672 = n18671 ^ n17646;
  assign n18673 = n18657 & ~n18672;
  assign n18674 = ~n18481 & n18673;
  assign n18675 = ~n18650 & n18674;
  assign n18676 = n17710 & n18675;
  assign n18677 = ~n18649 & n18676;
  assign n18678 = ~n18646 & n18677;
  assign n18679 = n18645 & n18678;
  assign n18680 = ~n18475 & n18679;
  assign n18681 = n18680 ^ n15287;
  assign n18682 = n18681 ^ x731;
  assign n18683 = n17417 & n18092;
  assign n18684 = n17377 & ~n18683;
  assign n18685 = n17419 & ~n17428;
  assign n18686 = ~n17375 & n18685;
  assign n18687 = ~n17380 & n18686;
  assign n18688 = n17394 & ~n18687;
  assign n18689 = ~n18684 & ~n18688;
  assign n18690 = ~n17380 & ~n18342;
  assign n18691 = n17383 & ~n18690;
  assign n18692 = ~n17388 & ~n17411;
  assign n18693 = n17377 & ~n18692;
  assign n18694 = ~n17424 & n18355;
  assign n18695 = ~n17409 & n18694;
  assign n18696 = ~n17411 & n18695;
  assign n18697 = n17304 & ~n18696;
  assign n18698 = ~n18693 & ~n18697;
  assign n18699 = ~n18691 & n18698;
  assign n18700 = n18689 & n18699;
  assign n18701 = ~n17397 & n18700;
  assign n18702 = n18329 & n18701;
  assign n18703 = n18085 & n18702;
  assign n18704 = ~n17376 & n18703;
  assign n18705 = n18704 ^ n16697;
  assign n18706 = n18705 ^ x733;
  assign n18707 = n18682 & ~n18706;
  assign n18708 = n18642 & n18707;
  assign n18709 = n18623 & n18708;
  assign n18710 = n18595 & n18622;
  assign n18711 = n18624 & n18641;
  assign n18712 = ~n18682 & n18706;
  assign n18713 = n18711 & n18712;
  assign n18714 = n18642 & n18712;
  assign n18715 = ~n18713 & ~n18714;
  assign n18716 = n18710 & ~n18715;
  assign n18717 = ~n18709 & ~n18716;
  assign n18718 = n18641 ^ n18624;
  assign n18719 = n18707 & n18718;
  assign n18720 = n18710 & n18719;
  assign n18721 = n18595 & ~n18622;
  assign n18722 = ~n18624 & n18641;
  assign n18723 = n18682 & n18706;
  assign n18724 = n18722 & n18723;
  assign n18725 = n18707 & n18711;
  assign n18726 = ~n18724 & ~n18725;
  assign n18727 = ~n18708 & n18726;
  assign n18728 = n18721 & ~n18727;
  assign n18729 = ~n18720 & ~n18728;
  assign n18730 = ~n18595 & ~n18622;
  assign n18731 = n18712 & n18722;
  assign n18732 = n18624 & ~n18641;
  assign n18733 = n18712 & n18732;
  assign n18734 = ~n18731 & ~n18733;
  assign n18735 = n18730 & ~n18734;
  assign n18736 = ~n18682 & ~n18706;
  assign n18737 = n18722 & n18736;
  assign n18738 = n18711 & n18736;
  assign n18739 = ~n18737 & ~n18738;
  assign n18740 = n18623 & ~n18739;
  assign n18741 = ~n18735 & ~n18740;
  assign n18742 = n18711 & n18723;
  assign n18743 = n18721 & n18742;
  assign n18744 = n18642 & n18736;
  assign n18745 = n18710 & n18744;
  assign n18746 = ~n18743 & ~n18745;
  assign n18747 = n18623 & n18713;
  assign n18748 = n18732 & n18736;
  assign n18749 = n18730 & n18748;
  assign n18750 = ~n18747 & ~n18749;
  assign n18751 = n18642 & n18723;
  assign n18752 = ~n18738 & ~n18748;
  assign n18753 = ~n18751 & n18752;
  assign n18754 = n18721 & ~n18753;
  assign n18755 = n18723 & n18732;
  assign n18756 = ~n18731 & ~n18755;
  assign n18757 = ~n18737 & n18756;
  assign n18758 = n18710 & ~n18757;
  assign n18759 = ~n18751 & ~n18755;
  assign n18760 = ~n18725 & n18759;
  assign n18761 = ~n18730 & n18760;
  assign n18762 = ~n18719 & ~n18751;
  assign n18763 = ~n18623 & n18762;
  assign n18764 = ~n18761 & ~n18763;
  assign n18765 = ~n18744 & ~n18764;
  assign n18766 = ~n18595 & ~n18765;
  assign n18767 = ~n18758 & ~n18766;
  assign n18768 = ~n18754 & n18767;
  assign n18769 = n18750 & n18768;
  assign n18770 = n18746 & n18769;
  assign n18771 = n18742 ^ n18595;
  assign n18772 = n18771 ^ n18742;
  assign n18773 = n18742 ^ n18731;
  assign n18774 = n18772 & n18773;
  assign n18775 = n18774 ^ n18742;
  assign n18776 = ~n18622 & n18775;
  assign n18777 = n18770 & ~n18776;
  assign n18778 = n18741 & n18777;
  assign n18779 = n18729 & n18778;
  assign n18780 = n18717 & n18779;
  assign n18781 = n18780 ^ n16785;
  assign n18782 = n18781 ^ x765;
  assign n18783 = ~n18594 & ~n18782;
  assign n18784 = n18455 & n18783;
  assign n18785 = n17494 & ~n17954;
  assign n18786 = n18454 & n18785;
  assign n18787 = n18594 & n18782;
  assign n18788 = n18786 & n18787;
  assign n18789 = n18183 & ~n18453;
  assign n18790 = n17955 & n18789;
  assign n18791 = n18594 & ~n18782;
  assign n18792 = n18790 & n18791;
  assign n18793 = ~n18788 & ~n18792;
  assign n18794 = ~n18784 & n18793;
  assign n18795 = ~n17494 & n17954;
  assign n18796 = n18789 & n18795;
  assign n18797 = ~n18782 & n18796;
  assign n18798 = n18183 & n18453;
  assign n18799 = n17955 & n18798;
  assign n18800 = ~n18594 & n18782;
  assign n18801 = ~n18791 & ~n18800;
  assign n18802 = n18799 & ~n18801;
  assign n18803 = ~n18797 & ~n18802;
  assign n18804 = n18454 & n18795;
  assign n18805 = ~n18594 & n18804;
  assign n18806 = ~n17494 & ~n17954;
  assign n18807 = n18789 & n18806;
  assign n18808 = n18800 & n18807;
  assign n18809 = ~n18805 & ~n18808;
  assign n18810 = n18454 & n18806;
  assign n18811 = ~n18183 & ~n18453;
  assign n18812 = n18806 & n18811;
  assign n18813 = ~n18810 & ~n18812;
  assign n18814 = n18787 & ~n18813;
  assign n18815 = n18453 ^ n18183;
  assign n18816 = n18183 ^ n17494;
  assign n18817 = n18816 ^ n18183;
  assign n18818 = ~n18815 & ~n18817;
  assign n18819 = n18818 ^ n18183;
  assign n18820 = ~n17954 & ~n18819;
  assign n18821 = ~n18791 & ~n18820;
  assign n18822 = n18798 & n18806;
  assign n18823 = n18785 & n18789;
  assign n18824 = ~n18810 & ~n18823;
  assign n18825 = ~n18822 & n18824;
  assign n18826 = ~n18455 & n18825;
  assign n18827 = ~n18800 & n18826;
  assign n18828 = ~n18821 & ~n18827;
  assign n18829 = ~n18801 & n18828;
  assign n18830 = n17954 & n18811;
  assign n18831 = n18795 & n18798;
  assign n18832 = ~n18790 & ~n18831;
  assign n18833 = ~n18830 & n18832;
  assign n18834 = n18787 & ~n18833;
  assign n18835 = n18785 & n18798;
  assign n18836 = ~n18812 & ~n18835;
  assign n18837 = ~n18807 & n18836;
  assign n18838 = ~n18822 & n18837;
  assign n18839 = n18783 & ~n18838;
  assign n18840 = ~n18834 & ~n18839;
  assign n18841 = ~n18829 & n18840;
  assign n18842 = ~n18814 & n18841;
  assign n18843 = n18809 & n18842;
  assign n18844 = n18803 & n18843;
  assign n18845 = ~n17494 & n18830;
  assign n18846 = n18782 ^ n18594;
  assign n18847 = n18845 & n18846;
  assign n18848 = n18844 & ~n18847;
  assign n18849 = n18794 & n18848;
  assign n18850 = n18823 ^ n18782;
  assign n18851 = n18850 ^ n18823;
  assign n18852 = n17494 & n18830;
  assign n18853 = n18852 ^ n18823;
  assign n18854 = ~n18851 & n18853;
  assign n18855 = n18854 ^ n18823;
  assign n18856 = ~n18846 & n18855;
  assign n18857 = n18849 & ~n18856;
  assign n18858 = n18857 ^ n17985;
  assign n18859 = ~n16903 & ~n17129;
  assign n18860 = n17449 ^ n17124;
  assign n18861 = n18860 ^ n17449;
  assign n18862 = n17456 ^ n17449;
  assign n18863 = n18861 & ~n18862;
  assign n18864 = n18863 ^ n17449;
  assign n18865 = ~n18859 & ~n18864;
  assign n18866 = n17446 & n18865;
  assign n18867 = n17486 ^ n17129;
  assign n18868 = ~n17124 & ~n18867;
  assign n18869 = n18868 ^ n17129;
  assign n18870 = n17448 & n18869;
  assign n18871 = ~n18866 & ~n18870;
  assign n18872 = n17445 ^ n17301;
  assign n18873 = n16539 & ~n17467;
  assign n18874 = ~n16539 & n17467;
  assign n18875 = n18874 ^ n17124;
  assign n18876 = n18875 ^ n18874;
  assign n18877 = n18874 ^ n16904;
  assign n18878 = n18877 ^ n18874;
  assign n18879 = n18876 & ~n18878;
  assign n18880 = n18879 ^ n18874;
  assign n18881 = ~n16190 & n18880;
  assign n18882 = n18881 ^ n18874;
  assign n18883 = ~n18873 & ~n18882;
  assign n18884 = n18883 ^ n17445;
  assign n18885 = n18884 ^ n18883;
  assign n18886 = n17483 & ~n18874;
  assign n18887 = n18886 ^ n18883;
  assign n18888 = n18885 & ~n18887;
  assign n18889 = n18888 ^ n18883;
  assign n18890 = ~n18872 & n18889;
  assign n18891 = n18871 & ~n18890;
  assign n18892 = n18891 ^ n16442;
  assign n18893 = n18892 ^ x750;
  assign n18894 = n17880 & n17900;
  assign n18895 = n17882 & n17917;
  assign n18896 = ~n18894 & ~n18895;
  assign n18897 = ~n17914 & n18896;
  assign n18898 = ~n17906 & ~n17915;
  assign n18899 = n17882 & ~n18898;
  assign n18900 = n17908 & ~n18899;
  assign n18901 = n17882 & n17923;
  assign n18902 = n17903 & n17905;
  assign n18903 = ~n18901 & ~n18902;
  assign n18904 = ~n17879 & n17922;
  assign n18905 = ~n17887 & n17916;
  assign n18906 = n17880 & ~n18905;
  assign n18907 = ~n17815 & ~n17924;
  assign n18908 = n17905 & ~n18907;
  assign n18909 = ~n18906 & ~n18908;
  assign n18910 = ~n18904 & n18909;
  assign n18911 = n17894 & ~n17929;
  assign n18912 = n17882 & ~n18911;
  assign n18913 = n17644 ^ n17608;
  assign n18914 = n18913 ^ n17644;
  assign n18915 = n18914 ^ n18913;
  assign n18916 = n18913 ^ n17813;
  assign n18917 = n18915 & n18916;
  assign n18918 = n18917 ^ n18913;
  assign n18919 = n17772 & n18918;
  assign n18920 = n18919 ^ n18913;
  assign n18921 = n17884 & n18920;
  assign n18922 = ~n18912 & ~n18921;
  assign n18923 = n18910 & n18922;
  assign n18924 = n17912 & n18923;
  assign n18925 = n18903 & n18924;
  assign n18926 = n18900 & n18925;
  assign n18927 = n18897 & n18926;
  assign n18928 = ~n17881 & n18927;
  assign n18929 = ~n17897 & n18928;
  assign n18930 = n18929 ^ n16472;
  assign n18931 = n18930 ^ x749;
  assign n18932 = n18893 & n18931;
  assign n18933 = n18297 ^ x724;
  assign n18934 = n18681 ^ x729;
  assign n18935 = ~n18933 & n18934;
  assign n18936 = n18621 ^ x728;
  assign n18937 = n18237 ^ x725;
  assign n18938 = ~n18936 & n18937;
  assign n18939 = n17558 & ~n18199;
  assign n18940 = n17569 & ~n18193;
  assign n18941 = ~n18939 & ~n18940;
  assign n18942 = n18202 & n18212;
  assign n18943 = ~n18205 & n18207;
  assign n18944 = ~n18942 & ~n18943;
  assign n18945 = n18941 & n18944;
  assign n18946 = n18945 ^ n15421;
  assign n18947 = n18946 ^ x726;
  assign n18948 = n15950 ^ n15598;
  assign n18949 = n15950 ^ n15750;
  assign n18950 = n18949 ^ n15950;
  assign n18951 = n18948 & ~n18950;
  assign n18952 = n18951 ^ n15950;
  assign n18953 = n16114 & n18952;
  assign n18954 = n16127 & n18953;
  assign n18955 = ~n16142 & ~n16178;
  assign n18956 = n15220 & ~n18955;
  assign n18957 = ~n16118 & ~n16139;
  assign n18958 = ~n16134 & ~n18957;
  assign n18959 = n16119 & n17859;
  assign n18960 = n16121 & ~n18959;
  assign n18961 = ~n18958 & ~n18960;
  assign n18962 = n15220 & ~n17849;
  assign n18963 = n16121 & ~n17848;
  assign n18964 = n16182 & ~n18963;
  assign n18965 = n15219 & ~n18964;
  assign n18966 = ~n18962 & ~n18965;
  assign n18967 = n18961 & n18966;
  assign n18968 = ~n18956 & n18967;
  assign n18969 = ~n18954 & n18968;
  assign n18970 = n17844 & n18969;
  assign n18971 = n18243 & n18970;
  assign n18972 = n16150 & n18971;
  assign n18973 = n18972 ^ n15517;
  assign n18974 = n18973 ^ x727;
  assign n18975 = ~n18947 & ~n18974;
  assign n18976 = n18938 & n18975;
  assign n18977 = n18936 & n18937;
  assign n18978 = n18947 & ~n18974;
  assign n18979 = n18977 & n18978;
  assign n18980 = ~n18976 & ~n18979;
  assign n18981 = n18935 & ~n18980;
  assign n18982 = ~n18936 & ~n18937;
  assign n18983 = ~n18947 & n18974;
  assign n18984 = n18982 & n18983;
  assign n18985 = n18935 & n18984;
  assign n18986 = n18938 & n18978;
  assign n18987 = n18933 & n18934;
  assign n18988 = n18986 & n18987;
  assign n18989 = ~n18985 & ~n18988;
  assign n18990 = n18938 & n18983;
  assign n18991 = n18947 & n18974;
  assign n18992 = n18938 & n18991;
  assign n18993 = n18975 & n18977;
  assign n18994 = ~n18992 & ~n18993;
  assign n18995 = n18936 & ~n18937;
  assign n18996 = n18978 & n18995;
  assign n18997 = ~n18984 & ~n18996;
  assign n18998 = n18991 & n18995;
  assign n18999 = n18975 & n18982;
  assign n19000 = ~n18998 & ~n18999;
  assign n19001 = n18997 & n19000;
  assign n19002 = n18994 & n19001;
  assign n19003 = ~n18990 & n19002;
  assign n19004 = n18987 & ~n19003;
  assign n19005 = ~n18933 & ~n18934;
  assign n19006 = n18982 & n18991;
  assign n19007 = n18975 & n18995;
  assign n19008 = ~n19006 & ~n19007;
  assign n19009 = n18977 & n18983;
  assign n19010 = ~n18992 & ~n19009;
  assign n19011 = n18997 & n19010;
  assign n19012 = ~n18993 & n19011;
  assign n19013 = n19008 & n19012;
  assign n19014 = ~n18986 & n19013;
  assign n19015 = n19005 & ~n19014;
  assign n19016 = ~n19004 & ~n19015;
  assign n19017 = n18934 ^ n18933;
  assign n19018 = n18983 & n18995;
  assign n19019 = ~n18990 & ~n19018;
  assign n19020 = n19008 & n19019;
  assign n19021 = ~n18996 & n19020;
  assign n19022 = n19021 ^ n18934;
  assign n19023 = n19022 ^ n19021;
  assign n19024 = ~n18979 & n18994;
  assign n19025 = n19001 & n19024;
  assign n19026 = ~n19018 & n19025;
  assign n19027 = n19026 ^ n19021;
  assign n19028 = ~n19023 & ~n19027;
  assign n19029 = n19028 ^ n19021;
  assign n19030 = n19017 & ~n19029;
  assign n19031 = n19016 & ~n19030;
  assign n19032 = n18989 & n19031;
  assign n19033 = ~n18981 & n19032;
  assign n19034 = n19033 ^ n16386;
  assign n19035 = n19034 ^ x752;
  assign n19036 = ~n18380 & ~n18419;
  assign n19037 = n18399 & ~n19036;
  assign n19038 = ~n18416 & ~n18428;
  assign n19039 = n18385 & ~n19038;
  assign n19040 = ~n19037 & ~n19039;
  assign n19041 = ~n18239 & ~n18399;
  assign n19042 = ~n18403 & n19041;
  assign n19043 = ~n18387 & n18397;
  assign n19044 = ~n18375 & n19043;
  assign n19045 = n18382 & ~n19044;
  assign n19046 = ~n18390 & ~n18436;
  assign n19047 = n18423 & n19046;
  assign n19048 = ~n18428 & n19047;
  assign n19049 = n18239 & ~n19048;
  assign n19050 = ~n19045 & ~n19049;
  assign n19051 = ~n19042 & n19050;
  assign n19052 = ~n18411 & ~n18436;
  assign n19053 = ~n18410 & n19052;
  assign n19054 = ~n18383 & n19053;
  assign n19055 = n19054 ^ n18419;
  assign n19056 = n19055 ^ n18419;
  assign n19057 = n18419 ^ n18217;
  assign n19058 = n19057 ^ n18419;
  assign n19059 = ~n19056 & n19058;
  assign n19060 = n19059 ^ n18419;
  assign n19061 = n18238 & n19060;
  assign n19062 = n19061 ^ n18419;
  assign n19063 = n19051 & ~n19062;
  assign n19064 = n18406 & n19063;
  assign n19065 = n19040 & n19064;
  assign n19066 = ~n18377 & n19065;
  assign n19067 = n19066 ^ n16425;
  assign n19068 = n19067 ^ x751;
  assign n19069 = ~n19035 & n19068;
  assign n19070 = n18932 & n19069;
  assign n19071 = n19035 & ~n19068;
  assign n19072 = n18932 & n19071;
  assign n19073 = ~n19070 & ~n19072;
  assign n19074 = n18108 & ~n18116;
  assign n19075 = n18110 & n18135;
  assign n19076 = ~n18131 & ~n18166;
  assign n19077 = n18119 & ~n19076;
  assign n19078 = ~n19075 & ~n19077;
  assign n19079 = ~n19074 & n19078;
  assign n19080 = n18119 & n18148;
  assign n19081 = n18110 & n18141;
  assign n19082 = ~n19080 & ~n19081;
  assign n19083 = n18108 & n18161;
  assign n19084 = n18119 & n18152;
  assign n19085 = ~n19083 & ~n19084;
  assign n19086 = n18119 & n18146;
  assign n19087 = n18107 ^ n18076;
  assign n19088 = n18126 & ~n19087;
  assign n19089 = ~n19086 & ~n19088;
  assign n19090 = n18110 & ~n18159;
  assign n19091 = ~n18134 & ~n18162;
  assign n19092 = n18108 & ~n19091;
  assign n19093 = n18136 & n18164;
  assign n19094 = n18123 & ~n19093;
  assign n19095 = ~n19092 & ~n19094;
  assign n19096 = ~n19090 & n19095;
  assign n19097 = n19089 & n19096;
  assign n19098 = n18128 & n19097;
  assign n19099 = n19085 & n19098;
  assign n19100 = n19082 & n19099;
  assign n19101 = n18139 & n19100;
  assign n19102 = n19079 & n19101;
  assign n19103 = n18118 & n19102;
  assign n19104 = n19103 ^ n16223;
  assign n19105 = n19104 ^ x753;
  assign n19106 = n16538 ^ x712;
  assign n19107 = n18268 ^ x717;
  assign n19108 = n19106 & ~n19107;
  assign n19109 = n17061 & n17065;
  assign n19110 = n17062 & ~n17617;
  assign n19111 = ~n19109 & ~n19110;
  assign n19112 = n17052 & ~n17090;
  assign n19113 = ~n17084 & ~n17096;
  assign n19114 = n17057 & ~n19113;
  assign n19115 = ~n17070 & ~n17104;
  assign n19116 = ~n17064 & n19115;
  assign n19117 = ~n17056 & n19116;
  assign n19118 = n17057 & ~n19117;
  assign n19119 = n17065 & ~n18608;
  assign n19120 = ~n19118 & ~n19119;
  assign n19121 = n17611 & n17617;
  assign n19122 = n17052 & ~n19121;
  assign n19123 = n17085 & ~n17096;
  assign n19124 = ~n17093 & n19123;
  assign n19125 = n17062 & ~n19124;
  assign n19126 = ~n19122 & ~n19125;
  assign n19127 = n19120 & n19126;
  assign n19128 = ~n19114 & n19127;
  assign n19129 = ~n19112 & n19128;
  assign n19130 = n19111 & n19129;
  assign n19131 = n17075 & n19130;
  assign n19132 = n17622 & n19131;
  assign n19133 = n18600 & n19132;
  assign n19134 = n19133 ^ n16256;
  assign n19135 = n19134 ^ x714;
  assign n19136 = n17646 & n17716;
  assign n19137 = n17727 & ~n17755;
  assign n19138 = ~n19136 & ~n19137;
  assign n19139 = ~n17724 & n18654;
  assign n19140 = n17648 & ~n19139;
  assign n19141 = ~n17728 & n18494;
  assign n19142 = n17647 & ~n19141;
  assign n19143 = ~n17735 & n17756;
  assign n19144 = n17713 & ~n19143;
  assign n19145 = ~n19142 & ~n19144;
  assign n19146 = n17648 & ~n18493;
  assign n19147 = ~n17733 & n18484;
  assign n19148 = ~n17722 & n19147;
  assign n19149 = n17702 & ~n19148;
  assign n19150 = ~n19146 & ~n19149;
  assign n19151 = n19145 & n19150;
  assign n19152 = ~n19140 & n19151;
  assign n19153 = n19138 & n19152;
  assign n19154 = n18479 & n19153;
  assign n19155 = ~n18650 & n19154;
  assign n19156 = ~n18475 & n19155;
  assign n19157 = n19156 ^ n16280;
  assign n19158 = n19157 ^ x715;
  assign n19159 = n19135 & ~n19158;
  assign n19160 = n18216 ^ x716;
  assign n19161 = n17444 ^ x713;
  assign n19162 = n19160 & n19161;
  assign n19163 = n19159 & n19162;
  assign n19164 = n19108 & n19163;
  assign n19165 = ~n19135 & n19158;
  assign n19166 = n19160 & ~n19161;
  assign n19167 = n19165 & n19166;
  assign n19168 = n19108 & n19167;
  assign n19169 = n19106 & n19107;
  assign n19170 = ~n19160 & ~n19161;
  assign n19171 = n19159 & n19170;
  assign n19172 = n19169 & n19171;
  assign n19173 = ~n19168 & ~n19172;
  assign n19174 = ~n19164 & n19173;
  assign n19175 = ~n19160 & n19161;
  assign n19176 = n19159 & n19175;
  assign n19177 = n19108 & n19176;
  assign n19178 = ~n19106 & ~n19107;
  assign n19179 = ~n19135 & ~n19158;
  assign n19180 = n19161 & n19179;
  assign n19181 = ~n19160 & n19180;
  assign n19182 = ~n19163 & ~n19181;
  assign n19183 = n19178 & ~n19182;
  assign n19184 = ~n19177 & ~n19183;
  assign n19185 = ~n19106 & n19107;
  assign n19186 = n19167 & n19185;
  assign n19187 = n19159 & n19166;
  assign n19188 = n19135 & n19158;
  assign n19189 = n19166 & n19188;
  assign n19190 = ~n19187 & ~n19189;
  assign n19191 = n19178 & ~n19190;
  assign n19192 = ~n19186 & ~n19191;
  assign n19193 = n19165 & n19170;
  assign n19194 = n19185 & n19193;
  assign n19195 = n19108 & n19171;
  assign n19196 = n19167 & n19169;
  assign n19197 = ~n19195 & ~n19196;
  assign n19198 = ~n19194 & n19197;
  assign n19199 = n19185 & n19187;
  assign n19200 = n19169 & n19193;
  assign n19201 = ~n19199 & ~n19200;
  assign n19202 = n19165 & n19175;
  assign n19203 = ~n19107 & n19202;
  assign n19204 = n19170 & n19188;
  assign n19205 = n19178 & n19204;
  assign n19206 = ~n19203 & ~n19205;
  assign n19207 = n19170 & n19179;
  assign n19208 = n19185 & n19207;
  assign n19209 = n19162 & n19188;
  assign n19210 = ~n19176 & ~n19209;
  assign n19211 = ~n19180 & n19210;
  assign n19212 = n19169 & ~n19211;
  assign n19213 = ~n19208 & ~n19212;
  assign n19214 = n19206 & n19213;
  assign n19215 = n19162 & n19165;
  assign n19216 = ~n19106 & n19215;
  assign n19218 = ~n19108 & ~n19185;
  assign n19217 = n19166 & n19179;
  assign n19219 = n19218 ^ n19217;
  assign n19220 = n19219 ^ n19217;
  assign n19221 = n19160 & n19180;
  assign n19222 = n19175 & n19188;
  assign n19223 = ~n19221 & ~n19222;
  assign n19224 = ~n19189 & n19223;
  assign n19225 = n19224 ^ n19217;
  assign n19226 = ~n19220 & ~n19225;
  assign n19227 = n19226 ^ n19217;
  assign n19228 = ~n19216 & ~n19227;
  assign n19229 = n19214 & n19228;
  assign n19230 = n19201 & n19229;
  assign n19231 = n19198 & n19230;
  assign n19232 = n19192 & n19231;
  assign n19233 = n19184 & n19232;
  assign n19234 = n19174 & n19233;
  assign n19235 = n19234 ^ n16359;
  assign n19236 = n19235 ^ x748;
  assign n19237 = ~n19105 & ~n19236;
  assign n19238 = ~n19073 & n19237;
  assign n19239 = ~n19035 & ~n19068;
  assign n19240 = n18932 & n19239;
  assign n19241 = n19105 & n19236;
  assign n19242 = n19240 & n19241;
  assign n19243 = n18893 & ~n18931;
  assign n19244 = n19071 & n19243;
  assign n19245 = ~n18893 & ~n18931;
  assign n19246 = n19239 & n19245;
  assign n19247 = ~n19244 & ~n19246;
  assign n19248 = n19105 & ~n19236;
  assign n19249 = ~n19247 & n19248;
  assign n19250 = ~n19242 & ~n19249;
  assign n19251 = n19069 & n19245;
  assign n19252 = ~n19246 & ~n19251;
  assign n19253 = n19237 & ~n19252;
  assign n19254 = n19035 & n19068;
  assign n19255 = n19243 & n19254;
  assign n19256 = n19241 & n19255;
  assign n19257 = ~n18893 & n18931;
  assign n19258 = n19069 & n19257;
  assign n19259 = ~n19072 & ~n19258;
  assign n19260 = n19248 & ~n19259;
  assign n19261 = ~n19256 & ~n19260;
  assign n19262 = n19245 & n19254;
  assign n19263 = n19241 & n19262;
  assign n19264 = n19254 & n19257;
  assign n19265 = n19236 ^ n19105;
  assign n19266 = n19264 & n19265;
  assign n19267 = ~n19263 & ~n19266;
  assign n19268 = n19239 & n19243;
  assign n19269 = ~n19105 & n19236;
  assign n19270 = ~n19241 & ~n19269;
  assign n19271 = n19268 & ~n19270;
  assign n19272 = n18932 & n19254;
  assign n19273 = n19239 & n19257;
  assign n19274 = ~n19272 & ~n19273;
  assign n19275 = n19274 ^ n19236;
  assign n19276 = n19275 ^ n19274;
  assign n19277 = ~n19255 & ~n19262;
  assign n19278 = ~n19240 & n19277;
  assign n19279 = n19278 ^ n19274;
  assign n19280 = n19279 ^ n19274;
  assign n19281 = ~n19276 & ~n19280;
  assign n19282 = n19281 ^ n19274;
  assign n19283 = ~n19265 & ~n19282;
  assign n19284 = n19283 ^ n19274;
  assign n19285 = ~n19271 & n19284;
  assign n19286 = n19069 & n19243;
  assign n19287 = n19071 & n19245;
  assign n19288 = ~n19286 & ~n19287;
  assign n19289 = n19269 & ~n19288;
  assign n19290 = n19071 & n19257;
  assign n19291 = ~n19070 & ~n19290;
  assign n19292 = ~n19273 & n19291;
  assign n19293 = n19241 & ~n19292;
  assign n19294 = ~n19289 & ~n19293;
  assign n19295 = n19290 ^ n19236;
  assign n19296 = n19295 ^ n19290;
  assign n19297 = n19290 ^ n19286;
  assign n19298 = n19297 ^ n19290;
  assign n19299 = ~n19296 & n19298;
  assign n19300 = n19299 ^ n19290;
  assign n19301 = n19105 & n19300;
  assign n19302 = n19301 ^ n19290;
  assign n19303 = n19294 & ~n19302;
  assign n19304 = n19285 & n19303;
  assign n19305 = n19267 & n19304;
  assign n19306 = n19261 & n19305;
  assign n19307 = ~n19253 & n19306;
  assign n19308 = n19250 & n19307;
  assign n19309 = ~n19238 & n19308;
  assign n19310 = n19251 ^ n19105;
  assign n19311 = n19310 ^ n19251;
  assign n19312 = n19251 ^ n19244;
  assign n19313 = ~n19311 & n19312;
  assign n19314 = n19313 ^ n19251;
  assign n19315 = n19236 & n19314;
  assign n19316 = n19309 & ~n19315;
  assign n19317 = n19316 ^ n16538;
  assign n19318 = n19317 ^ x808;
  assign n19319 = n17475 & ~n18865;
  assign n19320 = n17464 & n18869;
  assign n19321 = ~n19319 & ~n19320;
  assign n19322 = ~n17482 & ~n18874;
  assign n19323 = n19322 ^ n17445;
  assign n19324 = n19323 ^ n19322;
  assign n19325 = n19322 ^ n18883;
  assign n19326 = n19324 & n19325;
  assign n19327 = n19326 ^ n19322;
  assign n19328 = n18872 & ~n19327;
  assign n19329 = n19321 & ~n19328;
  assign n19330 = ~n17477 & n19329;
  assign n19331 = n19330 ^ n14782;
  assign n19332 = n19331 ^ x783;
  assign n19333 = ~n18122 & ~n18126;
  assign n19334 = n18110 & ~n19333;
  assign n19335 = ~n18131 & n18136;
  assign n19336 = n18108 & ~n19335;
  assign n19337 = ~n19334 & ~n19336;
  assign n19338 = n18123 & n18152;
  assign n19339 = ~n18141 & ~n18161;
  assign n19340 = ~n19087 & ~n19339;
  assign n19341 = ~n19338 & ~n19340;
  assign n19342 = ~n18115 & n18136;
  assign n19343 = n18119 & ~n19342;
  assign n19346 = ~n18112 & n18164;
  assign n19344 = ~n18075 & n18163;
  assign n19345 = ~n18166 & n19344;
  assign n19347 = n19346 ^ n19345;
  assign n19348 = n19346 ^ n18107;
  assign n19349 = n19348 ^ n19346;
  assign n19350 = n19347 & n19349;
  assign n19351 = n19350 ^ n19346;
  assign n19352 = n18076 & ~n19351;
  assign n19353 = ~n19343 & ~n19352;
  assign n19354 = n19341 & n19353;
  assign n19355 = n18148 ^ n18108;
  assign n19356 = n18147 ^ n18110;
  assign n19357 = n18147 ^ n18108;
  assign n19358 = n19357 ^ n18147;
  assign n19359 = ~n19356 & ~n19358;
  assign n19360 = n19359 ^ n18147;
  assign n19361 = n19355 & n19360;
  assign n19362 = n19361 ^ n18148;
  assign n19363 = n19354 & ~n19362;
  assign n19364 = n19337 & n19363;
  assign n19365 = n19079 & n19364;
  assign n19366 = n18129 & n19365;
  assign n19367 = n19366 ^ n15218;
  assign n19368 = n19367 ^ x778;
  assign n19369 = ~n19332 & ~n19368;
  assign n19370 = n18978 & n18982;
  assign n19371 = ~n19007 & ~n19370;
  assign n19372 = n18933 & ~n19371;
  assign n19373 = n19001 & n19010;
  assign n19374 = n18935 & ~n19373;
  assign n19375 = n18933 & ~n18934;
  assign n19376 = ~n18976 & n19012;
  assign n19377 = n19375 & ~n19376;
  assign n19378 = ~n19374 & ~n19377;
  assign n19379 = ~n19372 & n19378;
  assign n19380 = ~n18999 & n19019;
  assign n19381 = n19024 & n19380;
  assign n19382 = n19381 ^ n18934;
  assign n19383 = n19382 ^ n19381;
  assign n19384 = n19381 ^ n19026;
  assign n19385 = ~n19383 & ~n19384;
  assign n19386 = n19385 ^ n19381;
  assign n19387 = ~n19017 & ~n19386;
  assign n19388 = n19379 & ~n19387;
  assign n19389 = ~n18981 & n19388;
  assign n19390 = n19389 ^ n15597;
  assign n19391 = n19390 ^ x782;
  assign n19392 = n17880 & n17924;
  assign n19393 = ~n17815 & ~n17923;
  assign n19394 = n17905 & ~n19393;
  assign n19395 = ~n19392 & ~n19394;
  assign n19396 = n17884 & n17913;
  assign n19397 = n17882 & n17887;
  assign n19398 = ~n19396 & ~n19397;
  assign n19399 = ~n17893 & ~n17922;
  assign n19400 = n17882 & ~n19399;
  assign n19401 = ~n17909 & ~n17922;
  assign n19402 = n17918 & n19401;
  assign n19403 = ~n17897 & n19402;
  assign n19404 = n17880 & ~n19403;
  assign n19405 = ~n19400 & ~n19404;
  assign n19406 = n17894 & ~n17906;
  assign n19407 = ~n17887 & n19406;
  assign n19408 = n17905 & ~n19407;
  assign n19409 = ~n17917 & ~n17924;
  assign n19410 = ~n17903 & n19409;
  assign n19411 = n17916 & n19410;
  assign n19412 = ~n17929 & n19411;
  assign n19413 = n17884 & ~n19412;
  assign n19414 = ~n19408 & ~n19413;
  assign n19415 = n19405 & n19414;
  assign n19416 = n17889 & n19415;
  assign n19417 = ~n17902 & n19416;
  assign n19418 = n19398 & n19417;
  assign n19419 = n19395 & n19418;
  assign n19420 = n18903 & n19419;
  assign n19421 = n18897 & n19420;
  assign n19422 = ~n17881 & n19421;
  assign n19423 = n19422 ^ n16113;
  assign n19424 = n19423 ^ x781;
  assign n19425 = ~n19391 & n19424;
  assign n19426 = n18518 & n18549;
  assign n19427 = n18473 ^ n18472;
  assign n19428 = n19427 ^ n18509;
  assign n19429 = n18509 ^ n18473;
  assign n19430 = n18507 ^ n18473;
  assign n19431 = n19430 ^ n18473;
  assign n19432 = n19429 & n19431;
  assign n19433 = n19432 ^ n18473;
  assign n19434 = n19428 & n19433;
  assign n19435 = n18512 & n19434;
  assign n19436 = ~n19426 & ~n19435;
  assign n19437 = ~n18515 & ~n18534;
  assign n19438 = ~n18512 & n19437;
  assign n19439 = n19438 ^ n18547;
  assign n19440 = n19438 ^ n18569;
  assign n19441 = n19440 ^ n18569;
  assign n19442 = n18569 ^ n18550;
  assign n19443 = ~n19441 & ~n19442;
  assign n19444 = n19443 ^ n18569;
  assign n19445 = ~n19439 & n19444;
  assign n19446 = n19445 ^ n18547;
  assign n19447 = ~n18521 & n18569;
  assign n19448 = n18518 & ~n19447;
  assign n19451 = ~n18548 & ~n18560;
  assign n19449 = n18545 & ~n18556;
  assign n19450 = ~n18549 & n19449;
  assign n19452 = n19451 ^ n19450;
  assign n19453 = n19451 ^ n18458;
  assign n19454 = n19451 & n19453;
  assign n19455 = n19454 ^ n19451;
  assign n19456 = n19452 & n19455;
  assign n19457 = n19456 ^ n19454;
  assign n19458 = n19457 ^ n19451;
  assign n19459 = n19458 ^ n18458;
  assign n19460 = ~n19448 & n19459;
  assign n19461 = n19460 ^ n19448;
  assign n19462 = ~n19446 & ~n19461;
  assign n19463 = n19436 & n19462;
  assign n19464 = n18534 ^ n18457;
  assign n19465 = n19464 ^ n18534;
  assign n19466 = n18545 ^ n18534;
  assign n19467 = n19465 & ~n19466;
  assign n19468 = n19467 ^ n18534;
  assign n19469 = n18456 & n19468;
  assign n19470 = n19463 & ~n19469;
  assign n19471 = ~n18563 & n19470;
  assign n19472 = ~n18591 & n19471;
  assign n19473 = n18558 & n19472;
  assign n19474 = ~n18536 & n19473;
  assign n19475 = n19474 ^ n15749;
  assign n19476 = n19475 ^ x780;
  assign n19477 = n18239 & n18419;
  assign n19478 = ~n18396 & ~n18422;
  assign n19479 = ~n18238 & ~n19478;
  assign n19480 = ~n19477 & ~n19479;
  assign n19481 = ~n18383 & ~n18402;
  assign n19482 = ~n19041 & ~n19481;
  assign n19483 = ~n18375 & ~n18436;
  assign n19484 = n18385 & ~n19483;
  assign n19485 = ~n18372 & n18391;
  assign n19486 = n18399 & ~n19485;
  assign n19487 = ~n18387 & n19052;
  assign n19488 = ~n18401 & n19487;
  assign n19489 = n18382 & ~n19488;
  assign n19490 = ~n19486 & ~n19489;
  assign n19491 = ~n19484 & n19490;
  assign n19492 = ~n19482 & n19491;
  assign n19493 = n19480 & n19492;
  assign n19494 = n18418 & n19493;
  assign n19495 = ~n18413 & n19494;
  assign n19496 = n18393 & n19495;
  assign n19497 = n19040 & n19496;
  assign n19498 = ~n18381 & n19497;
  assign n19499 = ~n18377 & n19498;
  assign n19500 = n19499 ^ n15949;
  assign n19501 = n19500 ^ x779;
  assign n19502 = n19476 & ~n19501;
  assign n19503 = n19425 & n19502;
  assign n19504 = n19391 & n19424;
  assign n19505 = ~n19476 & ~n19501;
  assign n19506 = n19504 & n19505;
  assign n19507 = ~n19503 & ~n19506;
  assign n19508 = n19369 & ~n19507;
  assign n19509 = n19332 & ~n19368;
  assign n19510 = ~n19391 & ~n19424;
  assign n19511 = ~n19476 & n19501;
  assign n19512 = n19510 & n19511;
  assign n19513 = n19391 & ~n19424;
  assign n19514 = n19501 & n19513;
  assign n19515 = n19476 & n19514;
  assign n19516 = n19476 & n19501;
  assign n19517 = n19425 & n19516;
  assign n19518 = ~n19515 & ~n19517;
  assign n19519 = ~n19512 & n19518;
  assign n19520 = n19509 & ~n19519;
  assign n19521 = n19425 & n19511;
  assign n19522 = n19504 & n19516;
  assign n19523 = ~n19521 & ~n19522;
  assign n19524 = n19369 & ~n19523;
  assign n19525 = n19505 & n19513;
  assign n19526 = ~n19503 & ~n19525;
  assign n19527 = n19509 & ~n19526;
  assign n19528 = ~n19524 & ~n19527;
  assign n19529 = ~n19332 & n19368;
  assign n19530 = n19521 & n19529;
  assign n19531 = n19332 & n19368;
  assign n19532 = ~n19476 & n19514;
  assign n19533 = n19510 & n19516;
  assign n19534 = ~n19532 & ~n19533;
  assign n19535 = n19531 & ~n19534;
  assign n19536 = ~n19530 & ~n19535;
  assign n19537 = n19502 & n19510;
  assign n19538 = n19531 & n19537;
  assign n19539 = ~n19512 & ~n19515;
  assign n19540 = n19529 & ~n19539;
  assign n19541 = ~n19538 & ~n19540;
  assign n19542 = n19504 & n19511;
  assign n19543 = n19368 & n19542;
  assign n19544 = n19502 & n19513;
  assign n19545 = n19523 & ~n19544;
  assign n19546 = n19509 & ~n19545;
  assign n19547 = n19505 & n19510;
  assign n19548 = ~n19525 & ~n19547;
  assign n19549 = n19534 & n19548;
  assign n19550 = n19369 & ~n19549;
  assign n19551 = n19502 & n19504;
  assign n19552 = n19425 & n19505;
  assign n19553 = ~n19551 & ~n19552;
  assign n19554 = ~n19529 & n19553;
  assign n19555 = ~n19503 & n19554;
  assign n19556 = ~n19537 & ~n19544;
  assign n19557 = ~n19551 & n19556;
  assign n19558 = ~n19531 & n19557;
  assign n19559 = ~n19555 & ~n19558;
  assign n19560 = ~n19547 & ~n19559;
  assign n19561 = n19368 & ~n19560;
  assign n19562 = ~n19550 & ~n19561;
  assign n19563 = ~n19546 & n19562;
  assign n19564 = ~n19543 & n19563;
  assign n19565 = n19541 & n19564;
  assign n19566 = n19536 & n19565;
  assign n19567 = n19528 & n19566;
  assign n19568 = ~n19520 & n19567;
  assign n19569 = ~n19508 & n19568;
  assign n19570 = n19569 ^ n18268;
  assign n19571 = n19570 ^ x813;
  assign n19572 = ~n19318 & n19571;
  assign n19573 = n17953 ^ x759;
  assign n19651 = n19034 ^ x754;
  assign n19609 = ~n18641 & n18707;
  assign n19610 = ~n18725 & ~n19609;
  assign n19611 = n18734 & n19610;
  assign n19612 = n18721 & ~n19611;
  assign n19613 = n18710 & n18748;
  assign n19614 = n18641 & n18723;
  assign n19615 = ~n18733 & ~n19614;
  assign n19616 = ~n18714 & n19615;
  assign n19617 = ~n18755 & n19616;
  assign n19618 = n18623 & ~n19617;
  assign n19619 = ~n19613 & ~n19618;
  assign n19620 = ~n19612 & n19619;
  assign n19621 = ~n18721 & ~n18730;
  assign n19622 = ~n18713 & ~n18737;
  assign n19623 = ~n19621 & ~n19622;
  assign n19624 = ~n18710 & ~n18730;
  assign n19625 = ~n18730 & n19609;
  assign n19626 = n19625 ^ n18707;
  assign n19627 = n18726 & ~n19626;
  assign n19628 = ~n18710 & n19610;
  assign n19629 = ~n19627 & ~n19628;
  assign n19630 = ~n18751 & ~n19629;
  assign n19631 = ~n19624 & ~n19630;
  assign n19632 = ~n19623 & ~n19631;
  assign n19633 = n19620 & n19632;
  assign n19634 = n18746 & n19633;
  assign n19635 = n18741 & n19634;
  assign n19636 = n18717 & n19635;
  assign n19637 = n19636 ^ n17547;
  assign n19638 = n19637 ^ x757;
  assign n19574 = n19108 & n19204;
  assign n19575 = n19171 & n19178;
  assign n19576 = ~n19574 & ~n19575;
  assign n19577 = n19189 & n19218;
  assign n19578 = ~n19176 & ~n19215;
  assign n19579 = n19185 & ~n19578;
  assign n19580 = ~n19577 & ~n19579;
  assign n19581 = n19576 & n19580;
  assign n19582 = n19207 & ~n19218;
  assign n19583 = n19178 & n19193;
  assign n19584 = ~n19582 & ~n19583;
  assign n19585 = n19108 & n19215;
  assign n19586 = ~n19204 & ~n19217;
  assign n19587 = n19169 & ~n19586;
  assign n19588 = ~n19585 & ~n19587;
  assign n19589 = n19108 & n19187;
  assign n19590 = ~n19107 & ~n19223;
  assign n19591 = ~n19589 & ~n19590;
  assign n19592 = n19169 & ~n19182;
  assign n19593 = n19202 & n19218;
  assign n19594 = ~n19202 & ~n19209;
  assign n19595 = ~n19217 & n19594;
  assign n19596 = ~n19189 & n19595;
  assign n19597 = n19185 & ~n19596;
  assign n19598 = ~n19593 & ~n19597;
  assign n19599 = ~n19592 & n19598;
  assign n19600 = n19591 & n19599;
  assign n19601 = n19588 & n19600;
  assign n19602 = n19584 & n19601;
  assign n19603 = n19173 & n19602;
  assign n19604 = n19201 & n19603;
  assign n19605 = n19184 & n19604;
  assign n19606 = n19581 & n19605;
  assign n19607 = n19606 ^ n17525;
  assign n19608 = n19607 ^ x756;
  assign n19639 = n19638 ^ n19608;
  assign n19640 = n18593 ^ x758;
  assign n19641 = n19640 ^ n19608;
  assign n19642 = n19641 ^ n19640;
  assign n19643 = n19104 ^ x755;
  assign n19644 = n19643 ^ n19638;
  assign n19645 = n19644 ^ n19640;
  assign n19646 = n19645 ^ n19640;
  assign n19647 = ~n19642 & ~n19646;
  assign n19648 = n19647 ^ n19640;
  assign n19649 = n19639 & n19648;
  assign n19650 = n19649 ^ n19644;
  assign n19652 = n19651 ^ n19650;
  assign n19653 = n19652 ^ n19650;
  assign n19654 = ~n19638 & ~n19643;
  assign n19655 = ~n19608 & n19654;
  assign n19656 = n19640 ^ n19638;
  assign n19657 = n19656 ^ n19643;
  assign n19658 = n19657 ^ n19656;
  assign n19659 = n19608 & ~n19640;
  assign n19660 = n19638 & n19659;
  assign n19661 = ~n19608 & n19640;
  assign n19662 = ~n19660 & ~n19661;
  assign n19663 = n19662 ^ n19656;
  assign n19664 = ~n19658 & n19663;
  assign n19665 = n19664 ^ n19656;
  assign n19666 = ~n19655 & n19665;
  assign n19667 = n19666 ^ n19650;
  assign n19668 = n19653 & ~n19667;
  assign n19669 = n19668 ^ n19650;
  assign n19670 = ~n19573 & ~n19669;
  assign n19671 = n19608 & n19640;
  assign n19672 = n19654 & n19671;
  assign n19673 = ~n19608 & ~n19640;
  assign n19674 = ~n19643 & n19673;
  assign n19675 = ~n19672 & ~n19674;
  assign n19676 = n19638 & ~n19643;
  assign n19677 = ~n19608 & n19676;
  assign n19678 = n19673 ^ n19643;
  assign n19679 = n19671 ^ n19638;
  assign n19680 = n19679 ^ n19673;
  assign n19681 = ~n19673 & n19680;
  assign n19682 = n19681 ^ n19673;
  assign n19683 = ~n19678 & ~n19682;
  assign n19684 = n19683 ^ n19681;
  assign n19685 = n19684 ^ n19673;
  assign n19686 = n19685 ^ n19679;
  assign n19687 = ~n19671 & n19686;
  assign n19688 = n19687 ^ n19679;
  assign n19689 = ~n19677 & n19688;
  assign n19690 = n19675 & n19689;
  assign n19691 = n19690 ^ n19651;
  assign n19692 = n19691 ^ n19690;
  assign n19693 = n19659 & n19676;
  assign n19694 = n19638 & n19643;
  assign n19695 = ~n19608 & n19694;
  assign n19696 = ~n19693 & ~n19695;
  assign n19697 = n19640 & n19654;
  assign n19698 = ~n19671 & ~n19673;
  assign n19699 = ~n19638 & ~n19698;
  assign n19700 = ~n19697 & ~n19699;
  assign n19701 = n19696 & n19700;
  assign n19702 = n19701 ^ n19690;
  assign n19703 = ~n19692 & n19702;
  assign n19704 = n19703 ^ n19690;
  assign n19705 = n19573 & ~n19704;
  assign n19706 = ~n19670 & ~n19705;
  assign n19707 = n19706 ^ n18216;
  assign n19708 = n19707 ^ x812;
  assign n19709 = ~n18524 & ~n18560;
  assign n19710 = n18518 & ~n19709;
  assign n19711 = n18566 & ~n19710;
  assign n19712 = ~n19434 & n19449;
  assign n19713 = n18458 & ~n19712;
  assign n19714 = n18550 & ~n18553;
  assign n19715 = ~n18527 & n19714;
  assign n19716 = n18518 & ~n19715;
  assign n19717 = ~n19713 & ~n19716;
  assign n19718 = n18521 & n18547;
  assign n19719 = ~n18534 & ~n18548;
  assign n19720 = ~n18544 & ~n18549;
  assign n19721 = ~n18547 & n19720;
  assign n19722 = ~n18512 & n18545;
  assign n19723 = ~n19721 & ~n19722;
  assign n19724 = n19719 & ~n19723;
  assign n19725 = ~n18567 & n19724;
  assign n19726 = ~n18456 & ~n19725;
  assign n19727 = ~n19718 & ~n19726;
  assign n19728 = n19717 & n19727;
  assign n19729 = n19711 & n19728;
  assign n19730 = ~n18591 & n19729;
  assign n19731 = ~n18562 & n19730;
  assign n19732 = n18558 & n19731;
  assign n19733 = n19732 ^ n17011;
  assign n19734 = n19733 ^ x744;
  assign n19735 = n18984 & n19375;
  assign n19736 = n18986 & n19005;
  assign n19737 = ~n19735 & ~n19736;
  assign n19738 = n18993 & n19375;
  assign n19739 = n18947 ^ n18936;
  assign n19740 = n19739 ^ n18937;
  assign n19741 = n19740 ^ n18974;
  assign n19742 = n18937 ^ n18936;
  assign n19743 = n18974 ^ n18936;
  assign n19744 = n19743 ^ n18936;
  assign n19745 = ~n19742 & ~n19744;
  assign n19746 = n19745 ^ n18936;
  assign n19747 = ~n19741 & n19746;
  assign n19748 = ~n18976 & ~n19747;
  assign n19749 = n19010 & n19748;
  assign n19750 = n19005 & ~n19749;
  assign n19751 = ~n18998 & ~n19006;
  assign n19752 = n19371 & n19751;
  assign n19753 = n19017 & ~n19752;
  assign n19754 = n18935 & ~n19024;
  assign n19755 = ~n19753 & ~n19754;
  assign n19756 = ~n18979 & ~n18990;
  assign n19757 = n18933 & ~n19756;
  assign n19758 = ~n19006 & ~n19747;
  assign n19759 = n18987 & ~n19758;
  assign n19760 = ~n19757 & ~n19759;
  assign n19761 = n19755 & n19760;
  assign n19762 = ~n19750 & n19761;
  assign n19763 = ~n19738 & n19762;
  assign n19764 = n18989 & n19763;
  assign n19765 = n19737 & n19764;
  assign n19766 = n19765 ^ n16942;
  assign n19767 = n19766 ^ x745;
  assign n19768 = n18708 & n18730;
  assign n19769 = n18623 & n18742;
  assign n19770 = ~n18715 & n18721;
  assign n19771 = ~n19769 & ~n19770;
  assign n19772 = ~n19768 & n19771;
  assign n19773 = ~n18742 & n18752;
  assign n19774 = n18726 & n19773;
  assign n19775 = n18734 & n19774;
  assign n19776 = n18730 & ~n19775;
  assign n19777 = n18710 & n19614;
  assign n19778 = n18739 & ~n18755;
  assign n19779 = n18721 & ~n19778;
  assign n19780 = ~n19777 & ~n19779;
  assign n19781 = ~n19776 & n19780;
  assign n19782 = n18707 & n18722;
  assign n19783 = n18759 & ~n19782;
  assign n19784 = n18623 & ~n19783;
  assign n19785 = n18714 ^ n18622;
  assign n19787 = n18734 & ~n18748;
  assign n19786 = ~n18744 & n18752;
  assign n19788 = n19787 ^ n19786;
  assign n19789 = n19787 ^ n18595;
  assign n19790 = n19789 ^ n19787;
  assign n19791 = n19788 & ~n19790;
  assign n19792 = n19791 ^ n19787;
  assign n19793 = n19792 ^ n18714;
  assign n19794 = ~n19785 & ~n19793;
  assign n19795 = n19794 ^ n19791;
  assign n19796 = n19795 ^ n19787;
  assign n19797 = n19796 ^ n18622;
  assign n19798 = ~n18714 & n19797;
  assign n19799 = n19798 ^ n18714;
  assign n19800 = n19799 ^ n18622;
  assign n19801 = ~n19784 & n19800;
  assign n19802 = n19781 & n19801;
  assign n19803 = n19772 & n19802;
  assign n19804 = n18729 & n19803;
  assign n19805 = n19804 ^ n16981;
  assign n19806 = n19805 ^ x743;
  assign n19807 = n19767 & n19806;
  assign n19808 = n19235 ^ x746;
  assign n19809 = n19807 & n19808;
  assign n19810 = ~n19734 & n19809;
  assign n19811 = n18930 ^ x747;
  assign n19812 = ~n18375 & n19052;
  assign n19813 = n18382 & ~n19812;
  assign n19814 = ~n18416 & ~n18422;
  assign n19815 = n18399 & ~n19814;
  assign n19816 = ~n18402 & n18423;
  assign n19817 = n18239 & ~n19816;
  assign n19818 = ~n19815 & ~n19817;
  assign n19819 = n18385 & ~n19487;
  assign n19820 = n19481 & ~n19819;
  assign n19821 = ~n18428 & n19820;
  assign n19822 = ~n18396 & n19821;
  assign n19823 = n19041 & ~n19822;
  assign n19824 = n19818 & ~n19823;
  assign n19825 = ~n19037 & n19824;
  assign n19826 = ~n18381 & n19825;
  assign n19827 = ~n19813 & n19826;
  assign n19828 = n18372 ^ n18217;
  assign n19829 = n19828 ^ n18372;
  assign n19830 = n18419 ^ n18372;
  assign n19831 = n19830 ^ n18372;
  assign n19832 = ~n19829 & n19831;
  assign n19833 = n19832 ^ n18372;
  assign n19834 = n18238 & n19833;
  assign n19835 = n19834 ^ n18372;
  assign n19836 = n19827 & ~n19835;
  assign n19837 = n18401 ^ n18399;
  assign n19838 = n19046 ^ n18239;
  assign n19839 = n18401 ^ n18239;
  assign n19840 = n19839 ^ n18239;
  assign n19841 = n19838 & ~n19840;
  assign n19842 = n19841 ^ n18239;
  assign n19843 = n19837 & n19842;
  assign n19844 = n19843 ^ n18399;
  assign n19845 = n19836 & ~n19844;
  assign n19846 = n18409 & n19845;
  assign n19847 = n19846 ^ n17050;
  assign n19848 = n19847 ^ x742;
  assign n19849 = n19811 & n19848;
  assign n19850 = n19810 & n19849;
  assign n19851 = n19734 & ~n19808;
  assign n19852 = n19807 & n19851;
  assign n19853 = n19811 & ~n19848;
  assign n19854 = n19852 & n19853;
  assign n19855 = ~n19850 & ~n19854;
  assign n19856 = ~n19811 & n19848;
  assign n19857 = n19852 & n19856;
  assign n19858 = n19734 & n19809;
  assign n19859 = n19853 & n19858;
  assign n19860 = ~n19857 & ~n19859;
  assign n19861 = n19767 & ~n19806;
  assign n19862 = ~n19767 & n19808;
  assign n19863 = n19734 & n19862;
  assign n19864 = n19806 & n19863;
  assign n19865 = ~n19861 & ~n19864;
  assign n19866 = n19856 & ~n19865;
  assign n19867 = ~n19767 & n19851;
  assign n19868 = n19806 & n19867;
  assign n19869 = ~n19810 & ~n19868;
  assign n19870 = n19853 & ~n19869;
  assign n19871 = ~n19806 & n19863;
  assign n19872 = ~n19734 & ~n19808;
  assign n19873 = ~n19767 & n19872;
  assign n19874 = ~n19806 & n19873;
  assign n19875 = ~n19871 & ~n19874;
  assign n19876 = ~n19856 & ~n19875;
  assign n19877 = ~n19734 & n19862;
  assign n19878 = n19806 & n19877;
  assign n19879 = ~n19868 & ~n19878;
  assign n19880 = n19848 & ~n19879;
  assign n19881 = ~n19876 & ~n19880;
  assign n19882 = ~n19806 & n19877;
  assign n19883 = n19851 & n19861;
  assign n19884 = ~n19852 & ~n19883;
  assign n19885 = ~n19882 & n19884;
  assign n19886 = n19849 & ~n19885;
  assign n19887 = ~n19811 & ~n19848;
  assign n19888 = n19806 & n19873;
  assign n19889 = n19808 & n19861;
  assign n19890 = ~n19734 & n19889;
  assign n19891 = ~n19806 & n19867;
  assign n19892 = ~n19890 & ~n19891;
  assign n19893 = ~n19888 & n19892;
  assign n19894 = ~n19810 & n19893;
  assign n19895 = n19887 & ~n19894;
  assign n19896 = ~n19886 & ~n19895;
  assign n19897 = n19881 & n19896;
  assign n19898 = ~n19870 & n19897;
  assign n19899 = ~n19866 & n19898;
  assign n19900 = n19807 & n19872;
  assign n19901 = ~n19864 & ~n19900;
  assign n19902 = n19901 ^ n19811;
  assign n19903 = n19902 ^ n19901;
  assign n19904 = n19861 & n19872;
  assign n19905 = ~n19882 & ~n19904;
  assign n19906 = n19905 ^ n19901;
  assign n19907 = n19903 & n19906;
  assign n19908 = n19907 ^ n19901;
  assign n19909 = ~n19848 & ~n19908;
  assign n19910 = n19899 & ~n19909;
  assign n19911 = n19860 & n19910;
  assign n19912 = n19855 & n19911;
  assign n19913 = n19912 ^ n19134;
  assign n19914 = n19913 ^ x810;
  assign n19915 = ~n19708 & ~n19914;
  assign n19916 = n17493 ^ x766;
  assign n19917 = n19185 & n19204;
  assign n19918 = n19187 ^ n19106;
  assign n19919 = n19918 ^ n19187;
  assign n19920 = n19207 ^ n19187;
  assign n19921 = n19920 ^ n19187;
  assign n19922 = ~n19919 & n19921;
  assign n19923 = n19922 ^ n19187;
  assign n19924 = ~n19107 & n19923;
  assign n19925 = n19924 ^ n19187;
  assign n19926 = ~n19917 & ~n19925;
  assign n19927 = n19218 & ~n19578;
  assign n19928 = n19185 & ~n19211;
  assign n19929 = ~n19927 & ~n19928;
  assign n19930 = n19178 & n19180;
  assign n19931 = n19169 & ~n19594;
  assign n19932 = ~n19222 & n19594;
  assign n19933 = ~n19217 & n19932;
  assign n19934 = n19108 & ~n19933;
  assign n19935 = ~n19931 & ~n19934;
  assign n19936 = ~n19930 & n19935;
  assign n19937 = n19929 & n19936;
  assign n19938 = n19588 & n19937;
  assign n19939 = n19584 & n19938;
  assign n19940 = n19926 & n19939;
  assign n19941 = n19192 & n19940;
  assign n19942 = n19174 & n19941;
  assign n19943 = n19942 ^ n17241;
  assign n19944 = n19943 ^ x771;
  assign n19945 = ~n19916 & ~n19944;
  assign n19946 = n18977 & n18991;
  assign n19947 = ~n18990 & ~n19946;
  assign n19948 = ~n18993 & n19947;
  assign n19949 = n19005 & ~n19948;
  assign n19950 = ~n19008 & n19375;
  assign n19951 = ~n19949 & ~n19950;
  assign n19952 = n18997 & ~n19370;
  assign n19953 = n18987 & ~n19952;
  assign n19954 = n18935 & n18993;
  assign n19955 = ~n18979 & n19010;
  assign n19956 = ~n18986 & n19955;
  assign n19957 = n18935 & n18983;
  assign n19958 = ~n19375 & ~n19957;
  assign n19959 = ~n19956 & ~n19958;
  assign n19960 = ~n18976 & n19948;
  assign n19961 = n18987 & ~n19960;
  assign n19962 = ~n18996 & n19000;
  assign n19963 = ~n19006 & n19962;
  assign n19964 = n19005 & ~n19963;
  assign n19965 = ~n19961 & ~n19964;
  assign n19966 = ~n19959 & n19965;
  assign n19967 = ~n19954 & n19966;
  assign n19968 = ~n18981 & n19967;
  assign n19969 = ~n19953 & n19968;
  assign n19970 = n19018 ^ n18935;
  assign n19971 = ~n18986 & n19751;
  assign n19972 = n19971 ^ n18933;
  assign n19973 = n18935 ^ n18933;
  assign n19974 = n19973 ^ n18933;
  assign n19975 = n19972 & n19974;
  assign n19976 = n19975 ^ n18933;
  assign n19977 = n19970 & ~n19976;
  assign n19978 = n19977 ^ n19018;
  assign n19979 = n19969 & ~n19978;
  assign n19980 = n19951 & n19979;
  assign n19981 = n19737 & n19980;
  assign n19982 = n19981 ^ n17669;
  assign n19983 = n19982 ^ x768;
  assign n19984 = n17900 & n17905;
  assign n19985 = ~n17903 & n19401;
  assign n19986 = ~n17923 & n19985;
  assign n19987 = n17884 & ~n19986;
  assign n19988 = ~n19984 & ~n19987;
  assign n19989 = n17880 & n17929;
  assign n19990 = ~n17923 & n19410;
  assign n19991 = n17882 & ~n19990;
  assign n19992 = n17897 ^ n17879;
  assign n19994 = ~n17917 & n19399;
  assign n19993 = n18898 & n19401;
  assign n19995 = n19994 ^ n19993;
  assign n19996 = n19994 ^ n17840;
  assign n19997 = n19996 ^ n19994;
  assign n19998 = n19995 & n19997;
  assign n19999 = n19998 ^ n19994;
  assign n20000 = n19999 ^ n17897;
  assign n20001 = n19992 & ~n20000;
  assign n20002 = n20001 ^ n19998;
  assign n20003 = n20002 ^ n19994;
  assign n20004 = n20003 ^ n17879;
  assign n20005 = ~n17897 & ~n20004;
  assign n20006 = n20005 ^ n17897;
  assign n20007 = n20006 ^ n17879;
  assign n20008 = ~n19991 & ~n20007;
  assign n20009 = ~n19989 & n20008;
  assign n20010 = n19988 & n20009;
  assign n20011 = n19398 & n20010;
  assign n20012 = n19395 & n20011;
  assign n20013 = n17896 & n20012;
  assign n20014 = n18900 & n20013;
  assign n20015 = n20014 ^ n17697;
  assign n20016 = n20015 ^ x769;
  assign n20017 = n19983 & ~n20016;
  assign n20018 = ~n18456 & n18510;
  assign n20019 = ~n18538 & n19719;
  assign n20020 = n18518 & ~n20019;
  assign n20021 = ~n18527 & ~n18534;
  assign n20022 = n18547 & ~n20021;
  assign n20023 = ~n18536 & n18568;
  assign n20024 = ~n18548 & n20023;
  assign n20025 = n18512 & ~n20024;
  assign n20026 = ~n20022 & ~n20025;
  assign n20027 = ~n20020 & n20026;
  assign n20028 = ~n20018 & n20027;
  assign n20029 = ~n18515 & ~n18538;
  assign n20030 = ~n18544 & n20029;
  assign n20031 = n18547 & ~n20030;
  assign n20032 = ~n18547 & n18550;
  assign n20033 = n18528 & n20032;
  assign n20034 = ~n18556 & n20033;
  assign n20035 = n18458 & ~n20034;
  assign n20036 = ~n20031 & ~n20035;
  assign n20037 = n20028 & n20036;
  assign n20038 = ~n18554 & n20037;
  assign n20039 = n18517 & n20038;
  assign n20040 = ~n19469 & n20039;
  assign n20041 = n19711 & n20040;
  assign n20042 = ~n18563 & n20041;
  assign n20043 = ~n18562 & n20042;
  assign n20044 = n20043 ^ n17160;
  assign n20045 = n20044 ^ x770;
  assign n20046 = n18781 ^ x767;
  assign n20047 = ~n20045 & ~n20046;
  assign n20048 = n20017 & n20047;
  assign n20049 = n19945 & n20048;
  assign n20050 = n19916 & ~n19944;
  assign n20051 = ~n19983 & ~n20016;
  assign n20052 = n20047 & n20051;
  assign n20053 = n20045 & ~n20046;
  assign n20054 = n20017 & n20053;
  assign n20055 = ~n20052 & ~n20054;
  assign n20056 = n20050 & ~n20055;
  assign n20057 = ~n20049 & ~n20056;
  assign n20058 = n19916 & n19944;
  assign n20059 = n19983 & n20016;
  assign n20060 = ~n20045 & n20046;
  assign n20061 = n20059 & n20060;
  assign n20062 = n20045 & n20046;
  assign n20063 = n20051 & n20062;
  assign n20064 = ~n19983 & n20016;
  assign n20065 = n20060 & n20064;
  assign n20066 = ~n20063 & ~n20065;
  assign n20067 = ~n20061 & n20066;
  assign n20068 = n20058 & ~n20067;
  assign n20069 = n20053 & n20059;
  assign n20070 = n20050 & n20069;
  assign n20071 = n20053 & n20064;
  assign n20072 = ~n20052 & ~n20071;
  assign n20073 = n20047 & n20064;
  assign n20074 = ~n20054 & ~n20073;
  assign n20075 = n20072 & n20074;
  assign n20076 = n20058 & ~n20075;
  assign n20077 = ~n19916 & n19944;
  assign n20078 = n20051 & n20053;
  assign n20079 = ~n20073 & ~n20078;
  assign n20080 = n20055 & n20079;
  assign n20081 = n20077 & ~n20080;
  assign n20082 = ~n20076 & ~n20081;
  assign n20083 = n19944 ^ n19916;
  assign n20086 = n20062 & n20064;
  assign n20090 = n20067 & ~n20086;
  assign n20084 = n20059 & n20062;
  assign n20085 = n20017 & n20060;
  assign n20087 = ~n20061 & ~n20086;
  assign n20088 = ~n20085 & n20087;
  assign n20089 = ~n20084 & n20088;
  assign n20091 = n20090 ^ n20089;
  assign n20092 = n20090 ^ n19944;
  assign n20093 = n20092 ^ n20090;
  assign n20094 = n20091 & n20093;
  assign n20095 = n20094 ^ n20090;
  assign n20096 = n20083 & ~n20095;
  assign n20097 = n20082 & ~n20096;
  assign n20105 = n20017 & n20062;
  assign n20098 = n20051 & n20060;
  assign n20099 = n20047 & n20059;
  assign n20100 = ~n20069 & ~n20099;
  assign n20101 = ~n20085 & n20100;
  assign n20102 = n20066 & n20101;
  assign n20103 = ~n20071 & n20102;
  assign n20104 = ~n20098 & n20103;
  assign n20106 = n20105 ^ n20104;
  assign n20107 = n20106 ^ n20105;
  assign n20108 = n20105 ^ n19944;
  assign n20109 = n20108 ^ n20105;
  assign n20110 = ~n20107 & ~n20109;
  assign n20111 = n20110 ^ n20105;
  assign n20112 = ~n19916 & n20111;
  assign n20113 = n20112 ^ n20105;
  assign n20114 = n20097 & ~n20113;
  assign n20115 = ~n20070 & n20114;
  assign n20116 = ~n20068 & n20115;
  assign n20117 = n20057 & n20116;
  assign n20118 = n20117 ^ n19157;
  assign n20119 = n20118 ^ x811;
  assign n20120 = n19390 ^ x736;
  assign n20121 = n19805 ^ x741;
  assign n20122 = n20120 & n20121;
  assign n20123 = n18108 & n18166;
  assign n20124 = n18119 & n18141;
  assign n20125 = ~n20123 & ~n20124;
  assign n20126 = n18110 & ~n18153;
  assign n20127 = n18028 ^ n17986;
  assign n20128 = n20127 ^ n17987;
  assign n20129 = n20128 ^ n18073;
  assign n20130 = n18073 ^ n17987;
  assign n20131 = n20130 ^ n17987;
  assign n20132 = n17987 ^ n17986;
  assign n20133 = n20132 ^ n17987;
  assign n20134 = ~n20131 & ~n20133;
  assign n20135 = n20134 ^ n17987;
  assign n20136 = n20129 & ~n20135;
  assign n20137 = n18123 & n20136;
  assign n20138 = ~n18135 & ~n18147;
  assign n20139 = ~n18166 & n20138;
  assign n20140 = ~n19087 & ~n20139;
  assign n20141 = ~n20137 & ~n20140;
  assign n20142 = ~n20126 & n20141;
  assign n20143 = n20125 & n20142;
  assign n20144 = n19085 & n20143;
  assign n20145 = n19082 & n20144;
  assign n20146 = n18145 & n20145;
  assign n20147 = n19337 & n20146;
  assign n20148 = n18129 & n20147;
  assign n20149 = n18118 & n20148;
  assign n20150 = n20149 ^ n17369;
  assign n20151 = n20150 ^ x738;
  assign n20152 = n19182 & n19223;
  assign n20153 = n19108 & ~n20152;
  assign n20154 = ~n19221 & n19595;
  assign n20155 = n19178 & ~n20154;
  assign n20156 = ~n20153 & ~n20155;
  assign n20157 = n19215 ^ n19106;
  assign n20158 = n20157 ^ n19215;
  assign n20159 = ~n19181 & n19932;
  assign n20160 = ~n19171 & n20159;
  assign n20161 = n20160 ^ n19215;
  assign n20162 = n20161 ^ n19215;
  assign n20163 = n20158 & ~n20162;
  assign n20164 = n20163 ^ n19215;
  assign n20165 = n19107 & n20164;
  assign n20166 = n20165 ^ n19215;
  assign n20167 = n20156 & ~n20166;
  assign n20168 = n19217 ^ n19185;
  assign n20169 = n19217 ^ n19108;
  assign n20170 = n20169 ^ n19108;
  assign n20171 = ~n19158 & n19162;
  assign n20172 = n20171 ^ n19108;
  assign n20173 = ~n20170 & ~n20172;
  assign n20174 = n20173 ^ n19108;
  assign n20175 = n20168 & n20174;
  assign n20176 = n20175 ^ n19185;
  assign n20177 = n20167 & ~n20176;
  assign n20178 = n19926 & n20177;
  assign n20179 = n19198 & n20178;
  assign n20180 = n19581 & n20179;
  assign n20181 = n20180 ^ n17338;
  assign n20182 = n20181 ^ x739;
  assign n20183 = ~n20151 & n20182;
  assign n20184 = n19331 ^ x737;
  assign n20185 = n19847 ^ x740;
  assign n20186 = n20184 & n20185;
  assign n20187 = n20183 & n20186;
  assign n20188 = n20122 & n20187;
  assign n20189 = ~n20151 & ~n20182;
  assign n20190 = n20184 & ~n20185;
  assign n20191 = n20189 & n20190;
  assign n20192 = n20122 & n20191;
  assign n20193 = ~n20188 & ~n20192;
  assign n20194 = ~n20120 & n20121;
  assign n20195 = n20151 & ~n20182;
  assign n20196 = ~n20184 & n20185;
  assign n20197 = n20195 & n20196;
  assign n20198 = n20194 & n20197;
  assign n20199 = n20151 & n20182;
  assign n20200 = n20196 & n20199;
  assign n20201 = ~n20184 & ~n20185;
  assign n20202 = n20189 & n20201;
  assign n20203 = ~n20200 & ~n20202;
  assign n20204 = n20122 & ~n20203;
  assign n20205 = ~n20198 & ~n20204;
  assign n20206 = ~n20120 & ~n20121;
  assign n20207 = n20189 & n20196;
  assign n20208 = n20195 & n20201;
  assign n20209 = ~n20207 & ~n20208;
  assign n20210 = n20206 & ~n20209;
  assign n20211 = n20120 & ~n20121;
  assign n20212 = n20183 & n20196;
  assign n20213 = n20211 & n20212;
  assign n20214 = n20120 & n20208;
  assign n20215 = ~n20213 & ~n20214;
  assign n20216 = n20122 & n20199;
  assign n20217 = n20186 & n20216;
  assign n20218 = n20190 & n20216;
  assign n20219 = n20184 ^ n20182;
  assign n20220 = n20219 ^ n20185;
  assign n20221 = n20220 ^ n20182;
  assign n20222 = n20221 ^ n20220;
  assign n20223 = n20220 ^ n20185;
  assign n20224 = n20222 & ~n20223;
  assign n20225 = n20224 ^ n20220;
  assign n20226 = ~n20151 & n20225;
  assign n20227 = n20226 ^ n20220;
  assign n20228 = n20206 & n20227;
  assign n20229 = ~n20218 & ~n20228;
  assign n20230 = ~n20197 & ~n20207;
  assign n20231 = n20184 & n20199;
  assign n20232 = n20186 & n20195;
  assign n20233 = ~n20231 & ~n20232;
  assign n20234 = ~n20191 & n20233;
  assign n20235 = n20230 & n20234;
  assign n20236 = n20211 & ~n20235;
  assign n20237 = n20122 & n20207;
  assign n20238 = n20183 & n20201;
  assign n20239 = ~n20200 & ~n20238;
  assign n20240 = n20183 & n20190;
  assign n20241 = n20186 & n20189;
  assign n20242 = n20190 & n20195;
  assign n20243 = n20190 & n20199;
  assign n20244 = ~n20242 & ~n20243;
  assign n20245 = ~n20241 & n20244;
  assign n20246 = ~n20240 & n20245;
  assign n20247 = n20239 & n20246;
  assign n20248 = ~n20232 & n20247;
  assign n20249 = n20194 & ~n20248;
  assign n20250 = ~n20237 & ~n20249;
  assign n20251 = ~n20236 & n20250;
  assign n20252 = n20229 & n20251;
  assign n20253 = ~n20217 & n20252;
  assign n20254 = n20215 & n20253;
  assign n20255 = ~n20210 & n20254;
  assign n20256 = n20205 & n20255;
  assign n20257 = n20193 & n20256;
  assign n20258 = n20257 ^ n17444;
  assign n20259 = n20258 ^ x809;
  assign n20260 = n20119 & n20259;
  assign n20261 = n19915 & n20260;
  assign n20262 = n19572 & n20261;
  assign n20263 = n19318 & ~n19571;
  assign n20264 = ~n20119 & n20259;
  assign n20265 = n19915 & n20264;
  assign n20266 = n19708 & n19914;
  assign n20267 = ~n20119 & ~n20259;
  assign n20268 = n20266 & n20267;
  assign n20269 = ~n20265 & ~n20268;
  assign n20270 = n20263 & ~n20269;
  assign n20271 = ~n20262 & ~n20270;
  assign n20272 = ~n19708 & n19914;
  assign n20273 = n20119 & ~n20259;
  assign n20274 = n20272 & n20273;
  assign n20275 = n19572 & n20274;
  assign n20276 = ~n19318 & ~n19571;
  assign n20277 = n20265 & n20276;
  assign n20278 = n19571 ^ n19318;
  assign n20279 = n19708 & ~n19914;
  assign n20280 = n20267 & n20279;
  assign n20281 = ~n20278 & n20280;
  assign n20282 = ~n20277 & ~n20281;
  assign n20283 = n20260 & n20266;
  assign n20284 = n20264 & n20272;
  assign n20285 = ~n20283 & ~n20284;
  assign n20286 = n20276 & ~n20285;
  assign n20287 = n20282 & ~n20286;
  assign n20288 = n20263 & n20283;
  assign n20289 = n19915 & n20267;
  assign n20290 = n19572 & n20289;
  assign n20291 = ~n20288 & ~n20290;
  assign n20292 = n20264 & n20266;
  assign n20293 = n19572 & n20292;
  assign n20294 = n19318 & n19571;
  assign n20295 = n20289 & n20294;
  assign n20296 = ~n20293 & ~n20295;
  assign n20297 = n20264 & n20279;
  assign n20298 = n20294 & n20297;
  assign n20299 = n19572 & n20280;
  assign n20300 = ~n20298 & ~n20299;
  assign n20301 = n20268 & ~n20278;
  assign n20302 = n20274 & n20276;
  assign n20303 = ~n20301 & ~n20302;
  assign n20304 = n20260 & n20279;
  assign n20305 = n20260 & n20272;
  assign n20306 = ~n20304 & ~n20305;
  assign n20307 = n19572 & ~n20306;
  assign n20308 = n20266 & n20273;
  assign n20309 = n19915 & n20273;
  assign n20310 = ~n20308 & ~n20309;
  assign n20311 = ~n20284 & n20310;
  assign n20312 = ~n20304 & n20311;
  assign n20313 = n20294 & ~n20312;
  assign n20314 = n20273 & n20279;
  assign n20315 = n20267 & n20272;
  assign n20316 = ~n20314 & ~n20315;
  assign n20317 = ~n20308 & n20316;
  assign n20318 = ~n20297 & n20317;
  assign n20319 = ~n20261 & n20318;
  assign n20320 = n20263 & ~n20319;
  assign n20321 = ~n20313 & ~n20320;
  assign n20322 = ~n20307 & n20321;
  assign n20323 = n20303 & n20322;
  assign n20324 = n20300 & n20323;
  assign n20325 = n20296 & n20324;
  assign n20326 = n20291 & n20325;
  assign n20327 = n20314 ^ n19571;
  assign n20328 = n20327 ^ n20314;
  assign n20329 = n20314 ^ n20306;
  assign n20330 = ~n20328 & ~n20329;
  assign n20331 = n20330 ^ n20314;
  assign n20332 = ~n19318 & n20331;
  assign n20333 = n20326 & ~n20332;
  assign n20334 = n20287 & n20333;
  assign n20335 = ~n20275 & n20334;
  assign n20336 = n20271 & n20335;
  assign n20337 = n20336 ^ n19235;
  assign n20338 = n19734 & n19889;
  assign n20339 = ~n19904 & ~n20338;
  assign n20340 = n19856 & ~n20339;
  assign n20341 = n19849 & n19891;
  assign n20342 = n19853 & n19888;
  assign n20343 = ~n20341 & ~n20342;
  assign n20344 = ~n20340 & n20343;
  assign n20345 = n19883 & n19887;
  assign n20346 = ~n19874 & ~n19890;
  assign n20347 = ~n19882 & n20346;
  assign n20348 = ~n19849 & ~n19887;
  assign n20349 = ~n20347 & ~n20348;
  assign n20350 = ~n19852 & n19901;
  assign n20351 = ~n19878 & n20350;
  assign n20352 = n19887 & ~n20351;
  assign n20353 = n19808 ^ n19806;
  assign n20354 = n19767 ^ n19734;
  assign n20355 = n20354 ^ n19808;
  assign n20356 = n20355 ^ n20354;
  assign n20357 = n20354 ^ n19734;
  assign n20358 = n20357 ^ n20354;
  assign n20359 = n20356 & n20358;
  assign n20360 = n20359 ^ n20354;
  assign n20361 = n20353 & n20360;
  assign n20362 = n20361 ^ n20354;
  assign n20363 = n19853 & n20362;
  assign n20364 = ~n20352 & ~n20363;
  assign n20365 = n19856 & ~n19875;
  assign n20366 = ~n19856 & n20350;
  assign n20367 = ~n19849 & ~n19900;
  assign n20368 = n19879 & n20367;
  assign n20369 = ~n19858 & n20368;
  assign n20370 = ~n20366 & ~n20369;
  assign n20371 = n19848 & n20370;
  assign n20372 = ~n20365 & ~n20371;
  assign n20373 = n20364 & n20372;
  assign n20374 = n19855 & n20373;
  assign n20375 = ~n20349 & n20374;
  assign n20376 = ~n20345 & n20375;
  assign n20377 = n20344 & n20376;
  assign n20378 = n20377 ^ n17123;
  assign n20379 = n20378 ^ x801;
  assign n20380 = n18858 ^ x796;
  assign n20381 = ~n20379 & n20380;
  assign n20382 = n17448 & n17473;
  assign n20383 = ~n17133 & n17475;
  assign n20384 = ~n20382 & ~n20383;
  assign n20385 = ~n17461 & n17464;
  assign n20386 = n17446 & ~n17489;
  assign n20387 = ~n20385 & ~n20386;
  assign n20388 = n20384 & n20387;
  assign n20389 = n20388 ^ n17174;
  assign n20390 = n20389 ^ x774;
  assign n20391 = n19367 ^ x776;
  assign n20392 = n20390 & ~n20391;
  assign n20393 = ~n18725 & n18753;
  assign n20394 = n18734 & n20393;
  assign n20395 = n18623 & ~n20394;
  assign n20396 = ~n18719 & n18726;
  assign n20397 = ~n18748 & n20396;
  assign n20398 = n18721 & ~n20397;
  assign n20399 = n18733 & ~n19624;
  assign n20400 = n18707 & n18732;
  assign n20401 = ~n18737 & ~n20400;
  assign n20402 = n18727 & n20401;
  assign n20403 = n18710 & ~n20402;
  assign n20404 = n18739 & ~n18744;
  assign n20405 = n18759 & n20404;
  assign n20406 = n18730 & ~n20405;
  assign n20407 = ~n20403 & ~n20406;
  assign n20408 = ~n20399 & n20407;
  assign n20409 = ~n20398 & n20408;
  assign n20410 = ~n20395 & n20409;
  assign n20411 = ~n18776 & n20410;
  assign n20412 = n19772 & n20411;
  assign n20413 = n18717 & n20412;
  assign n20414 = n20413 ^ n17204;
  assign n20415 = n20414 ^ x775;
  assign n20416 = n19943 ^ x773;
  assign n20417 = n20415 & ~n20416;
  assign n20418 = n20392 & n20417;
  assign n20419 = n20044 ^ x772;
  assign n20420 = n19500 ^ x777;
  assign n20421 = ~n20419 & n20420;
  assign n20422 = ~n20419 & ~n20420;
  assign n20423 = ~n20421 & ~n20422;
  assign n20424 = n20418 & ~n20423;
  assign n20425 = n20419 & n20420;
  assign n20426 = ~n20390 & n20391;
  assign n20427 = ~n20415 & n20416;
  assign n20428 = n20426 & n20427;
  assign n20429 = ~n20390 & ~n20391;
  assign n20430 = n20415 & n20416;
  assign n20431 = n20429 & n20430;
  assign n20432 = ~n20428 & ~n20431;
  assign n20433 = n20425 & ~n20432;
  assign n20434 = ~n20424 & ~n20433;
  assign n20435 = n20417 & n20429;
  assign n20436 = n20421 & n20435;
  assign n20437 = ~n20422 & ~n20425;
  assign n20438 = n20392 & ~n20437;
  assign n20439 = n20427 & n20438;
  assign n20440 = ~n20436 & ~n20439;
  assign n20441 = n20392 & n20430;
  assign n20442 = n20425 & n20441;
  assign n20443 = n20427 & n20429;
  assign n20444 = n20421 & n20443;
  assign n20445 = ~n20442 & ~n20444;
  assign n20446 = n20390 & n20391;
  assign n20447 = n20417 & n20446;
  assign n20448 = ~n20415 & ~n20416;
  assign n20449 = n20446 & n20448;
  assign n20450 = n20429 & n20448;
  assign n20451 = ~n20449 & ~n20450;
  assign n20452 = ~n20447 & n20451;
  assign n20453 = n20425 & ~n20452;
  assign n20454 = n20426 & n20448;
  assign n20455 = ~n20419 & n20454;
  assign n20456 = n20427 & n20446;
  assign n20457 = ~n20431 & ~n20456;
  assign n20458 = ~n20449 & n20457;
  assign n20459 = n20421 & ~n20458;
  assign n20460 = ~n20455 & ~n20459;
  assign n20461 = ~n20453 & n20460;
  assign n20462 = n20419 & ~n20420;
  assign n20463 = n20417 & n20426;
  assign n20464 = ~n20450 & ~n20463;
  assign n20465 = ~n20456 & n20464;
  assign n20466 = n20415 ^ n20391;
  assign n20467 = n20415 ^ n20390;
  assign n20468 = n20467 ^ n20416;
  assign n20469 = n20466 & n20468;
  assign n20470 = n20465 & ~n20469;
  assign n20471 = ~n20447 & n20470;
  assign n20472 = n20462 & n20471;
  assign n20473 = n20426 & n20430;
  assign n20474 = ~n20469 & ~n20473;
  assign n20475 = n20422 & ~n20474;
  assign n20476 = ~n20472 & ~n20475;
  assign n20477 = n20461 & n20476;
  assign n20478 = n20435 ^ n20419;
  assign n20479 = n20478 ^ n20435;
  assign n20480 = n20463 ^ n20435;
  assign n20481 = ~n20479 & n20480;
  assign n20482 = n20481 ^ n20435;
  assign n20483 = n20420 & n20482;
  assign n20484 = n20477 & ~n20483;
  assign n20485 = n20445 & n20484;
  assign n20486 = n20440 & n20485;
  assign n20487 = n20434 & n20486;
  assign n20488 = n20487 ^ n17300;
  assign n20489 = n20488 ^ x800;
  assign n20490 = n19945 & n20086;
  assign n20491 = ~n20061 & ~n20063;
  assign n20492 = n20050 & ~n20491;
  assign n20493 = ~n20490 & ~n20492;
  assign n20494 = ~n20065 & ~n20084;
  assign n20495 = n19945 & ~n20494;
  assign n20496 = ~n19916 & n20085;
  assign n20497 = ~n20050 & ~n20077;
  assign n20498 = n20098 & ~n20497;
  assign n20499 = ~n20496 & ~n20498;
  assign n20500 = n20050 & n20086;
  assign n20501 = ~n20084 & ~n20105;
  assign n20502 = n20077 & ~n20501;
  assign n20503 = ~n20048 & n20066;
  assign n20504 = ~n20069 & ~n20085;
  assign n20505 = n20503 & n20504;
  assign n20506 = n20055 & n20505;
  assign n20507 = ~n20084 & n20506;
  assign n20508 = n20058 & ~n20507;
  assign n20509 = n20079 & n20100;
  assign n20510 = n20050 & ~n20509;
  assign n20511 = n19945 & ~n20072;
  assign n20512 = ~n20071 & ~n20073;
  assign n20513 = n20077 & ~n20512;
  assign n20514 = ~n20511 & ~n20513;
  assign n20515 = ~n20099 & n20514;
  assign n20516 = ~n20054 & n20515;
  assign n20517 = ~n19916 & ~n20516;
  assign n20518 = ~n20510 & ~n20517;
  assign n20519 = ~n20508 & n20518;
  assign n20520 = ~n20502 & n20519;
  assign n20521 = ~n20500 & n20520;
  assign n20522 = n20499 & n20521;
  assign n20523 = ~n20495 & n20522;
  assign n20524 = n20493 & n20523;
  assign n20525 = n20524 ^ n18506;
  assign n20526 = n20525 ^ x799;
  assign n20527 = n20489 & n20526;
  assign n20528 = n19573 & n19651;
  assign n20529 = n19643 ^ n19640;
  assign n20530 = n20529 ^ n19608;
  assign n20531 = n19642 & ~n19656;
  assign n20532 = n20531 ^ n19640;
  assign n20533 = ~n20530 & ~n20532;
  assign n20534 = n20533 ^ n19640;
  assign n20535 = n20528 & ~n20534;
  assign n20536 = ~n19573 & n19651;
  assign n20537 = n19643 & ~n19662;
  assign n20538 = n19654 ^ n19608;
  assign n20539 = n20538 ^ n19654;
  assign n20540 = n19656 ^ n19654;
  assign n20541 = ~n20539 & ~n20540;
  assign n20542 = n20541 ^ n19654;
  assign n20543 = ~n20537 & ~n20542;
  assign n20544 = n20536 & n20543;
  assign n20545 = ~n20535 & ~n20544;
  assign n20546 = n19644 & n19661;
  assign n20547 = n19573 & n20546;
  assign n20548 = n19573 & ~n19651;
  assign n20549 = n19643 & n19656;
  assign n20550 = n19675 & ~n20549;
  assign n20551 = n20548 & ~n20550;
  assign n20552 = ~n20547 & ~n20551;
  assign n20553 = ~n19573 & ~n19651;
  assign n20554 = ~n19640 & n19654;
  assign n20555 = n19671 & n19676;
  assign n20556 = ~n20554 & ~n20555;
  assign n20557 = ~n19638 & n19673;
  assign n20558 = n19694 & n19698;
  assign n20559 = ~n20557 & ~n20558;
  assign n20560 = n20556 & n20559;
  assign n20561 = n19675 & n20560;
  assign n20562 = n20553 & ~n20561;
  assign n20563 = n20552 & ~n20562;
  assign n20564 = n20545 & n20563;
  assign n20565 = n20564 ^ n18471;
  assign n20566 = n20565 ^ x798;
  assign n20567 = n20122 & n20240;
  assign n20568 = ~n20207 & ~n20238;
  assign n20569 = n20194 & ~n20568;
  assign n20570 = ~n20217 & ~n20569;
  assign n20571 = n20206 & n20240;
  assign n20572 = ~n20198 & ~n20571;
  assign n20573 = n20122 & ~n20230;
  assign n20574 = n20211 & ~n20239;
  assign n20575 = ~n20573 & ~n20574;
  assign n20576 = n20201 & n20216;
  assign n20577 = n20199 & n20201;
  assign n20578 = ~n20212 & ~n20577;
  assign n20579 = ~n20207 & n20578;
  assign n20580 = n20206 & ~n20579;
  assign n20581 = ~n20576 & ~n20580;
  assign n20582 = n20186 & n20199;
  assign n20583 = ~n20187 & ~n20582;
  assign n20584 = n20203 & n20583;
  assign n20585 = n20194 & ~n20584;
  assign n20586 = ~n20192 & ~n20242;
  assign n20587 = ~n20211 & n20586;
  assign n20588 = ~n20206 & n20587;
  assign n20589 = ~n20122 & ~n20206;
  assign n20590 = ~n20241 & n20589;
  assign n20591 = ~n20191 & ~n20211;
  assign n20592 = ~n20590 & ~n20591;
  assign n20593 = n20244 & ~n20592;
  assign n20594 = ~n20232 & n20593;
  assign n20595 = ~n20588 & ~n20594;
  assign n20596 = ~n20585 & ~n20595;
  assign n20597 = n20581 & n20596;
  assign n20598 = n20575 & n20597;
  assign n20599 = n20572 & n20598;
  assign n20600 = n20215 & n20599;
  assign n20601 = n20570 & n20600;
  assign n20602 = ~n20567 & n20601;
  assign n20603 = n20602 ^ n18106;
  assign n20604 = n20603 ^ x797;
  assign n20605 = n20566 & n20604;
  assign n20606 = n20527 & n20605;
  assign n20607 = n20381 & n20606;
  assign n20608 = n20379 & ~n20380;
  assign n20609 = n20489 & ~n20526;
  assign n20610 = ~n20566 & ~n20604;
  assign n20611 = n20609 & n20610;
  assign n20612 = n20608 & n20611;
  assign n20613 = ~n20607 & ~n20612;
  assign n20614 = ~n20381 & ~n20608;
  assign n20615 = n20605 & n20609;
  assign n20616 = n20614 & n20615;
  assign n20617 = ~n20379 & ~n20380;
  assign n20618 = n20566 & ~n20604;
  assign n20619 = n20527 & n20618;
  assign n20620 = ~n20489 & ~n20526;
  assign n20621 = n20618 & n20620;
  assign n20622 = ~n20619 & ~n20621;
  assign n20623 = n20617 & ~n20622;
  assign n20624 = ~n20616 & ~n20623;
  assign n20625 = n20613 & n20624;
  assign n20626 = ~n20489 & n20526;
  assign n20627 = ~n20566 & n20604;
  assign n20628 = n20626 & n20627;
  assign n20629 = n20618 & n20626;
  assign n20630 = ~n20628 & ~n20629;
  assign n20631 = ~n20380 & ~n20630;
  assign n20632 = n20527 & n20627;
  assign n20633 = n20527 & n20610;
  assign n20634 = ~n20632 & ~n20633;
  assign n20635 = n20617 & ~n20634;
  assign n20636 = ~n20631 & ~n20635;
  assign n20637 = ~n20606 & ~n20628;
  assign n20638 = n20637 ^ n20380;
  assign n20639 = n20638 ^ n20637;
  assign n20640 = n20609 & n20618;
  assign n20641 = n20610 & n20620;
  assign n20642 = ~n20640 & ~n20641;
  assign n20643 = n20642 ^ n20637;
  assign n20644 = ~n20639 & n20643;
  assign n20645 = n20644 ^ n20637;
  assign n20646 = n20379 & ~n20645;
  assign n20647 = n20636 & ~n20646;
  assign n20648 = n20379 & n20380;
  assign n20649 = n20620 & n20627;
  assign n20650 = n20610 & n20626;
  assign n20651 = ~n20619 & ~n20650;
  assign n20652 = ~n20649 & n20651;
  assign n20653 = ~n20621 & n20652;
  assign n20654 = n20648 & ~n20653;
  assign n20655 = ~n20611 & n20642;
  assign n20656 = ~n20650 & n20655;
  assign n20657 = n20381 & ~n20656;
  assign n20658 = ~n20654 & ~n20657;
  assign n20659 = n20609 & n20627;
  assign n20660 = n20659 ^ n20614;
  assign n20661 = n20660 ^ n20659;
  assign n20662 = n20605 & n20620;
  assign n20663 = n20605 & n20626;
  assign n20664 = ~n20632 & ~n20663;
  assign n20665 = ~n20662 & n20664;
  assign n20666 = n20665 ^ n20659;
  assign n20667 = ~n20661 & ~n20666;
  assign n20668 = n20667 ^ n20659;
  assign n20669 = n20658 & ~n20668;
  assign n20670 = n20647 & n20669;
  assign n20671 = n20625 & n20670;
  assign n20672 = n20671 ^ n18593;
  assign n20673 = n19237 & n19244;
  assign n20674 = n19248 & n19287;
  assign n20675 = ~n19072 & ~n19273;
  assign n20676 = n19241 & ~n20675;
  assign n20677 = ~n20674 & ~n20676;
  assign n20678 = ~n20673 & n20677;
  assign n20679 = ~n19105 & n19262;
  assign n20680 = n19248 & n19251;
  assign n20681 = ~n20679 & ~n20680;
  assign n20682 = n19255 & n19269;
  assign n20683 = ~n19246 & ~n19268;
  assign n20684 = n19237 & ~n20683;
  assign n20685 = ~n20682 & ~n20684;
  assign n20686 = n20681 & n20685;
  assign n20687 = ~n19258 & ~n19268;
  assign n20688 = n19241 & ~n20687;
  assign n20689 = ~n19244 & ~n19286;
  assign n20690 = n19265 & ~n20689;
  assign n20691 = n19237 & n19264;
  assign n20692 = n19237 & n19273;
  assign n20693 = n19277 & ~n19286;
  assign n20694 = ~n19246 & n20693;
  assign n20695 = n19241 & ~n20694;
  assign n20696 = n19035 ^ n18893;
  assign n20697 = n20696 ^ n19068;
  assign n20698 = n18931 & n20697;
  assign n20699 = n19265 & n20698;
  assign n20700 = ~n20695 & ~n20699;
  assign n20701 = ~n20692 & n20700;
  assign n20702 = ~n20691 & n20701;
  assign n20703 = ~n19238 & n20702;
  assign n20704 = ~n20690 & n20703;
  assign n20705 = ~n20688 & n20704;
  assign n20706 = n20686 & n20705;
  assign n20707 = n20678 & n20706;
  assign n20708 = n20707 ^ n18297;
  assign n20709 = n20608 & n20621;
  assign n20710 = ~n20659 & ~n20662;
  assign n20711 = n20381 & ~n20710;
  assign n20712 = ~n20709 & ~n20711;
  assign n20713 = ~n20380 & n20640;
  assign n20714 = n20608 & n20650;
  assign n20715 = ~n20713 & ~n20714;
  assign n20716 = n20611 & n20617;
  assign n20717 = ~n20649 & n20664;
  assign n20718 = n20614 & ~n20717;
  assign n20719 = ~n20716 & ~n20718;
  assign n20720 = n20715 & n20719;
  assign n20721 = n20381 & n20628;
  assign n20722 = n20526 ^ n20489;
  assign n20723 = n20610 & ~n20722;
  assign n20724 = ~n20621 & ~n20723;
  assign n20725 = ~n20619 & n20724;
  assign n20726 = n20648 & ~n20725;
  assign n20727 = ~n20629 & ~n20649;
  assign n20728 = n20637 & n20727;
  assign n20729 = ~n20381 & n20728;
  assign n20730 = ~n20629 & n20651;
  assign n20731 = ~n20611 & n20730;
  assign n20732 = ~n20608 & n20731;
  assign n20733 = ~n20729 & ~n20732;
  assign n20734 = ~n20614 & n20733;
  assign n20735 = ~n20726 & ~n20734;
  assign n20736 = ~n20721 & n20735;
  assign n20737 = n20720 & n20736;
  assign n20738 = n20712 & n20737;
  assign n20739 = n20625 & n20738;
  assign n20740 = n20739 ^ n20044;
  assign n20741 = ~n20456 & ~n20473;
  assign n20742 = n20421 & ~n20741;
  assign n20743 = n20392 & n20448;
  assign n20744 = n20425 & n20743;
  assign n20745 = n20422 & n20471;
  assign n20746 = ~n20454 & n20465;
  assign n20747 = n20432 & n20746;
  assign n20748 = n20425 & ~n20747;
  assign n20749 = ~n20745 & ~n20748;
  assign n20750 = ~n20435 & ~n20441;
  assign n20751 = n20452 & n20750;
  assign n20752 = n20421 & ~n20751;
  assign n20753 = ~n20454 & ~n20743;
  assign n20754 = n20474 & n20753;
  assign n20755 = ~n20443 & n20754;
  assign n20756 = n20462 & ~n20755;
  assign n20757 = ~n20752 & ~n20756;
  assign n20758 = n20749 & n20757;
  assign n20759 = ~n20744 & n20758;
  assign n20760 = n20445 & n20759;
  assign n20761 = ~n20742 & n20760;
  assign n20762 = n20761 ^ n17839;
  assign n20763 = n20708 ^ x820;
  assign n20764 = n20054 & n20077;
  assign n20765 = ~n20511 & ~n20764;
  assign n20766 = ~n19944 & n20078;
  assign n20767 = ~n20072 & n20077;
  assign n20768 = ~n20766 & ~n20767;
  assign n20769 = n20099 & ~n20497;
  assign n20770 = ~n20098 & ~n20105;
  assign n20771 = ~n20083 & ~n20770;
  assign n20772 = ~n20069 & n20503;
  assign n20773 = ~n20073 & n20772;
  assign n20774 = ~n20086 & n20773;
  assign n20775 = n20058 & ~n20774;
  assign n20776 = ~n20071 & n20088;
  assign n20777 = n20050 & ~n20776;
  assign n20778 = n20067 & ~n20085;
  assign n20779 = n20077 & ~n20778;
  assign n20780 = ~n20777 & ~n20779;
  assign n20781 = ~n20775 & n20780;
  assign n20782 = ~n20495 & n20781;
  assign n20783 = ~n20771 & n20782;
  assign n20784 = ~n20769 & n20783;
  assign n20785 = n20768 & n20784;
  assign n20786 = n20765 & n20785;
  assign n20787 = n20057 & n20786;
  assign n20788 = n20787 ^ n18681;
  assign n20789 = n20788 ^ x825;
  assign n20790 = n20763 & n20789;
  assign n20791 = n19650 & n20548;
  assign n20792 = ~n19666 & n20528;
  assign n20793 = ~n20791 & ~n20792;
  assign n20794 = ~n19690 & n20536;
  assign n20795 = ~n19701 & n20553;
  assign n20796 = ~n20794 & ~n20795;
  assign n20797 = n20793 & n20796;
  assign n20798 = n20797 ^ n18946;
  assign n20799 = n20798 ^ x822;
  assign n20800 = n18791 & n18804;
  assign n20801 = n18783 & n18822;
  assign n20802 = ~n20800 & ~n20801;
  assign n20803 = n18787 & n18807;
  assign n20804 = n18783 & n18845;
  assign n20805 = ~n20803 & ~n20804;
  assign n20806 = n18783 & n18786;
  assign n20807 = n18787 & ~n18836;
  assign n20808 = ~n20806 & ~n20807;
  assign n20809 = ~n18455 & ~n18831;
  assign n20810 = ~n18790 & ~n18804;
  assign n20811 = n20809 & n20810;
  assign n20812 = n18787 & ~n20811;
  assign n20813 = n18785 & n18811;
  assign n20814 = n18813 & ~n20813;
  assign n20815 = ~n18455 & n20814;
  assign n20816 = n18791 & ~n20815;
  assign n20817 = ~n20812 & ~n20816;
  assign n20818 = ~n18810 & ~n18835;
  assign n20819 = ~n18830 & n20818;
  assign n20820 = n18800 & ~n20819;
  assign n20821 = n18783 & n18804;
  assign n20822 = ~n18796 & ~n18799;
  assign n20823 = n18791 & ~n20822;
  assign n20824 = ~n20821 & ~n20823;
  assign n20825 = ~n18801 & n18831;
  assign n20826 = ~n18807 & ~n20813;
  assign n20827 = ~n18790 & n20826;
  assign n20828 = ~n18594 & ~n20827;
  assign n20829 = ~n20825 & ~n20828;
  assign n20830 = n20824 & n20829;
  assign n20831 = ~n20820 & n20830;
  assign n20832 = n20817 & n20831;
  assign n20833 = n20808 & n20832;
  assign n20834 = n20805 & n20833;
  assign n20835 = n20802 & n20834;
  assign n20836 = ~n18856 & n20835;
  assign n20837 = n20836 ^ n18237;
  assign n20838 = n20837 ^ x821;
  assign n20839 = ~n20799 & n20838;
  assign n20840 = n19849 & n19874;
  assign n20841 = n19853 & n20338;
  assign n20842 = ~n20840 & ~n20841;
  assign n20843 = ~n19810 & ~n19900;
  assign n20844 = ~n19878 & n20843;
  assign n20845 = n19856 & ~n20844;
  assign n20846 = ~n19858 & ~n19888;
  assign n20847 = ~n20348 & ~n20846;
  assign n20848 = ~n19871 & ~n19883;
  assign n20849 = n19905 & n20848;
  assign n20850 = n19887 & ~n20849;
  assign n20851 = n19879 & n19901;
  assign n20852 = n19853 & ~n20851;
  assign n20853 = ~n20850 & ~n20852;
  assign n20854 = ~n20847 & n20853;
  assign n20855 = n19892 ^ n19848;
  assign n20856 = ~n19874 & ~n20338;
  assign n20857 = n20856 ^ n20848;
  assign n20858 = n20848 ^ n19811;
  assign n20859 = n20858 ^ n20848;
  assign n20860 = n20857 & ~n20859;
  assign n20861 = n20860 ^ n20848;
  assign n20862 = n20861 ^ n19892;
  assign n20863 = n20855 & n20862;
  assign n20864 = n20863 ^ n20860;
  assign n20865 = n20864 ^ n20848;
  assign n20866 = n20865 ^ n19848;
  assign n20867 = n19892 & n20866;
  assign n20868 = n20867 ^ n19892;
  assign n20869 = n20868 ^ n19848;
  assign n20870 = n20854 & ~n20869;
  assign n20871 = ~n20845 & n20870;
  assign n20872 = n20842 & n20871;
  assign n20873 = ~n19857 & n20872;
  assign n20874 = ~n19909 & n20873;
  assign n20875 = n19855 & n20874;
  assign n20876 = n20875 ^ n18621;
  assign n20877 = n20876 ^ x824;
  assign n20878 = n20839 & n20877;
  assign n20879 = n19369 & n19512;
  assign n20880 = n19509 & n19551;
  assign n20881 = ~n20879 & ~n20880;
  assign n20882 = n19517 & n19531;
  assign n20883 = n19509 & n19552;
  assign n20884 = ~n20882 & ~n20883;
  assign n20885 = n19531 & n19532;
  assign n20886 = ~n19542 & n19556;
  assign n20887 = ~n19547 & n20886;
  assign n20888 = ~n19506 & n20887;
  assign n20889 = n19369 & ~n20888;
  assign n20890 = ~n20885 & ~n20889;
  assign n20891 = ~n19523 & n19529;
  assign n20892 = n19518 & n19534;
  assign n20893 = n19509 & ~n20892;
  assign n20894 = ~n19506 & n19554;
  assign n20895 = ~n19537 & n20894;
  assign n20896 = n19507 & ~n19525;
  assign n20897 = ~n19544 & n20896;
  assign n20898 = ~n19531 & n20897;
  assign n20899 = ~n20895 & ~n20898;
  assign n20900 = n19539 & ~n20899;
  assign n20901 = n19368 & ~n20900;
  assign n20902 = ~n20893 & ~n20901;
  assign n20903 = ~n20891 & n20902;
  assign n20904 = n20890 & n20903;
  assign n20905 = n20884 & n20904;
  assign n20906 = n19528 & n20905;
  assign n20907 = n20881 & n20906;
  assign n20908 = n20907 ^ n18973;
  assign n20909 = n20908 ^ x823;
  assign n20910 = n20878 & ~n20909;
  assign n20911 = n20790 & n20910;
  assign n20912 = ~n20763 & n20789;
  assign n20913 = ~n20799 & ~n20838;
  assign n20914 = n20877 & n20913;
  assign n20915 = n20909 & n20914;
  assign n20916 = n20912 & n20915;
  assign n20917 = n20763 & ~n20789;
  assign n20918 = n20799 & ~n20838;
  assign n20919 = n20877 & n20918;
  assign n20920 = ~n20909 & n20919;
  assign n20921 = n20917 & n20920;
  assign n20922 = ~n20916 & ~n20921;
  assign n20923 = ~n20911 & n20922;
  assign n20924 = ~n20877 & n20909;
  assign n20925 = n20839 & n20924;
  assign n20926 = n20790 & n20925;
  assign n20927 = n20799 & n20838;
  assign n20928 = n20924 & n20927;
  assign n20929 = n20877 & n20927;
  assign n20930 = ~n20909 & n20929;
  assign n20931 = ~n20928 & ~n20930;
  assign n20932 = n20790 & ~n20931;
  assign n20933 = ~n20877 & ~n20909;
  assign n20934 = n20927 & n20933;
  assign n20935 = ~n20910 & ~n20934;
  assign n20936 = n20912 & ~n20935;
  assign n20937 = ~n20932 & ~n20936;
  assign n20938 = ~n20926 & n20937;
  assign n20939 = n20918 & n20933;
  assign n20940 = n20790 & n20939;
  assign n20941 = n20918 & n20924;
  assign n20942 = ~n20909 & n20914;
  assign n20943 = ~n20941 & ~n20942;
  assign n20944 = n20912 & ~n20943;
  assign n20945 = ~n20940 & ~n20944;
  assign n20946 = n20789 ^ n20763;
  assign n20947 = n20909 & n20929;
  assign n20948 = ~n20925 & ~n20947;
  assign n20949 = n20946 & ~n20948;
  assign n20950 = n20909 & n20919;
  assign n20951 = n20913 & n20933;
  assign n20952 = ~n20920 & ~n20951;
  assign n20953 = ~n20950 & n20952;
  assign n20954 = n20790 & ~n20953;
  assign n20955 = ~n20934 & ~n20951;
  assign n20956 = n20943 & n20955;
  assign n20957 = ~n20930 & n20956;
  assign n20958 = n20917 & ~n20957;
  assign n20959 = ~n20954 & ~n20958;
  assign n20960 = ~n20949 & n20959;
  assign n20961 = ~n20942 & ~n20950;
  assign n20962 = ~n20910 & ~n20925;
  assign n20963 = ~n20941 & n20962;
  assign n20964 = ~n20930 & n20963;
  assign n20965 = n20961 & n20964;
  assign n20966 = ~n20915 & n20965;
  assign n20967 = n20966 ^ n20912;
  assign n20968 = n20967 ^ n20912;
  assign n20969 = ~n20763 & ~n20789;
  assign n20970 = n20969 ^ n20912;
  assign n20971 = n20970 ^ n20912;
  assign n20972 = n20968 & n20971;
  assign n20973 = n20972 ^ n20912;
  assign n20974 = ~n20939 & n20973;
  assign n20975 = n20974 ^ n20912;
  assign n20976 = n20960 & ~n20975;
  assign n20977 = n20945 & n20976;
  assign n20978 = n20938 & n20977;
  assign n20979 = n20923 & n20978;
  assign n20980 = n20979 ^ n19390;
  assign n20981 = n20421 & n20428;
  assign n20982 = n20422 & ~n20451;
  assign n20983 = ~n20981 & ~n20982;
  assign n20984 = n20430 & n20446;
  assign n20985 = n20425 & n20984;
  assign n20986 = n20456 & n20462;
  assign n20987 = ~n20985 & ~n20986;
  assign n20988 = n20425 & ~n20457;
  assign n20989 = ~n20441 & ~n20456;
  assign n20990 = n20421 & ~n20989;
  assign n20991 = ~n20441 & ~n20473;
  assign n20992 = ~n20984 & n20991;
  assign n20993 = ~n20443 & n20992;
  assign n20994 = n20422 & ~n20993;
  assign n20995 = ~n20418 & ~n20463;
  assign n20996 = n20451 & n20995;
  assign n20997 = n20425 & ~n20996;
  assign n20998 = ~n20994 & ~n20997;
  assign n20999 = n20418 & ~n20422;
  assign n21000 = ~n20447 & n20753;
  assign n21001 = n20437 & ~n21000;
  assign n21002 = ~n20999 & ~n21001;
  assign n21003 = n20998 & n21002;
  assign n21004 = ~n20990 & n21003;
  assign n21005 = ~n20988 & n21004;
  assign n21006 = n20463 ^ n20419;
  assign n21007 = n21006 ^ n20463;
  assign n21008 = n20432 & ~n20435;
  assign n21009 = n21008 ^ n20463;
  assign n21010 = n21007 & ~n21009;
  assign n21011 = n21010 ^ n20463;
  assign n21012 = ~n20420 & n21011;
  assign n21013 = n21005 & ~n21012;
  assign n21014 = n20987 & n21013;
  assign n21015 = n20983 & n21014;
  assign n21016 = n20440 & n21015;
  assign n21017 = n21016 ^ n18027;
  assign n21018 = n20913 & n20924;
  assign n21019 = ~n20920 & ~n21018;
  assign n21020 = n20912 & ~n21019;
  assign n21021 = n20839 & n20933;
  assign n21022 = n21021 ^ n20969;
  assign n21023 = n21021 ^ n20790;
  assign n21024 = n21023 ^ n20790;
  assign n21025 = n20948 ^ n20790;
  assign n21026 = ~n21024 & n21025;
  assign n21027 = n21026 ^ n20790;
  assign n21028 = n21022 & n21027;
  assign n21029 = n21028 ^ n20969;
  assign n21030 = ~n21020 & ~n21029;
  assign n21031 = n20939 & n20969;
  assign n21032 = n20917 ^ n20909;
  assign n21033 = n21032 ^ n20917;
  assign n21034 = n20917 ^ n20790;
  assign n21035 = n21033 & n21034;
  assign n21036 = n21035 ^ n20917;
  assign n21037 = n20878 & n21036;
  assign n21038 = ~n21031 & ~n21037;
  assign n21039 = n20878 & n20909;
  assign n21040 = n20969 & n21039;
  assign n21041 = n20917 & n20941;
  assign n21042 = ~n21040 & ~n21041;
  assign n21043 = n20934 & n20969;
  assign n21044 = ~n20790 & ~n20969;
  assign n21045 = ~n20961 & ~n21044;
  assign n21046 = ~n21043 & ~n21045;
  assign n21047 = n20917 & ~n20931;
  assign n21048 = n20912 & ~n20964;
  assign n21049 = ~n21047 & ~n21048;
  assign n21050 = ~n20928 & ~n21018;
  assign n21051 = ~n20939 & n21050;
  assign n21052 = n20790 & ~n21051;
  assign n21053 = n20909 ^ n20877;
  assign n21054 = n21053 ^ n20877;
  assign n21055 = n20917 ^ n20877;
  assign n21056 = n21054 & ~n21055;
  assign n21057 = n21056 ^ n20877;
  assign n21058 = n20913 & ~n21057;
  assign n21059 = n21044 & n21058;
  assign n21060 = ~n21052 & ~n21059;
  assign n21061 = n21049 & n21060;
  assign n21062 = n21046 & n21061;
  assign n21063 = n21042 & n21062;
  assign n21064 = n21038 & n21063;
  assign n21065 = n20923 & n21064;
  assign n21066 = n21030 & n21065;
  assign n21067 = n21066 ^ n19766;
  assign n21068 = n19531 & ~n19548;
  assign n21069 = ~n19532 & n19539;
  assign n21070 = ~n19522 & n21069;
  assign n21071 = n19509 & ~n21070;
  assign n21072 = ~n21068 & ~n21071;
  assign n21073 = n19552 ^ n19332;
  assign n21074 = n21073 ^ n19552;
  assign n21075 = n19552 ^ n19537;
  assign n21076 = n21075 ^ n19552;
  assign n21077 = ~n21074 & n21076;
  assign n21078 = n21077 ^ n19552;
  assign n21079 = ~n19368 & n21078;
  assign n21080 = n21079 ^ n19552;
  assign n21081 = n21072 & ~n21080;
  assign n21082 = n19368 ^ n19332;
  assign n21083 = n19551 & ~n21082;
  assign n21084 = ~n19506 & n19556;
  assign n21085 = n19529 & ~n21084;
  assign n21086 = n19369 & n19514;
  assign n21087 = n19518 & ~n19533;
  assign n21088 = n19531 & ~n21087;
  assign n21089 = n19507 & ~n19537;
  assign n21090 = n19509 & ~n21089;
  assign n21091 = ~n21088 & ~n21090;
  assign n21092 = ~n21086 & n21091;
  assign n21093 = ~n19512 & ~n19517;
  assign n21094 = ~n19542 & n21093;
  assign n21095 = ~n19522 & n21094;
  assign n21096 = n21095 ^ n19521;
  assign n21097 = n21096 ^ n19521;
  assign n21098 = n19521 ^ n19368;
  assign n21099 = n21098 ^ n19521;
  assign n21100 = ~n21097 & n21099;
  assign n21101 = n21100 ^ n19521;
  assign n21102 = n21082 & n21101;
  assign n21103 = n21102 ^ n19521;
  assign n21104 = n21092 & ~n21103;
  assign n21105 = n20881 & n21104;
  assign n21106 = ~n21085 & n21105;
  assign n21107 = ~n21083 & n21106;
  assign n21108 = n21081 & n21107;
  assign n21109 = ~n19508 & n21108;
  assign n21110 = n21109 ^ n16189;
  assign n21111 = ~n20534 & n20536;
  assign n21112 = n20548 & n20561;
  assign n21113 = ~n21111 & ~n21112;
  assign n21114 = ~n20550 & n20553;
  assign n21115 = n20528 & ~n20543;
  assign n21116 = ~n21114 & ~n21115;
  assign n21117 = n21113 & n21116;
  assign n21118 = ~n20546 & n21117;
  assign n21119 = n21118 ^ n17607;
  assign n21120 = n21119 ^ x831;
  assign n21121 = n20876 ^ x826;
  assign n21122 = n21120 & n21121;
  assign n21123 = ~n19255 & ~n19272;
  assign n21124 = ~n19251 & n21123;
  assign n21125 = n19248 & ~n21124;
  assign n21126 = n19264 & ~n19270;
  assign n21127 = ~n19070 & ~n19287;
  assign n21128 = n19241 & ~n21127;
  assign n21129 = n19288 & n19291;
  assign n21130 = n19237 & ~n21129;
  assign n21131 = ~n21128 & ~n21130;
  assign n21132 = ~n21126 & n21131;
  assign n21133 = n19248 & n19268;
  assign n21134 = ~n19272 & n20675;
  assign n21135 = ~n19262 & n21134;
  assign n21136 = ~n19258 & n21135;
  assign n21137 = n19269 & ~n21136;
  assign n21138 = ~n21133 & ~n21137;
  assign n21139 = n21132 & n21138;
  assign n21140 = n19261 & n21139;
  assign n21141 = ~n19253 & n21140;
  assign n21142 = ~n21125 & n21141;
  assign n21143 = n20678 & n21142;
  assign n21144 = ~n20691 & n21143;
  assign n21145 = ~n19315 & n21144;
  assign n21146 = ~n19246 & n21145;
  assign n21147 = n21146 ^ n18640;
  assign n21148 = n21147 ^ x828;
  assign n21149 = n20788 ^ x827;
  assign n21150 = ~n21148 & ~n21149;
  assign n21151 = n20762 ^ x830;
  assign n21152 = n20121 & n20208;
  assign n21153 = n20122 & n20232;
  assign n21154 = n20191 & n20211;
  assign n21155 = ~n21153 & ~n21154;
  assign n21156 = ~n21152 & n21155;
  assign n21157 = n20120 & n20197;
  assign n21158 = n20122 & ~n20239;
  assign n21159 = ~n21157 & ~n21158;
  assign n21160 = ~n20202 & n20245;
  assign n21161 = ~n20582 & n21160;
  assign n21162 = ~n20212 & n21161;
  assign n21163 = n20194 & ~n21162;
  assign n21164 = n20203 & n20233;
  assign n21165 = n21164 ^ n20120;
  assign n21166 = n21165 ^ n21164;
  assign n21167 = n20246 & n20578;
  assign n21168 = n21167 ^ n21164;
  assign n21169 = n21166 & n21168;
  assign n21170 = n21169 ^ n21164;
  assign n21171 = ~n20121 & ~n21170;
  assign n21172 = ~n21163 & ~n21171;
  assign n21173 = n21159 & n21172;
  assign n21174 = n20572 & n21173;
  assign n21175 = n21156 & n21174;
  assign n21176 = ~n20210 & n21175;
  assign n21177 = n20193 & n21176;
  assign n21178 = ~n20567 & n21177;
  assign n21179 = n21178 ^ n18705;
  assign n21180 = n21179 ^ x829;
  assign n21181 = ~n21151 & ~n21180;
  assign n21182 = n21150 & n21181;
  assign n21183 = n21122 & n21182;
  assign n21184 = ~n21120 & n21121;
  assign n21185 = ~n21148 & n21149;
  assign n21186 = n21151 & ~n21180;
  assign n21187 = n21185 & n21186;
  assign n21188 = n21184 & n21187;
  assign n21189 = ~n21120 & ~n21121;
  assign n21190 = n21150 & n21186;
  assign n21191 = n21148 & ~n21149;
  assign n21192 = n21181 & n21191;
  assign n21193 = ~n21190 & ~n21192;
  assign n21194 = n21189 & ~n21193;
  assign n21195 = ~n21188 & ~n21194;
  assign n21196 = ~n21183 & n21195;
  assign n21197 = ~n21151 & n21180;
  assign n21198 = n21185 & n21197;
  assign n21199 = n21184 & n21198;
  assign n21200 = n21120 & ~n21121;
  assign n21201 = n21192 & n21200;
  assign n21202 = ~n21199 & ~n21201;
  assign n21203 = n21148 & n21149;
  assign n21204 = n21180 ^ n21151;
  assign n21205 = n21203 & ~n21204;
  assign n21206 = n21122 & n21205;
  assign n21207 = n21202 & ~n21206;
  assign n21208 = n21198 & n21200;
  assign n21209 = n21182 & n21184;
  assign n21210 = ~n21208 & ~n21209;
  assign n21211 = n21151 & n21180;
  assign n21212 = n21203 & n21211;
  assign n21213 = ~n21198 & ~n21212;
  assign n21214 = n21189 & ~n21213;
  assign n21215 = n21191 & n21211;
  assign n21216 = n21184 & n21215;
  assign n21217 = n21197 & n21203;
  assign n21218 = n21122 & n21217;
  assign n21219 = ~n21216 & ~n21218;
  assign n21220 = n21186 & n21191;
  assign n21221 = n21200 & n21220;
  assign n21222 = ~n21122 & ~n21189;
  assign n21223 = n21181 & n21185;
  assign n21224 = ~n21222 & n21223;
  assign n21225 = ~n21180 & n21203;
  assign n21226 = n21191 & n21197;
  assign n21227 = ~n21190 & ~n21226;
  assign n21228 = ~n21225 & n21227;
  assign n21229 = n21184 & ~n21228;
  assign n21230 = ~n21224 & ~n21229;
  assign n21231 = n21185 & n21211;
  assign n21232 = ~n21121 & n21231;
  assign n21233 = n21151 & n21203;
  assign n21234 = n21227 & ~n21233;
  assign n21235 = n21200 & ~n21234;
  assign n21236 = n21121 ^ n21120;
  assign n21241 = ~n21220 & ~n21226;
  assign n21237 = n21150 & n21197;
  assign n21238 = n21150 & n21211;
  assign n21239 = ~n21220 & ~n21238;
  assign n21240 = ~n21237 & n21239;
  assign n21242 = n21241 ^ n21240;
  assign n21243 = n21241 ^ n21121;
  assign n21244 = n21243 ^ n21241;
  assign n21245 = n21242 & n21244;
  assign n21246 = n21245 ^ n21241;
  assign n21247 = ~n21236 & ~n21246;
  assign n21248 = ~n21235 & ~n21247;
  assign n21249 = ~n21232 & n21248;
  assign n21250 = n21230 & n21249;
  assign n21251 = ~n21221 & n21250;
  assign n21252 = n21219 & n21251;
  assign n21253 = ~n21214 & n21252;
  assign n21254 = n21210 & n21253;
  assign n21255 = n21207 & n21254;
  assign n21256 = n21196 & n21255;
  assign n21257 = n21256 ^ n19637;
  assign n21258 = ~n20187 & n20568;
  assign n21259 = ~n20242 & n21258;
  assign n21260 = ~n20232 & n21259;
  assign n21261 = n20211 & ~n21260;
  assign n21262 = n20230 & n21162;
  assign n21263 = n20206 & ~n21262;
  assign n21264 = ~n21261 & ~n21263;
  assign n21265 = n20578 ^ n20121;
  assign n21266 = n21265 ^ n20578;
  assign n21267 = n20578 ^ n20234;
  assign n21268 = n21267 ^ n20578;
  assign n21269 = n21266 & ~n21268;
  assign n21270 = n21269 ^ n20578;
  assign n21271 = ~n20120 & ~n21270;
  assign n21272 = n21271 ^ n20578;
  assign n21273 = n21264 & n21272;
  assign n21274 = n21156 & n21273;
  assign n21275 = n20205 & n21274;
  assign n21276 = n20570 & n21275;
  assign n21277 = ~n20567 & n21276;
  assign n21278 = n21277 ^ n18370;
  assign n21279 = n20762 ^ x784;
  assign n21280 = ~n19552 & n20896;
  assign n21281 = n19531 & ~n21280;
  assign n21282 = n19518 & ~n19525;
  assign n21283 = ~n19544 & n21282;
  assign n21284 = ~n19522 & n21283;
  assign n21285 = n19369 & ~n21284;
  assign n21286 = n19476 ^ n19424;
  assign n21287 = n19424 ^ n19391;
  assign n21288 = n21287 ^ n19501;
  assign n21289 = n21288 ^ n19501;
  assign n21290 = n21289 ^ n21288;
  assign n21291 = n21288 ^ n19476;
  assign n21292 = n21291 ^ n21288;
  assign n21293 = ~n21290 & ~n21292;
  assign n21294 = n21293 ^ n21288;
  assign n21295 = ~n21286 & n21294;
  assign n21296 = n21295 ^ n21288;
  assign n21297 = n19529 & n21296;
  assign n21298 = ~n21285 & ~n21297;
  assign n21299 = ~n21281 & n21298;
  assign n21300 = n20886 ^ n19522;
  assign n21301 = n21300 ^ n19522;
  assign n21302 = n19522 ^ n19332;
  assign n21303 = n21302 ^ n19522;
  assign n21304 = ~n21301 & n21303;
  assign n21305 = n21304 ^ n19522;
  assign n21306 = ~n19368 & n21305;
  assign n21307 = n21306 ^ n19522;
  assign n21308 = n21299 & ~n21307;
  assign n21309 = n19536 & n21308;
  assign n21310 = n20884 & n21309;
  assign n21311 = ~n19520 & n21310;
  assign n21312 = ~n19508 & n21311;
  assign n21313 = n20881 & n21312;
  assign n21314 = n21313 ^ n17878;
  assign n21315 = n21314 ^ x789;
  assign n21316 = ~n21279 & n21315;
  assign n21317 = n21119 ^ x785;
  assign n21318 = n18783 & n18823;
  assign n21319 = ~n18455 & ~n18852;
  assign n21320 = n18787 & ~n21319;
  assign n21321 = ~n21318 & ~n21320;
  assign n21322 = ~n18799 & ~n18831;
  assign n21323 = n18787 & ~n21322;
  assign n21324 = ~n18812 & ~n20813;
  assign n21325 = n18783 & ~n21324;
  assign n21326 = ~n21323 & ~n21325;
  assign n21327 = ~n18786 & ~n18807;
  assign n21328 = n18800 & ~n21327;
  assign n21329 = n18791 & n18852;
  assign n21330 = n18783 & ~n20809;
  assign n21331 = ~n21329 & ~n21330;
  assign n21332 = ~n18796 & n20810;
  assign n21333 = n18800 & ~n21332;
  assign n21334 = n18787 & ~n18825;
  assign n21335 = ~n21333 & ~n21334;
  assign n21336 = n21331 & n21335;
  assign n21337 = n20824 & n21336;
  assign n21338 = n20805 & n21337;
  assign n21339 = ~n18847 & n21338;
  assign n21340 = ~n21328 & n21339;
  assign n21341 = n21326 & n21340;
  assign n21342 = n18836 ^ n18791;
  assign n21343 = n18836 ^ n18823;
  assign n21344 = n21343 ^ n18823;
  assign n21345 = n18823 ^ n18800;
  assign n21346 = ~n21344 & ~n21345;
  assign n21347 = n21346 ^ n18823;
  assign n21348 = ~n21342 & ~n21347;
  assign n21349 = n21348 ^ n18791;
  assign n21350 = n21341 & ~n21349;
  assign n21351 = n21321 & n21350;
  assign n21352 = n20802 & n21351;
  assign n21353 = n21352 ^ n17812;
  assign n21354 = n21353 ^ x787;
  assign n21355 = n21317 & ~n21354;
  assign n21356 = ~n19916 & n20061;
  assign n21357 = n20084 & ~n20497;
  assign n21358 = ~n21356 & ~n21357;
  assign n21359 = n20050 & n20065;
  assign n21360 = ~n20065 & n20101;
  assign n21361 = n20072 & n21360;
  assign n21362 = n20058 & ~n21361;
  assign n21363 = n19945 & ~n20504;
  assign n21364 = ~n20054 & n20079;
  assign n21365 = ~n20085 & n21364;
  assign n21366 = n20050 & ~n21365;
  assign n21367 = n20045 ^ n19983;
  assign n21368 = n21367 ^ n19983;
  assign n21369 = n20046 ^ n19983;
  assign n21370 = n21369 ^ n19983;
  assign n21371 = ~n21368 & ~n21370;
  assign n21372 = n21371 ^ n19983;
  assign n21373 = ~n20016 & ~n21372;
  assign n21374 = ~n20099 & ~n21373;
  assign n21375 = n20077 & ~n21374;
  assign n21376 = ~n21366 & ~n21375;
  assign n21377 = ~n21363 & n21376;
  assign n21378 = n20765 & n21377;
  assign n21379 = ~n21362 & n21378;
  assign n21380 = ~n21359 & n21379;
  assign n21381 = n21358 & n21380;
  assign n21382 = n20493 & n21381;
  assign n21383 = ~n20771 & n21382;
  assign n21384 = n21383 ^ n17771;
  assign n21385 = n21384 ^ x788;
  assign n21386 = n19856 & n19874;
  assign n21387 = n19849 & n20338;
  assign n21388 = ~n21386 & ~n21387;
  assign n21389 = n19883 & ~n20348;
  assign n21390 = n19848 & n19882;
  assign n21391 = ~n19868 & ~n19900;
  assign n21392 = ~n19888 & n21391;
  assign n21393 = n19849 & ~n21392;
  assign n21394 = n20350 & n20848;
  assign n21395 = ~n19882 & n21394;
  assign n21396 = n19853 & ~n21395;
  assign n21397 = ~n21393 & ~n21396;
  assign n21398 = n19879 & n20843;
  assign n21399 = n19887 & ~n21398;
  assign n21400 = ~n19856 & ~n21399;
  assign n21401 = n21400 ^ n19887;
  assign n21402 = ~n19810 & ~n19864;
  assign n21403 = ~n19858 & n21402;
  assign n21404 = n21403 ^ n21400;
  assign n21405 = n21404 ^ n21403;
  assign n21406 = ~n19858 & n19875;
  assign n21407 = n21406 ^ n21403;
  assign n21408 = n21405 & ~n21407;
  assign n21409 = n21408 ^ n21403;
  assign n21410 = ~n21401 & ~n21409;
  assign n21411 = n21410 ^ n19887;
  assign n21412 = n21397 & ~n21411;
  assign n21413 = ~n19850 & n21412;
  assign n21414 = n19860 & n21413;
  assign n21415 = ~n21390 & n21414;
  assign n21416 = ~n21389 & n21415;
  assign n21417 = n21388 & n21416;
  assign n21418 = n20344 & n21417;
  assign n21419 = n21418 ^ n17643;
  assign n21420 = n21419 ^ x786;
  assign n21421 = ~n21385 & n21420;
  assign n21422 = n21355 & n21421;
  assign n21423 = n21316 & n21422;
  assign n21424 = n21279 & n21315;
  assign n21425 = ~n21317 & ~n21354;
  assign n21426 = n21385 & n21420;
  assign n21427 = n21425 & n21426;
  assign n21428 = ~n21317 & n21354;
  assign n21429 = ~n21385 & ~n21420;
  assign n21430 = n21428 & n21429;
  assign n21431 = ~n21427 & ~n21430;
  assign n21432 = n21424 & ~n21431;
  assign n21433 = ~n21423 & ~n21432;
  assign n21434 = n21421 & n21425;
  assign n21435 = n21424 & n21434;
  assign n21436 = n21385 & ~n21420;
  assign n21437 = n21425 & n21436;
  assign n21438 = ~n21315 & n21437;
  assign n21439 = ~n21435 & ~n21438;
  assign n21440 = n21424 & n21437;
  assign n21441 = n21428 & n21436;
  assign n21442 = ~n21315 & n21441;
  assign n21443 = ~n21440 & ~n21442;
  assign n21444 = ~n21279 & ~n21315;
  assign n21445 = n21426 & n21428;
  assign n21446 = n21355 & n21426;
  assign n21447 = n21317 & n21354;
  assign n21448 = n21421 & n21447;
  assign n21449 = n21436 & n21447;
  assign n21450 = ~n21448 & ~n21449;
  assign n21451 = ~n21422 & n21450;
  assign n21452 = ~n21446 & n21451;
  assign n21453 = ~n21430 & n21452;
  assign n21454 = ~n21445 & n21453;
  assign n21455 = n21444 & ~n21454;
  assign n21456 = n21279 & ~n21315;
  assign n21457 = n21425 & n21429;
  assign n21458 = n21355 & n21436;
  assign n21459 = n21426 & n21447;
  assign n21460 = n21429 & n21447;
  assign n21461 = ~n21459 & ~n21460;
  assign n21462 = ~n21458 & n21461;
  assign n21463 = ~n21457 & n21462;
  assign n21464 = ~n21434 & n21463;
  assign n21465 = ~n21448 & n21464;
  assign n21466 = n21456 & ~n21465;
  assign n21467 = ~n21455 & ~n21466;
  assign n21468 = ~n21446 & n21461;
  assign n21469 = n21316 & ~n21468;
  assign n21470 = n21424 ^ n21316;
  assign n21475 = n21355 & n21429;
  assign n21471 = n21421 & n21428;
  assign n21476 = ~n21446 & ~n21459;
  assign n21477 = ~n21471 & n21476;
  assign n21478 = ~n21475 & n21477;
  assign n21472 = ~n21441 & ~n21471;
  assign n21473 = ~n21445 & n21472;
  assign n21474 = ~n21457 & n21473;
  assign n21479 = n21478 ^ n21474;
  assign n21480 = n21478 ^ n21424;
  assign n21481 = n21480 ^ n21478;
  assign n21482 = ~n21479 & ~n21481;
  assign n21483 = n21482 ^ n21478;
  assign n21484 = n21470 & ~n21483;
  assign n21485 = n21484 ^ n21316;
  assign n21486 = ~n21469 & ~n21485;
  assign n21487 = n21467 & n21486;
  assign n21488 = n21443 & n21487;
  assign n21489 = n21439 & n21488;
  assign n21490 = n21433 & n21489;
  assign n21491 = n21490 ^ n20015;
  assign n21492 = n21424 & n21475;
  assign n21493 = n21316 & n21430;
  assign n21494 = ~n21492 & ~n21493;
  assign n21495 = ~n21315 & n21422;
  assign n21496 = n21428 ^ n21426;
  assign n21497 = n21444 & n21496;
  assign n21498 = ~n21495 & ~n21497;
  assign n21499 = n21450 & ~n21460;
  assign n21500 = n21456 & ~n21499;
  assign n21501 = n21452 & ~n21471;
  assign n21502 = ~n21437 & n21501;
  assign n21503 = n21316 & ~n21502;
  assign n21504 = ~n21500 & ~n21503;
  assign n21505 = n21498 & n21504;
  assign n21506 = n21424 & ~n21462;
  assign n21507 = n21445 ^ n21279;
  assign n21510 = ~n21427 & ~n21457;
  assign n21511 = ~n21471 & n21510;
  assign n21508 = ~n21434 & ~n21437;
  assign n21509 = ~n21475 & n21508;
  assign n21512 = n21511 ^ n21509;
  assign n21513 = n21511 ^ n21315;
  assign n21514 = n21513 ^ n21511;
  assign n21515 = n21512 & ~n21514;
  assign n21516 = n21515 ^ n21511;
  assign n21517 = n21516 ^ n21445;
  assign n21518 = ~n21507 & ~n21517;
  assign n21519 = n21518 ^ n21515;
  assign n21520 = n21519 ^ n21511;
  assign n21521 = n21520 ^ n21279;
  assign n21522 = ~n21445 & n21521;
  assign n21523 = n21522 ^ n21445;
  assign n21524 = n21523 ^ n21279;
  assign n21525 = ~n21506 & n21524;
  assign n21526 = n21505 & n21525;
  assign n21527 = n21445 ^ n21315;
  assign n21528 = n21527 ^ n21445;
  assign n21529 = n21475 ^ n21445;
  assign n21530 = ~n21528 & n21529;
  assign n21531 = n21530 ^ n21445;
  assign n21532 = ~n21279 & n21531;
  assign n21533 = n21526 & ~n21532;
  assign n21534 = n21494 & n21533;
  assign n21535 = n21534 ^ n19423;
  assign n21536 = n19246 & n19269;
  assign n21537 = n19288 & n21134;
  assign n21538 = n19241 & ~n21537;
  assign n21539 = ~n21536 & ~n21538;
  assign n21540 = n19265 & ~n19291;
  assign n21541 = ~n19251 & ~n19287;
  assign n21542 = n19237 & ~n21541;
  assign n21543 = ~n19255 & n20687;
  assign n21544 = ~n19105 & ~n21543;
  assign n21545 = ~n21542 & ~n21544;
  assign n21546 = ~n21540 & n21545;
  assign n21547 = n21539 & n21546;
  assign n21548 = n19250 & n21547;
  assign n21549 = n19267 & n21548;
  assign n21550 = ~n21125 & n21549;
  assign n21551 = ~n20691 & n21550;
  assign n21552 = ~n19238 & n21551;
  assign n21553 = ~n19315 & n21552;
  assign n21554 = n21553 ^ n18072;
  assign n21555 = n20642 & n20651;
  assign n21556 = ~n20615 & n21555;
  assign n21557 = n20648 & ~n21556;
  assign n21558 = n20610 ^ n20605;
  assign n21559 = ~n20722 & n21558;
  assign n21560 = n21559 ^ n20605;
  assign n21561 = n20637 & ~n21560;
  assign n21562 = n21561 ^ n20381;
  assign n21563 = n21562 ^ n21561;
  assign n21564 = ~n20632 & n20710;
  assign n21565 = n21564 ^ n21561;
  assign n21566 = n21565 ^ n21561;
  assign n21567 = ~n21563 & ~n21566;
  assign n21568 = n21567 ^ n21561;
  assign n21569 = ~n20608 & ~n21568;
  assign n21570 = n21569 ^ n21561;
  assign n21571 = ~n21557 & n21570;
  assign n21572 = n20723 ^ n20651;
  assign n21573 = n20380 ^ n20379;
  assign n21574 = n21573 ^ n20380;
  assign n21575 = n20651 ^ n20380;
  assign n21576 = n21574 & ~n21575;
  assign n21577 = n21576 ^ n20380;
  assign n21578 = ~n21572 & ~n21577;
  assign n21579 = n21578 ^ n20723;
  assign n21580 = n20727 & ~n21579;
  assign n21581 = ~n20640 & n21580;
  assign n21582 = ~n20379 & ~n21581;
  assign n21583 = n21571 & ~n21582;
  assign n21584 = n20712 & n21583;
  assign n21585 = n20613 & n21584;
  assign n21586 = n21585 ^ n19733;
  assign n21587 = n18791 & n18845;
  assign n21588 = ~n18801 & ~n20826;
  assign n21589 = ~n18799 & n20818;
  assign n21590 = n18791 & ~n21589;
  assign n21591 = ~n18796 & ~n18822;
  assign n21592 = n18787 & ~n21591;
  assign n21593 = ~n21590 & ~n21592;
  assign n21594 = ~n21588 & n21593;
  assign n21595 = n18783 & ~n20822;
  assign n21596 = ~n18812 & n20811;
  assign n21597 = ~n18822 & n21596;
  assign n21598 = n18800 & ~n21597;
  assign n21599 = ~n21595 & ~n21598;
  assign n21600 = n21594 & n21599;
  assign n21601 = ~n20804 & n21600;
  assign n21602 = ~n21587 & n21601;
  assign n21603 = n20808 & n21602;
  assign n21604 = n21321 & n21603;
  assign n21605 = n18794 & n21604;
  assign n21606 = n20802 & n21605;
  assign n21607 = ~n18856 & n21606;
  assign n21608 = n21607 ^ n16902;
  assign n21609 = n20263 & n20304;
  assign n21610 = n19572 & ~n20269;
  assign n21611 = ~n21609 & ~n21610;
  assign n21612 = ~n20261 & ~n20289;
  assign n21613 = n20263 & ~n21612;
  assign n21614 = n20263 & n20274;
  assign n21615 = ~n20265 & ~n20305;
  assign n21616 = ~n20292 & n21615;
  assign n21617 = n20294 & ~n21616;
  assign n21618 = ~n21614 & ~n21617;
  assign n21619 = ~n20278 & n20297;
  assign n21620 = ~n19571 & n20284;
  assign n21621 = ~n21619 & ~n21620;
  assign n21622 = ~n20283 & ~n20315;
  assign n21623 = n19572 & ~n21622;
  assign n21624 = ~n20309 & ~n20314;
  assign n21625 = ~n20308 & n21624;
  assign n21626 = ~n20268 & n21625;
  assign n21627 = n20294 & ~n21626;
  assign n21628 = n20310 & ~n20315;
  assign n21629 = ~n20280 & n21628;
  assign n21630 = n20276 & ~n21629;
  assign n21631 = ~n21627 & ~n21630;
  assign n21632 = ~n21623 & n21631;
  assign n21633 = n21621 & n21632;
  assign n21634 = n21618 & n21633;
  assign n21635 = ~n21613 & n21634;
  assign n21636 = n20291 & n21635;
  assign n21637 = ~n20332 & n21636;
  assign n21638 = n21611 & n21637;
  assign n21639 = ~n20275 & n21638;
  assign n21640 = n20271 & n21639;
  assign n21641 = n21640 ^ n19607;
  assign n21642 = ~n20423 & n20447;
  assign n21643 = ~n20443 & ~n20449;
  assign n21644 = ~n20463 & n21643;
  assign n21645 = n20425 & ~n21644;
  assign n21646 = ~n21642 & ~n21645;
  assign n21647 = n20432 & ~n20984;
  assign n21648 = n20422 & ~n21647;
  assign n21649 = n20392 & n20427;
  assign n21650 = ~n20425 & n21649;
  assign n21651 = n20991 & n20995;
  assign n21652 = ~n20454 & n21651;
  assign n21653 = ~n20435 & n21652;
  assign n21654 = n20462 & ~n21653;
  assign n21655 = ~n21650 & ~n21654;
  assign n21656 = ~n21648 & n21655;
  assign n21657 = n21646 & n21656;
  assign n21658 = ~n20444 & n21657;
  assign n21659 = ~n20483 & n21658;
  assign n21660 = ~n20744 & n21659;
  assign n21661 = n20987 & n21660;
  assign n21662 = n20983 & n21661;
  assign n21663 = ~n20742 & n21662;
  assign n21664 = n20434 & n21663;
  assign n21665 = n21664 ^ n18324;
  assign n21666 = n20912 & n20929;
  assign n21667 = ~n21018 & ~n21021;
  assign n21668 = n20931 & n21667;
  assign n21669 = ~n20914 & n21668;
  assign n21670 = n20969 & ~n21669;
  assign n21671 = n20917 & ~n20948;
  assign n21674 = ~n20950 & n21667;
  assign n21672 = n20955 & n20961;
  assign n21673 = ~n20941 & n21672;
  assign n21675 = n21674 ^ n21673;
  assign n21676 = n21675 ^ n21674;
  assign n21677 = n21674 ^ n20789;
  assign n21678 = n21677 ^ n21674;
  assign n21679 = ~n21676 & n21678;
  assign n21680 = n21679 ^ n21674;
  assign n21681 = ~n20946 & ~n21680;
  assign n21682 = n21681 ^ n21674;
  assign n21683 = ~n21671 & n21682;
  assign n21684 = ~n21670 & n21683;
  assign n21685 = ~n21666 & n21684;
  assign n21686 = n20922 & n21685;
  assign n21687 = n21042 & n21686;
  assign n21688 = n21038 & n21687;
  assign n21689 = n20937 & n21688;
  assign n21690 = n21689 ^ n19982;
  assign n21691 = n20637 & ~n20659;
  assign n21692 = n20617 & ~n21691;
  assign n21693 = ~n20619 & n21564;
  assign n21694 = n20381 & ~n21693;
  assign n21695 = ~n21692 & ~n21694;
  assign n21696 = ~n20640 & ~n20723;
  assign n21697 = ~n20650 & n21696;
  assign n21698 = n20608 & ~n21697;
  assign n21699 = ~n20606 & n20727;
  assign n21700 = n20648 & ~n21699;
  assign n21701 = ~n20650 & n20724;
  assign n21702 = n20381 & ~n21701;
  assign n21703 = n20648 & ~n21697;
  assign n21704 = ~n21702 & ~n21703;
  assign n21705 = n20637 & n20710;
  assign n21706 = n20608 & ~n21705;
  assign n21707 = ~n20611 & n20652;
  assign n21708 = n20617 & ~n21707;
  assign n21709 = ~n21706 & ~n21708;
  assign n21710 = n21704 & n21709;
  assign n21711 = ~n21700 & n21710;
  assign n21712 = ~n21698 & n21711;
  assign n21713 = n21695 & n21712;
  assign n21714 = ~n20616 & n21713;
  assign n21715 = n21714 ^ n19475;
  assign n21716 = n21200 & n21205;
  assign n21717 = ~n21215 & ~n21238;
  assign n21718 = n21184 & ~n21717;
  assign n21719 = ~n21221 & ~n21718;
  assign n21720 = n21122 & n21190;
  assign n21721 = n21182 & n21200;
  assign n21722 = n21186 & n21203;
  assign n21723 = ~n21223 & ~n21722;
  assign n21724 = n21184 & ~n21723;
  assign n21725 = ~n21721 & ~n21724;
  assign n21726 = ~n21720 & n21725;
  assign n21727 = n21189 & n21238;
  assign n21728 = n21184 & n21237;
  assign n21729 = n21122 & n21192;
  assign n21730 = ~n21728 & ~n21729;
  assign n21731 = ~n21727 & n21730;
  assign n21732 = ~n21217 & ~n21231;
  assign n21733 = ~n21238 & n21732;
  assign n21734 = n21122 & ~n21733;
  assign n21735 = ~n21222 & n21225;
  assign n21736 = ~n21187 & ~n21226;
  assign n21737 = n21200 & ~n21736;
  assign n21738 = ~n21735 & ~n21737;
  assign n21739 = ~n21734 & n21738;
  assign n21740 = n21215 ^ n21120;
  assign n21741 = n21740 ^ n21215;
  assign n21742 = n21217 ^ n21215;
  assign n21743 = n21742 ^ n21215;
  assign n21744 = ~n21741 & n21743;
  assign n21745 = n21744 ^ n21215;
  assign n21746 = n21121 & n21745;
  assign n21747 = n21746 ^ n21215;
  assign n21748 = n21739 & ~n21747;
  assign n21749 = ~n21214 & n21748;
  assign n21750 = n21210 & n21749;
  assign n21751 = n21731 & n21750;
  assign n21752 = n21726 & n21751;
  assign n21753 = n21719 & n21752;
  assign n21754 = ~n21716 & n21753;
  assign n21755 = n21196 & n21754;
  assign n21756 = n21755 ^ n19805;
  assign n21757 = n21554 ^ x792;
  assign n21758 = n21017 ^ x793;
  assign n21759 = n18858 ^ x794;
  assign n21760 = n21314 ^ x791;
  assign n21761 = n21759 & n21760;
  assign n21762 = ~n21758 & n21761;
  assign n21763 = ~n21757 & n21762;
  assign n21764 = n21384 ^ x790;
  assign n21765 = n20603 ^ x795;
  assign n21766 = ~n21764 & n21765;
  assign n21767 = n21763 & n21766;
  assign n21768 = n21757 & n21758;
  assign n21769 = ~n21760 & n21768;
  assign n21770 = n21759 & n21769;
  assign n21771 = n21764 & n21765;
  assign n21772 = n21770 & n21771;
  assign n21773 = ~n21767 & ~n21772;
  assign n21774 = n21761 & n21768;
  assign n21775 = n21766 & n21774;
  assign n21776 = ~n21764 & ~n21765;
  assign n21777 = n21770 & n21776;
  assign n21778 = n21764 & ~n21765;
  assign n21779 = ~n21758 & ~n21760;
  assign n21780 = ~n21757 & n21779;
  assign n21781 = ~n21759 & n21780;
  assign n21782 = n21757 & n21779;
  assign n21783 = n21759 & n21782;
  assign n21784 = ~n21781 & ~n21783;
  assign n21785 = n21778 & ~n21784;
  assign n21786 = ~n21777 & ~n21785;
  assign n21787 = ~n21775 & n21786;
  assign n21788 = n21759 & n21780;
  assign n21789 = n21776 & n21788;
  assign n21790 = ~n21757 & n21758;
  assign n21791 = ~n21760 & n21790;
  assign n21792 = ~n21759 & n21791;
  assign n21793 = ~n21770 & ~n21792;
  assign n21794 = n21778 & ~n21793;
  assign n21795 = ~n21789 & ~n21794;
  assign n21796 = n21759 & n21791;
  assign n21797 = n21771 & n21796;
  assign n21798 = ~n21759 & n21760;
  assign n21799 = n21790 & n21798;
  assign n21800 = ~n21758 & n21798;
  assign n21801 = n21757 & n21800;
  assign n21802 = ~n21799 & ~n21801;
  assign n21803 = n21766 & ~n21802;
  assign n21804 = n21757 & n21762;
  assign n21805 = n21778 & n21804;
  assign n21806 = n21766 & ~n21784;
  assign n21807 = ~n21805 & ~n21806;
  assign n21808 = n21768 & n21798;
  assign n21809 = ~n21799 & ~n21804;
  assign n21810 = ~n21763 & n21809;
  assign n21811 = ~n21808 & n21810;
  assign n21812 = n21776 & ~n21811;
  assign n21813 = ~n21801 & n21810;
  assign n21814 = n21771 & ~n21813;
  assign n21815 = ~n21812 & ~n21814;
  assign n21816 = n21766 & n21791;
  assign n21817 = ~n21757 & n21800;
  assign n21818 = n21761 & n21790;
  assign n21819 = ~n21808 & ~n21818;
  assign n21820 = ~n21817 & n21819;
  assign n21821 = n21778 & ~n21820;
  assign n21822 = ~n21759 & n21769;
  assign n21823 = ~n21759 & n21782;
  assign n21824 = ~n21822 & ~n21823;
  assign n21825 = ~n21766 & ~n21778;
  assign n21826 = ~n21824 & n21825;
  assign n21827 = ~n21821 & ~n21826;
  assign n21828 = ~n21816 & n21827;
  assign n21829 = n21815 & n21828;
  assign n21830 = n21807 & n21829;
  assign n21831 = ~n21803 & n21830;
  assign n21832 = ~n21797 & n21831;
  assign n21833 = n21795 & n21832;
  assign n21834 = n21787 & n21833;
  assign n21835 = n21773 & n21834;
  assign n21836 = n21835 ^ n19104;
  assign n21837 = n21184 & n21212;
  assign n21838 = ~n21231 & n21241;
  assign n21839 = n21122 & ~n21838;
  assign n21840 = ~n21837 & ~n21839;
  assign n21841 = n21189 & ~n21732;
  assign n21842 = ~n21121 & ~n21723;
  assign n21843 = ~n21841 & ~n21842;
  assign n21844 = n21122 & n21187;
  assign n21845 = ~n21222 & n21237;
  assign n21846 = ~n21844 & ~n21845;
  assign n21847 = ~n21198 & n21717;
  assign n21848 = n21200 & ~n21847;
  assign n21849 = ~n21223 & n21241;
  assign n21850 = n21184 & ~n21849;
  assign n21851 = ~n21848 & ~n21850;
  assign n21852 = n21846 & n21851;
  assign n21853 = n21843 & n21852;
  assign n21854 = n21219 & n21853;
  assign n21855 = n21202 & n21854;
  assign n21856 = n21731 & n21855;
  assign n21857 = n21840 & n21856;
  assign n21858 = ~n21716 & n21857;
  assign n21859 = n21196 & n21858;
  assign n21860 = n21859 ^ n18781;
  assign n21861 = n19707 ^ x814;
  assign n21862 = n20837 ^ x819;
  assign n21863 = n21861 & n21862;
  assign n21864 = ~n21861 & ~n21862;
  assign n21865 = ~n21863 & ~n21864;
  assign n21866 = n21665 ^ x816;
  assign n21867 = n20708 ^ x818;
  assign n21868 = n21278 ^ x817;
  assign n21869 = n19570 ^ x815;
  assign n21870 = ~n21868 & ~n21869;
  assign n21871 = n21867 & n21870;
  assign n21872 = ~n21866 & n21871;
  assign n21873 = ~n21865 & n21872;
  assign n21874 = n21861 & ~n21862;
  assign n21875 = ~n21866 & ~n21867;
  assign n21876 = n21870 & n21875;
  assign n21877 = n21874 & n21876;
  assign n21878 = ~n21861 & n21862;
  assign n21879 = n21866 & ~n21867;
  assign n21880 = n21868 & n21869;
  assign n21881 = n21879 & n21880;
  assign n21882 = ~n21868 & n21869;
  assign n21883 = n21867 & n21882;
  assign n21884 = n21866 & n21883;
  assign n21885 = ~n21881 & ~n21884;
  assign n21886 = n21878 & ~n21885;
  assign n21887 = ~n21877 & ~n21886;
  assign n21888 = ~n21873 & n21887;
  assign n21889 = n21868 & ~n21869;
  assign n21890 = n21875 & n21889;
  assign n21891 = ~n21865 & n21890;
  assign n21892 = n21867 & n21889;
  assign n21893 = ~n21866 & n21892;
  assign n21894 = ~n21876 & ~n21893;
  assign n21895 = n21878 & ~n21894;
  assign n21896 = ~n21891 & ~n21895;
  assign n21897 = n21867 ^ n21866;
  assign n21898 = n21882 & n21897;
  assign n21899 = n21878 & n21898;
  assign n21900 = n21870 & n21879;
  assign n21901 = n21866 & n21892;
  assign n21902 = ~n21900 & ~n21901;
  assign n21903 = n21874 & ~n21902;
  assign n21904 = ~n21899 & ~n21903;
  assign n21905 = ~n21865 & ~n21902;
  assign n21906 = n21875 & n21882;
  assign n21907 = n21875 & n21880;
  assign n21908 = n21867 & n21880;
  assign n21909 = n21866 & n21908;
  assign n21910 = ~n21907 & ~n21909;
  assign n21911 = ~n21906 & n21910;
  assign n21912 = n21864 & ~n21911;
  assign n21915 = ~n21866 & n21908;
  assign n21916 = ~n21881 & ~n21915;
  assign n21917 = ~n21898 & n21916;
  assign n21913 = n21885 & ~n21906;
  assign n21914 = ~n21907 & n21913;
  assign n21918 = n21917 ^ n21914;
  assign n21919 = n21917 ^ n21862;
  assign n21920 = n21919 ^ n21917;
  assign n21921 = n21918 & n21920;
  assign n21922 = n21921 ^ n21917;
  assign n21923 = n21861 & ~n21922;
  assign n21924 = ~n21912 & ~n21923;
  assign n21925 = ~n21905 & n21924;
  assign n21928 = n21866 & n21871;
  assign n21926 = n21879 & n21889;
  assign n21927 = ~n21909 & ~n21926;
  assign n21929 = n21928 ^ n21927;
  assign n21930 = n21929 ^ n21928;
  assign n21931 = n21928 ^ n21861;
  assign n21932 = n21931 ^ n21928;
  assign n21933 = ~n21930 & ~n21932;
  assign n21934 = n21933 ^ n21928;
  assign n21935 = n21862 & n21934;
  assign n21936 = n21935 ^ n21928;
  assign n21937 = n21925 & ~n21936;
  assign n21938 = n21904 & n21937;
  assign n21939 = n21896 & n21938;
  assign n21940 = n21888 & n21939;
  assign n21941 = n21940 ^ n19500;
  assign n21942 = n21878 & n21881;
  assign n21943 = ~n21865 & n21871;
  assign n21944 = ~n21942 & ~n21943;
  assign n21945 = n21864 & n21926;
  assign n21946 = n21874 & n21893;
  assign n21947 = ~n21945 & ~n21946;
  assign n21948 = n21944 & n21947;
  assign n21949 = n21864 & ~n21885;
  assign n21950 = ~n21907 & ~n21915;
  assign n21951 = n21950 ^ n21863;
  assign n21952 = n21950 ^ n21864;
  assign n21953 = n21952 ^ n21864;
  assign n21954 = n21879 & n21882;
  assign n21955 = ~n21884 & ~n21954;
  assign n21956 = n21955 ^ n21864;
  assign n21957 = n21953 & n21956;
  assign n21958 = n21957 ^ n21864;
  assign n21959 = ~n21951 & n21958;
  assign n21960 = n21959 ^ n21863;
  assign n21961 = ~n21949 & ~n21960;
  assign n21962 = ~n21898 & n21910;
  assign n21963 = n21874 & ~n21962;
  assign n21964 = ~n21890 & n21902;
  assign n21965 = ~n21893 & n21964;
  assign n21966 = n21878 & ~n21965;
  assign n21967 = ~n21963 & ~n21966;
  assign n21968 = n21961 & n21967;
  assign n21969 = n21906 ^ n21863;
  assign n21970 = n21969 ^ n21906;
  assign n21971 = ~n21876 & ~n21890;
  assign n21972 = n21971 ^ n21906;
  assign n21973 = n21970 & ~n21972;
  assign n21974 = n21973 ^ n21906;
  assign n21975 = n21968 & ~n21974;
  assign n21976 = n21948 & n21975;
  assign n21977 = n21904 & n21976;
  assign n21978 = n21977 ^ n19847;
  assign n21979 = n20790 & n20915;
  assign n21980 = ~n20943 & ~n21044;
  assign n21981 = ~n21979 & ~n21980;
  assign n21982 = ~n20939 & n20966;
  assign n21983 = n20917 & n21982;
  assign n21984 = ~n20928 & ~n20950;
  assign n21985 = n21984 ^ n20789;
  assign n21986 = n21985 ^ n21984;
  assign n21987 = ~n20930 & n21019;
  assign n21988 = n21987 ^ n21984;
  assign n21989 = ~n21986 & n21988;
  assign n21990 = n21989 ^ n21984;
  assign n21991 = ~n20763 & ~n21990;
  assign n21992 = ~n21983 & ~n21991;
  assign n21993 = n21981 & n21992;
  assign n21994 = n20945 & n21993;
  assign n21995 = n20938 & n21994;
  assign n21996 = n21030 & n21995;
  assign n21997 = n21996 ^ n19034;
  assign n21998 = n20488 ^ x802;
  assign n22017 = n20258 ^ x807;
  assign n21999 = n19317 ^ x806;
  assign n22000 = n21110 ^ x805;
  assign n22001 = n21999 & ~n22000;
  assign n22002 = n20378 ^ x803;
  assign n22003 = n21608 ^ x804;
  assign n22004 = ~n22002 & ~n22003;
  assign n22005 = n22001 & n22004;
  assign n22006 = ~n22002 & n22003;
  assign n22007 = n22000 & n22006;
  assign n22008 = ~n21999 & n22000;
  assign n22009 = n22008 ^ n22003;
  assign n22010 = n22009 ^ n22003;
  assign n22011 = n22002 & n22003;
  assign n22012 = n22011 ^ n22003;
  assign n22013 = ~n22010 & ~n22012;
  assign n22014 = n22013 ^ n22003;
  assign n22015 = ~n22007 & n22014;
  assign n22016 = ~n22005 & n22015;
  assign n22018 = n22017 ^ n22016;
  assign n22019 = n22018 ^ n22016;
  assign n22020 = ~n22001 & n22006;
  assign n22021 = n21999 & n22000;
  assign n22022 = n22002 & ~n22003;
  assign n22023 = ~n22021 & n22022;
  assign n22024 = ~n22020 & ~n22023;
  assign n22025 = ~n21999 & ~n22000;
  assign n22026 = n22011 & n22025;
  assign n22027 = n22004 & n22021;
  assign n22028 = ~n22026 & ~n22027;
  assign n22029 = n22024 & n22028;
  assign n22030 = n22029 ^ n22016;
  assign n22031 = ~n22019 & n22030;
  assign n22032 = n22031 ^ n22016;
  assign n22033 = ~n21998 & ~n22032;
  assign n22034 = n22003 ^ n22002;
  assign n22035 = n22034 ^ n22002;
  assign n22036 = n22002 ^ n21999;
  assign n22037 = n22036 ^ n22003;
  assign n22038 = n22037 ^ n22002;
  assign n22039 = n22038 ^ n22002;
  assign n22040 = n22035 & n22039;
  assign n22041 = n22040 ^ n22002;
  assign n22042 = ~n22000 & n22041;
  assign n22043 = n22042 ^ n22037;
  assign n22044 = n22043 ^ n22017;
  assign n22045 = n22044 ^ n22043;
  assign n22046 = ~n22021 & ~n22025;
  assign n22047 = n22002 & ~n22046;
  assign n22048 = ~n22020 & ~n22047;
  assign n22049 = ~n22005 & n22048;
  assign n22050 = n22049 ^ n22043;
  assign n22051 = ~n22045 & ~n22050;
  assign n22052 = n22051 ^ n22043;
  assign n22053 = n21998 & ~n22052;
  assign n22054 = ~n22033 & ~n22053;
  assign n22055 = n22054 ^ n17493;
  assign n22056 = n21776 & ~n21809;
  assign n22057 = n21771 & n21801;
  assign n22058 = n21765 ^ n21764;
  assign n22059 = n21765 ^ n21763;
  assign n22060 = n22059 ^ n21763;
  assign n22061 = n21822 ^ n21763;
  assign n22062 = n22060 & n22061;
  assign n22063 = n22062 ^ n21763;
  assign n22064 = n22058 & n22063;
  assign n22065 = ~n22057 & ~n22064;
  assign n22066 = ~n22056 & n22065;
  assign n22067 = ~n21774 & ~n21817;
  assign n22068 = n21825 & ~n22067;
  assign n22069 = ~n21796 & ~n21823;
  assign n22070 = ~n21788 & ~n21792;
  assign n22071 = n22069 & n22070;
  assign n22072 = n21771 & ~n22071;
  assign n22073 = ~n22068 & ~n22072;
  assign n22074 = ~n21801 & ~n21808;
  assign n22075 = n21778 & ~n22074;
  assign n22076 = n21809 & n21819;
  assign n22077 = n21766 & ~n22076;
  assign n22078 = ~n21781 & n22069;
  assign n22079 = ~n21770 & n22078;
  assign n22080 = n21778 & ~n22079;
  assign n22081 = ~n21822 & n22070;
  assign n22082 = ~n21783 & n22081;
  assign n22083 = n21776 & ~n22082;
  assign n22084 = ~n22080 & ~n22083;
  assign n22085 = ~n22077 & n22084;
  assign n22086 = ~n22075 & n22085;
  assign n22087 = n22073 & n22086;
  assign n22088 = n22066 & n22087;
  assign n22089 = n21807 & n22088;
  assign n22090 = n21773 & n22089;
  assign n22091 = n22090 ^ n19367;
  assign n22092 = n20297 ^ n19318;
  assign n22093 = n22092 ^ n20297;
  assign n22094 = n20306 ^ n20297;
  assign n22095 = n22094 ^ n20297;
  assign n22096 = n22093 & ~n22095;
  assign n22097 = n22096 ^ n20297;
  assign n22098 = n19571 & n22097;
  assign n22099 = n22098 ^ n20297;
  assign n22100 = ~n20275 & ~n22099;
  assign n22101 = ~n20292 & n21624;
  assign n22102 = n20263 & ~n22101;
  assign n22103 = ~n20304 & n20316;
  assign n22104 = ~n20261 & n22103;
  assign n22105 = n20276 & ~n22104;
  assign n22106 = ~n22102 & ~n22105;
  assign n22107 = ~n19571 & n20274;
  assign n22108 = ~n20284 & ~n20308;
  assign n22109 = n19572 & ~n22108;
  assign n22110 = ~n20283 & n20317;
  assign n22111 = n20294 & ~n22110;
  assign n22112 = ~n22109 & ~n22111;
  assign n22113 = ~n22107 & n22112;
  assign n22114 = n22106 & n22113;
  assign n22115 = ~n20286 & n22114;
  assign n22116 = n20300 & n22115;
  assign n22117 = n20296 & n22116;
  assign n22118 = n22100 & n22117;
  assign n22119 = n21611 & n22118;
  assign n22120 = n20271 & n22119;
  assign n22121 = n22120 ^ n20181;
  assign n22122 = ~n21872 & ~n21900;
  assign n22123 = n21878 & ~n22122;
  assign n22124 = n21861 & n21872;
  assign n22125 = ~n21906 & ~n21915;
  assign n22126 = ~n21901 & n22125;
  assign n22127 = ~n21898 & n22126;
  assign n22128 = n21863 & ~n22127;
  assign n22129 = ~n22124 & ~n22128;
  assign n22130 = ~n21865 & n21926;
  assign n22131 = n21874 & ~n21964;
  assign n22132 = ~n22130 & ~n22131;
  assign n22133 = n22129 & n22132;
  assign n22134 = n21885 & n22125;
  assign n22135 = n21878 & ~n22134;
  assign n22136 = ~n21893 & ~n21928;
  assign n22137 = n21864 & ~n22136;
  assign n22138 = ~n21864 & n22125;
  assign n22139 = ~n21909 & n22138;
  assign n22140 = ~n21881 & n22139;
  assign n22141 = ~n21874 & ~n21883;
  assign n22142 = ~n22134 & ~n22141;
  assign n22143 = n21910 & ~n22142;
  assign n22144 = ~n21954 & n22143;
  assign n22145 = ~n22140 & ~n22144;
  assign n22146 = ~n21862 & n22145;
  assign n22147 = ~n22137 & ~n22146;
  assign n22148 = ~n22135 & n22147;
  assign n22149 = n22133 & n22148;
  assign n22150 = n21896 & n22149;
  assign n22151 = ~n22123 & n22150;
  assign n22152 = n22151 ^ n19067;
  assign n22153 = n21878 & n21907;
  assign n22154 = ~n21865 & n21900;
  assign n22155 = ~n22153 & ~n22154;
  assign n22156 = ~n21862 & n21893;
  assign n22157 = ~n21890 & ~n21901;
  assign n22158 = n21874 & ~n22157;
  assign n22159 = ~n22156 & ~n22158;
  assign n22160 = n22155 & n22159;
  assign n22161 = ~n21861 & n21883;
  assign n22162 = ~n21926 & ~n21928;
  assign n22163 = n21863 & ~n22162;
  assign n22164 = ~n21901 & ~n21926;
  assign n22165 = n21878 & ~n22164;
  assign n22166 = n21913 & ~n21954;
  assign n22167 = n21874 & ~n22166;
  assign n22168 = ~n21863 & n21885;
  assign n22169 = ~n22138 & ~n22168;
  assign n22170 = n21910 & ~n22169;
  assign n22171 = ~n21865 & ~n22170;
  assign n22172 = ~n22167 & ~n22171;
  assign n22173 = ~n22165 & n22172;
  assign n22174 = ~n22123 & n22173;
  assign n22175 = ~n22163 & n22174;
  assign n22176 = ~n22161 & n22175;
  assign n22177 = n22160 & n22176;
  assign n22178 = n21888 & n22177;
  assign n22179 = n22178 ^ n18452;
  assign n22180 = n21200 & ~n21733;
  assign n22181 = n21184 & ~n21193;
  assign n22182 = ~n22180 & ~n22181;
  assign n22183 = n21198 & ~n21222;
  assign n22184 = n21227 & n21723;
  assign n22185 = ~n21215 & n22184;
  assign n22186 = ~n21237 & n22185;
  assign n22187 = ~n21187 & n22186;
  assign n22188 = n21189 & ~n22187;
  assign n22189 = ~n22183 & ~n22188;
  assign n22190 = n22182 & n22189;
  assign n22191 = ~n21183 & n22190;
  assign n22192 = n21207 & n22191;
  assign n22193 = n21726 & n22192;
  assign n22194 = n21840 & n22193;
  assign n22195 = n21719 & n22194;
  assign n22196 = ~n21716 & n22195;
  assign n22197 = n22196 ^ n20414;
  assign n22198 = n21766 & ~n22070;
  assign n22199 = n21817 & ~n21825;
  assign n22200 = ~n22198 & ~n22199;
  assign n22201 = n21771 & n21774;
  assign n22202 = n21778 & ~n21802;
  assign n22203 = n21776 & ~n22074;
  assign n22204 = ~n21770 & ~n21822;
  assign n22205 = n21778 & ~n22204;
  assign n22206 = ~n21792 & ~n21817;
  assign n22207 = ~n21771 & n22206;
  assign n22208 = ~n21781 & ~n21796;
  assign n22209 = ~n21822 & n22208;
  assign n22210 = ~n21776 & n22209;
  assign n22211 = ~n22207 & ~n22210;
  assign n22212 = ~n21788 & ~n22211;
  assign n22213 = n21825 & ~n22212;
  assign n22214 = ~n22205 & ~n22213;
  assign n22215 = ~n22203 & n22214;
  assign n22216 = n21810 ^ n21778;
  assign n22217 = n22216 ^ n21810;
  assign n22218 = ~n21804 & ~n21818;
  assign n22219 = n22218 ^ n21810;
  assign n22220 = n22219 ^ n21810;
  assign n22221 = ~n22217 & ~n22220;
  assign n22222 = n22221 ^ n21810;
  assign n22223 = ~n21766 & ~n22222;
  assign n22224 = n22223 ^ n21810;
  assign n22225 = n22215 & n22224;
  assign n22226 = n21787 & n22225;
  assign n22227 = ~n22202 & n22226;
  assign n22228 = ~n22201 & n22227;
  assign n22229 = n22200 & n22228;
  assign n22230 = n22065 & n22229;
  assign n22231 = n22230 ^ n20150;
  assign n22232 = ~n21998 & n22017;
  assign n22233 = n22008 & n22011;
  assign n22234 = n22006 & n22025;
  assign n22235 = ~n22233 & ~n22234;
  assign n22236 = n21999 & n22006;
  assign n22237 = n22001 & n22002;
  assign n22238 = ~n22003 & n22008;
  assign n22239 = ~n22237 & ~n22238;
  assign n22240 = ~n22236 & n22239;
  assign n22241 = n22235 & n22240;
  assign n22242 = n22232 & ~n22241;
  assign n22243 = n21998 & n22017;
  assign n22244 = n22011 & ~n22025;
  assign n22245 = ~n22002 & n22025;
  assign n22246 = ~n22003 & n22021;
  assign n22247 = ~n22245 & ~n22246;
  assign n22248 = ~n22005 & n22247;
  assign n22249 = ~n22244 & n22248;
  assign n22250 = n22243 & ~n22249;
  assign n22251 = ~n22242 & ~n22250;
  assign n22252 = ~n21998 & ~n22017;
  assign n22253 = n22006 & n22008;
  assign n22254 = n22011 ^ n22001;
  assign n22255 = n22254 ^ n22011;
  assign n22256 = n22022 ^ n22011;
  assign n22257 = ~n22255 & n22256;
  assign n22258 = n22257 ^ n22011;
  assign n22259 = ~n22253 & ~n22258;
  assign n22260 = n22235 & n22259;
  assign n22261 = ~n22005 & n22260;
  assign n22262 = n22252 & n22261;
  assign n22263 = n21998 & ~n22017;
  assign n22264 = n22001 & n22022;
  assign n22265 = n22000 & n22004;
  assign n22266 = n22003 & ~n22046;
  assign n22267 = ~n22265 & ~n22266;
  assign n22268 = ~n22264 & n22267;
  assign n22269 = n22235 & n22268;
  assign n22270 = n22263 & n22269;
  assign n22271 = ~n22262 & ~n22270;
  assign n22272 = n22251 & n22271;
  assign n22273 = n22272 ^ n18892;
  assign n22274 = ~n21799 & n21819;
  assign n22275 = n21778 & ~n22274;
  assign n22276 = n21778 & n21779;
  assign n22277 = n21771 & ~n22081;
  assign n22278 = ~n22276 & ~n22277;
  assign n22279 = n21793 & n22069;
  assign n22280 = n21776 & ~n22279;
  assign n22281 = n21760 ^ n21758;
  assign n22282 = n21759 ^ n21758;
  assign n22283 = ~n22281 & n22282;
  assign n22284 = n22283 ^ n21758;
  assign n22285 = n21759 ^ n21757;
  assign n22286 = n22285 ^ n21760;
  assign n22287 = n22286 ^ n21758;
  assign n22288 = n22287 ^ n21759;
  assign n22289 = n22288 ^ n21760;
  assign n22290 = ~n22284 & ~n22289;
  assign n22291 = n22290 ^ n22286;
  assign n22292 = n21766 & ~n22291;
  assign n22293 = ~n22280 & ~n22292;
  assign n22294 = n22278 & n22293;
  assign n22295 = n21773 & n22294;
  assign n22296 = ~n22275 & n22295;
  assign n22297 = ~n21774 & ~n21801;
  assign n22298 = n22297 ^ n21765;
  assign n22299 = n22298 ^ n22297;
  assign n22300 = ~n21763 & n21819;
  assign n22301 = n22300 ^ n22297;
  assign n22302 = n22299 & n22301;
  assign n22303 = n22302 ^ n22297;
  assign n22304 = ~n22058 & ~n22303;
  assign n22305 = n22296 & ~n22304;
  assign n22306 = n22066 & n22305;
  assign n22307 = n22306 ^ n18182;
  assign n22308 = n22029 & n22232;
  assign n22309 = ~n22016 & n22252;
  assign n22310 = ~n22308 & ~n22309;
  assign n22311 = ~n22043 & n22263;
  assign n22312 = ~n22049 & n22243;
  assign n22313 = ~n22311 & ~n22312;
  assign n22314 = n22310 & n22313;
  assign n22315 = n22314 ^ n20389;
  assign n22316 = n21999 & n22011;
  assign n22317 = n22248 & ~n22316;
  assign n22318 = n22263 & ~n22317;
  assign n22319 = n22232 & ~n22261;
  assign n22320 = ~n22318 & ~n22319;
  assign n22321 = ~n22240 & n22252;
  assign n22322 = n22243 & ~n22269;
  assign n22323 = ~n22321 & ~n22322;
  assign n22324 = n22320 & n22323;
  assign n22325 = n22235 & n22324;
  assign n22326 = n22325 ^ n19331;
  assign n22327 = n21316 & ~n21510;
  assign n22328 = ~n21532 & ~n22327;
  assign n22329 = n21434 & n21444;
  assign n22330 = n21424 & ~n21472;
  assign n22331 = ~n22329 & ~n22330;
  assign n22332 = ~n21422 & n21461;
  assign n22333 = n21444 & ~n22332;
  assign n22334 = n21456 & ~n21511;
  assign n22335 = ~n21279 & n21441;
  assign n22336 = ~n21446 & ~n21458;
  assign n22337 = n21316 & ~n22336;
  assign n22338 = ~n22335 & ~n22337;
  assign n22339 = ~n21445 & ~n21460;
  assign n22340 = ~n21446 & n22339;
  assign n22341 = n21424 & ~n22340;
  assign n22342 = ~n21448 & ~n21456;
  assign n22343 = n21450 & ~n21459;
  assign n22344 = ~n21422 & n22343;
  assign n22345 = ~n22342 & ~n22344;
  assign n22346 = ~n22341 & ~n22345;
  assign n22347 = n22338 & n22346;
  assign n22348 = ~n22334 & n22347;
  assign n22349 = ~n22333 & n22348;
  assign n22350 = n21439 & n22349;
  assign n22351 = n21494 & n22350;
  assign n22352 = n22331 & n22351;
  assign n22353 = n22328 & n22352;
  assign n22354 = n22353 ^ n18930;
  assign n22355 = n21437 & n21456;
  assign n22356 = ~n21475 & n22343;
  assign n22357 = n21316 & ~n22356;
  assign n22358 = ~n21315 & ~n21473;
  assign n22359 = n21446 & n21456;
  assign n22360 = ~n21424 & ~n22359;
  assign n22361 = ~n21460 & n22336;
  assign n22362 = ~n22360 & ~n22361;
  assign n22363 = ~n22358 & ~n22362;
  assign n22364 = ~n21448 & n22336;
  assign n22365 = n21444 & ~n22364;
  assign n22366 = n21456 ^ n21422;
  assign n22367 = n21424 ^ n21422;
  assign n22368 = n22367 ^ n21424;
  assign n22369 = n21461 ^ n21424;
  assign n22370 = ~n22368 & n22369;
  assign n22371 = n22370 ^ n21424;
  assign n22372 = n22366 & n22371;
  assign n22373 = n22372 ^ n21456;
  assign n22374 = ~n22365 & ~n22373;
  assign n22375 = n22363 & n22374;
  assign n22376 = ~n22357 & n22375;
  assign n22377 = ~n22355 & n22376;
  assign n22378 = n22331 & n22377;
  assign n22379 = n21433 & n22378;
  assign n22380 = n22328 & n22379;
  assign n22381 = n22380 ^ n17953;
  assign n22382 = n20276 & ~n21624;
  assign n22383 = ~n20261 & n21628;
  assign n22384 = n20294 & ~n22383;
  assign n22385 = n20318 & n21616;
  assign n22386 = n19572 & ~n22385;
  assign n22387 = ~n22384 & ~n22386;
  assign n22388 = ~n22382 & n22387;
  assign n22389 = ~n20268 & n20310;
  assign n22390 = n20306 & n22389;
  assign n22391 = n22390 ^ n20292;
  assign n22392 = n22391 ^ n20292;
  assign n22393 = n20292 ^ n19571;
  assign n22394 = n22393 ^ n20292;
  assign n22395 = ~n22392 & ~n22394;
  assign n22396 = n22395 ^ n20292;
  assign n22397 = n20278 & n22396;
  assign n22398 = n22397 ^ n20292;
  assign n22399 = n22388 & ~n22398;
  assign n22400 = ~n21613 & n22399;
  assign n22401 = n20287 & n22400;
  assign n22402 = n22100 & n22401;
  assign n22403 = n22402 ^ n19943;
  assign y0 = n18858;
  assign y1 = n20337;
  assign y2 = n19317;
  assign y3 = n20672;
  assign y4 = n20708;
  assign y5 = n20740;
  assign y6 = n20762;
  assign y7 = n20980;
  assign y8 = n21017;
  assign y9 = n21067;
  assign y10 = n21110;
  assign y11 = n21257;
  assign y12 = n21278;
  assign y13 = n21491;
  assign y14 = n21179;
  assign y15 = n21535;
  assign y16 = n21554;
  assign y17 = n21586;
  assign y18 = n21608;
  assign y19 = n21641;
  assign y20 = n21665;
  assign y21 = n21690;
  assign y22 = n21147;
  assign y23 = n21715;
  assign y24 = n21314;
  assign y25 = n21756;
  assign y26 = n20378;
  assign y27 = n21836;
  assign y28 = n19570;
  assign y29 = n21860;
  assign y30 = n20788;
  assign y31 = n21941;
  assign y32 = n21384;
  assign y33 = n21978;
  assign y34 = n20488;
  assign y35 = n21997;
  assign y36 = n19707;
  assign y37 = ~n22055;
  assign y38 = n20876;
  assign y39 = n22091;
  assign y40 = n21353;
  assign y41 = n22121;
  assign y42 = n20525;
  assign y43 = n22152;
  assign y44 = n20118;
  assign y45 = n22179;
  assign y46 = n20908;
  assign y47 = n22197;
  assign y48 = n21419;
  assign y49 = n22231;
  assign y50 = n20565;
  assign y51 = ~n22273;
  assign y52 = n19913;
  assign y53 = n22307;
  assign y54 = n20798;
  assign y55 = n22315;
  assign y56 = n21119;
  assign y57 = n22326;
  assign y58 = n20603;
  assign y59 = n22354;
  assign y60 = n20258;
  assign y61 = n22381;
  assign y62 = n20837;
  assign y63 = n22403;
endmodule
